// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Feb 24 2020 16:35:41

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    TX,
    SDA,
    SCL,
    RX,
    NEOPXL,
    LED,
    INLC,
    INLB,
    INLA,
    INHC,
    INHB,
    INHA,
    HALL3,
    HALL2,
    HALL1,
    FAULT_N,
    ENCODER1_B,
    ENCODER1_A,
    ENCODER0_B,
    ENCODER0_A,
    DE,
    CS_MISO,
    CS_CLK,
    CS,
    CLK);

    inout USBPU;
    inout TX;
    inout SDA;
    inout SCL;
    inout RX;
    output NEOPXL;
    output LED;
    inout INLC;
    inout INLB;
    inout INLA;
    inout INHC;
    inout INHB;
    inout INHA;
    inout HALL3;
    inout HALL2;
    inout HALL1;
    inout FAULT_N;
    inout ENCODER1_B;
    inout ENCODER1_A;
    inout ENCODER0_B;
    inout ENCODER0_A;
    inout DE;
    inout CS_MISO;
    inout CS_CLK;
    inout CS;
    input CLK;

    wire N__51103;
    wire N__51102;
    wire N__51101;
    wire N__51094;
    wire N__51093;
    wire N__51092;
    wire N__51085;
    wire N__51084;
    wire N__51083;
    wire N__51076;
    wire N__51075;
    wire N__51074;
    wire N__51067;
    wire N__51066;
    wire N__51065;
    wire N__51058;
    wire N__51057;
    wire N__51056;
    wire N__51049;
    wire N__51048;
    wire N__51047;
    wire N__51040;
    wire N__51039;
    wire N__51038;
    wire N__51031;
    wire N__51030;
    wire N__51029;
    wire N__51022;
    wire N__51021;
    wire N__51020;
    wire N__51013;
    wire N__51012;
    wire N__51011;
    wire N__51004;
    wire N__51003;
    wire N__51002;
    wire N__50995;
    wire N__50994;
    wire N__50993;
    wire N__50986;
    wire N__50985;
    wire N__50984;
    wire N__50977;
    wire N__50976;
    wire N__50975;
    wire N__50968;
    wire N__50967;
    wire N__50966;
    wire N__50959;
    wire N__50958;
    wire N__50957;
    wire N__50950;
    wire N__50949;
    wire N__50948;
    wire N__50941;
    wire N__50940;
    wire N__50939;
    wire N__50932;
    wire N__50931;
    wire N__50930;
    wire N__50923;
    wire N__50922;
    wire N__50921;
    wire N__50914;
    wire N__50913;
    wire N__50912;
    wire N__50905;
    wire N__50904;
    wire N__50903;
    wire N__50896;
    wire N__50895;
    wire N__50894;
    wire N__50887;
    wire N__50886;
    wire N__50885;
    wire N__50878;
    wire N__50877;
    wire N__50876;
    wire N__50859;
    wire N__50856;
    wire N__50853;
    wire N__50850;
    wire N__50847;
    wire N__50844;
    wire N__50841;
    wire N__50838;
    wire N__50835;
    wire N__50832;
    wire N__50829;
    wire N__50826;
    wire N__50823;
    wire N__50820;
    wire N__50817;
    wire N__50816;
    wire N__50815;
    wire N__50812;
    wire N__50809;
    wire N__50806;
    wire N__50803;
    wire N__50800;
    wire N__50797;
    wire N__50790;
    wire N__50787;
    wire N__50784;
    wire N__50781;
    wire N__50778;
    wire N__50777;
    wire N__50774;
    wire N__50773;
    wire N__50772;
    wire N__50771;
    wire N__50770;
    wire N__50767;
    wire N__50762;
    wire N__50761;
    wire N__50760;
    wire N__50759;
    wire N__50758;
    wire N__50757;
    wire N__50756;
    wire N__50755;
    wire N__50754;
    wire N__50753;
    wire N__50752;
    wire N__50749;
    wire N__50744;
    wire N__50739;
    wire N__50734;
    wire N__50731;
    wire N__50730;
    wire N__50727;
    wire N__50726;
    wire N__50723;
    wire N__50722;
    wire N__50721;
    wire N__50718;
    wire N__50715;
    wire N__50714;
    wire N__50713;
    wire N__50712;
    wire N__50709;
    wire N__50706;
    wire N__50703;
    wire N__50696;
    wire N__50691;
    wire N__50688;
    wire N__50687;
    wire N__50684;
    wire N__50675;
    wire N__50670;
    wire N__50665;
    wire N__50662;
    wire N__50659;
    wire N__50656;
    wire N__50653;
    wire N__50648;
    wire N__50645;
    wire N__50642;
    wire N__50633;
    wire N__50616;
    wire N__50615;
    wire N__50612;
    wire N__50611;
    wire N__50608;
    wire N__50607;
    wire N__50604;
    wire N__50599;
    wire N__50596;
    wire N__50595;
    wire N__50590;
    wire N__50587;
    wire N__50584;
    wire N__50579;
    wire N__50574;
    wire N__50573;
    wire N__50570;
    wire N__50569;
    wire N__50568;
    wire N__50567;
    wire N__50566;
    wire N__50565;
    wire N__50564;
    wire N__50563;
    wire N__50562;
    wire N__50559;
    wire N__50558;
    wire N__50557;
    wire N__50556;
    wire N__50555;
    wire N__50554;
    wire N__50551;
    wire N__50548;
    wire N__50545;
    wire N__50544;
    wire N__50541;
    wire N__50538;
    wire N__50537;
    wire N__50536;
    wire N__50535;
    wire N__50534;
    wire N__50533;
    wire N__50532;
    wire N__50531;
    wire N__50528;
    wire N__50525;
    wire N__50520;
    wire N__50517;
    wire N__50512;
    wire N__50509;
    wire N__50506;
    wire N__50503;
    wire N__50500;
    wire N__50499;
    wire N__50496;
    wire N__50493;
    wire N__50492;
    wire N__50491;
    wire N__50490;
    wire N__50487;
    wire N__50482;
    wire N__50479;
    wire N__50476;
    wire N__50473;
    wire N__50470;
    wire N__50467;
    wire N__50462;
    wire N__50459;
    wire N__50454;
    wire N__50449;
    wire N__50446;
    wire N__50445;
    wire N__50444;
    wire N__50437;
    wire N__50434;
    wire N__50429;
    wire N__50424;
    wire N__50421;
    wire N__50418;
    wire N__50411;
    wire N__50398;
    wire N__50393;
    wire N__50388;
    wire N__50385;
    wire N__50378;
    wire N__50369;
    wire N__50358;
    wire N__50357;
    wire N__50356;
    wire N__50355;
    wire N__50354;
    wire N__50353;
    wire N__50352;
    wire N__50349;
    wire N__50348;
    wire N__50347;
    wire N__50346;
    wire N__50345;
    wire N__50344;
    wire N__50343;
    wire N__50342;
    wire N__50339;
    wire N__50338;
    wire N__50337;
    wire N__50336;
    wire N__50335;
    wire N__50334;
    wire N__50333;
    wire N__50332;
    wire N__50329;
    wire N__50328;
    wire N__50327;
    wire N__50322;
    wire N__50317;
    wire N__50316;
    wire N__50315;
    wire N__50310;
    wire N__50305;
    wire N__50298;
    wire N__50295;
    wire N__50292;
    wire N__50289;
    wire N__50288;
    wire N__50287;
    wire N__50286;
    wire N__50285;
    wire N__50284;
    wire N__50281;
    wire N__50272;
    wire N__50269;
    wire N__50266;
    wire N__50265;
    wire N__50264;
    wire N__50263;
    wire N__50262;
    wire N__50257;
    wire N__50256;
    wire N__50253;
    wire N__50250;
    wire N__50247;
    wire N__50244;
    wire N__50241;
    wire N__50236;
    wire N__50231;
    wire N__50224;
    wire N__50217;
    wire N__50212;
    wire N__50209;
    wire N__50206;
    wire N__50205;
    wire N__50204;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50188;
    wire N__50185;
    wire N__50182;
    wire N__50173;
    wire N__50164;
    wire N__50159;
    wire N__50154;
    wire N__50147;
    wire N__50130;
    wire N__50129;
    wire N__50128;
    wire N__50127;
    wire N__50126;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50116;
    wire N__50113;
    wire N__50110;
    wire N__50107;
    wire N__50104;
    wire N__50099;
    wire N__50094;
    wire N__50089;
    wire N__50086;
    wire N__50079;
    wire N__50078;
    wire N__50077;
    wire N__50076;
    wire N__50075;
    wire N__50072;
    wire N__50069;
    wire N__50068;
    wire N__50067;
    wire N__50066;
    wire N__50063;
    wire N__50060;
    wire N__50057;
    wire N__50054;
    wire N__50051;
    wire N__50048;
    wire N__50045;
    wire N__50044;
    wire N__50041;
    wire N__50038;
    wire N__50035;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50023;
    wire N__50020;
    wire N__50017;
    wire N__50016;
    wire N__50015;
    wire N__50014;
    wire N__50011;
    wire N__50008;
    wire N__50007;
    wire N__50006;
    wire N__50005;
    wire N__50002;
    wire N__50001;
    wire N__50000;
    wire N__49999;
    wire N__49996;
    wire N__49993;
    wire N__49990;
    wire N__49987;
    wire N__49986;
    wire N__49985;
    wire N__49984;
    wire N__49979;
    wire N__49974;
    wire N__49971;
    wire N__49968;
    wire N__49965;
    wire N__49962;
    wire N__49957;
    wire N__49956;
    wire N__49955;
    wire N__49954;
    wire N__49951;
    wire N__49948;
    wire N__49943;
    wire N__49942;
    wire N__49941;
    wire N__49934;
    wire N__49931;
    wire N__49924;
    wire N__49923;
    wire N__49920;
    wire N__49915;
    wire N__49906;
    wire N__49903;
    wire N__49898;
    wire N__49893;
    wire N__49890;
    wire N__49885;
    wire N__49878;
    wire N__49875;
    wire N__49868;
    wire N__49851;
    wire N__49850;
    wire N__49847;
    wire N__49844;
    wire N__49843;
    wire N__49842;
    wire N__49839;
    wire N__49838;
    wire N__49835;
    wire N__49834;
    wire N__49831;
    wire N__49830;
    wire N__49829;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49819;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49811;
    wire N__49808;
    wire N__49807;
    wire N__49804;
    wire N__49803;
    wire N__49800;
    wire N__49797;
    wire N__49796;
    wire N__49793;
    wire N__49790;
    wire N__49787;
    wire N__49784;
    wire N__49779;
    wire N__49776;
    wire N__49775;
    wire N__49774;
    wire N__49773;
    wire N__49772;
    wire N__49771;
    wire N__49768;
    wire N__49765;
    wire N__49762;
    wire N__49759;
    wire N__49758;
    wire N__49757;
    wire N__49754;
    wire N__49753;
    wire N__49752;
    wire N__49751;
    wire N__49750;
    wire N__49749;
    wire N__49746;
    wire N__49743;
    wire N__49738;
    wire N__49735;
    wire N__49730;
    wire N__49723;
    wire N__49722;
    wire N__49719;
    wire N__49716;
    wire N__49713;
    wire N__49704;
    wire N__49701;
    wire N__49698;
    wire N__49697;
    wire N__49694;
    wire N__49691;
    wire N__49688;
    wire N__49685;
    wire N__49680;
    wire N__49677;
    wire N__49674;
    wire N__49665;
    wire N__49662;
    wire N__49659;
    wire N__49656;
    wire N__49649;
    wire N__49646;
    wire N__49643;
    wire N__49638;
    wire N__49633;
    wire N__49620;
    wire N__49615;
    wire N__49602;
    wire N__49601;
    wire N__49600;
    wire N__49597;
    wire N__49594;
    wire N__49593;
    wire N__49590;
    wire N__49589;
    wire N__49588;
    wire N__49585;
    wire N__49582;
    wire N__49581;
    wire N__49580;
    wire N__49577;
    wire N__49574;
    wire N__49571;
    wire N__49570;
    wire N__49567;
    wire N__49564;
    wire N__49561;
    wire N__49558;
    wire N__49555;
    wire N__49554;
    wire N__49553;
    wire N__49548;
    wire N__49545;
    wire N__49542;
    wire N__49539;
    wire N__49536;
    wire N__49533;
    wire N__49528;
    wire N__49527;
    wire N__49526;
    wire N__49525;
    wire N__49524;
    wire N__49521;
    wire N__49518;
    wire N__49517;
    wire N__49516;
    wire N__49511;
    wire N__49510;
    wire N__49509;
    wire N__49508;
    wire N__49503;
    wire N__49498;
    wire N__49495;
    wire N__49490;
    wire N__49489;
    wire N__49484;
    wire N__49481;
    wire N__49478;
    wire N__49475;
    wire N__49472;
    wire N__49469;
    wire N__49466;
    wire N__49463;
    wire N__49460;
    wire N__49455;
    wire N__49450;
    wire N__49447;
    wire N__49444;
    wire N__49435;
    wire N__49426;
    wire N__49413;
    wire N__49412;
    wire N__49411;
    wire N__49410;
    wire N__49407;
    wire N__49406;
    wire N__49403;
    wire N__49396;
    wire N__49393;
    wire N__49390;
    wire N__49387;
    wire N__49384;
    wire N__49381;
    wire N__49378;
    wire N__49375;
    wire N__49368;
    wire N__49365;
    wire N__49362;
    wire N__49359;
    wire N__49356;
    wire N__49353;
    wire N__49350;
    wire N__49349;
    wire N__49346;
    wire N__49343;
    wire N__49340;
    wire N__49337;
    wire N__49334;
    wire N__49331;
    wire N__49326;
    wire N__49323;
    wire N__49320;
    wire N__49317;
    wire N__49314;
    wire N__49311;
    wire N__49308;
    wire N__49305;
    wire N__49302;
    wire N__49299;
    wire N__49296;
    wire N__49293;
    wire N__49290;
    wire N__49287;
    wire N__49284;
    wire N__49283;
    wire N__49280;
    wire N__49277;
    wire N__49272;
    wire N__49269;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49259;
    wire N__49256;
    wire N__49253;
    wire N__49250;
    wire N__49247;
    wire N__49242;
    wire N__49239;
    wire N__49236;
    wire N__49233;
    wire N__49230;
    wire N__49227;
    wire N__49226;
    wire N__49223;
    wire N__49220;
    wire N__49217;
    wire N__49214;
    wire N__49211;
    wire N__49208;
    wire N__49203;
    wire N__49200;
    wire N__49197;
    wire N__49194;
    wire N__49191;
    wire N__49188;
    wire N__49187;
    wire N__49184;
    wire N__49181;
    wire N__49178;
    wire N__49175;
    wire N__49172;
    wire N__49169;
    wire N__49166;
    wire N__49163;
    wire N__49160;
    wire N__49157;
    wire N__49152;
    wire N__49149;
    wire N__49146;
    wire N__49145;
    wire N__49144;
    wire N__49143;
    wire N__49142;
    wire N__49141;
    wire N__49138;
    wire N__49133;
    wire N__49130;
    wire N__49127;
    wire N__49124;
    wire N__49123;
    wire N__49120;
    wire N__49113;
    wire N__49110;
    wire N__49107;
    wire N__49102;
    wire N__49095;
    wire N__49092;
    wire N__49091;
    wire N__49088;
    wire N__49085;
    wire N__49082;
    wire N__49079;
    wire N__49076;
    wire N__49073;
    wire N__49068;
    wire N__49065;
    wire N__49062;
    wire N__49059;
    wire N__49056;
    wire N__49053;
    wire N__49050;
    wire N__49049;
    wire N__49048;
    wire N__49045;
    wire N__49044;
    wire N__49043;
    wire N__49042;
    wire N__49041;
    wire N__49040;
    wire N__49037;
    wire N__49034;
    wire N__49033;
    wire N__49032;
    wire N__49031;
    wire N__49030;
    wire N__49021;
    wire N__49018;
    wire N__49017;
    wire N__49016;
    wire N__49015;
    wire N__49014;
    wire N__49011;
    wire N__49008;
    wire N__49005;
    wire N__49004;
    wire N__49003;
    wire N__49002;
    wire N__49001;
    wire N__49000;
    wire N__48999;
    wire N__48998;
    wire N__48997;
    wire N__48996;
    wire N__48995;
    wire N__48994;
    wire N__48993;
    wire N__48992;
    wire N__48989;
    wire N__48986;
    wire N__48985;
    wire N__48984;
    wire N__48979;
    wire N__48976;
    wire N__48973;
    wire N__48970;
    wire N__48969;
    wire N__48968;
    wire N__48967;
    wire N__48964;
    wire N__48961;
    wire N__48956;
    wire N__48955;
    wire N__48950;
    wire N__48947;
    wire N__48940;
    wire N__48937;
    wire N__48928;
    wire N__48925;
    wire N__48922;
    wire N__48921;
    wire N__48920;
    wire N__48919;
    wire N__48914;
    wire N__48913;
    wire N__48910;
    wire N__48907;
    wire N__48902;
    wire N__48895;
    wire N__48894;
    wire N__48891;
    wire N__48884;
    wire N__48877;
    wire N__48874;
    wire N__48869;
    wire N__48862;
    wire N__48859;
    wire N__48854;
    wire N__48849;
    wire N__48846;
    wire N__48845;
    wire N__48844;
    wire N__48843;
    wire N__48842;
    wire N__48839;
    wire N__48836;
    wire N__48829;
    wire N__48826;
    wire N__48819;
    wire N__48810;
    wire N__48803;
    wire N__48794;
    wire N__48787;
    wire N__48774;
    wire N__48773;
    wire N__48770;
    wire N__48767;
    wire N__48764;
    wire N__48761;
    wire N__48756;
    wire N__48753;
    wire N__48750;
    wire N__48747;
    wire N__48746;
    wire N__48743;
    wire N__48740;
    wire N__48737;
    wire N__48734;
    wire N__48731;
    wire N__48728;
    wire N__48723;
    wire N__48720;
    wire N__48717;
    wire N__48714;
    wire N__48711;
    wire N__48708;
    wire N__48705;
    wire N__48702;
    wire N__48701;
    wire N__48700;
    wire N__48699;
    wire N__48698;
    wire N__48697;
    wire N__48696;
    wire N__48695;
    wire N__48692;
    wire N__48691;
    wire N__48686;
    wire N__48683;
    wire N__48682;
    wire N__48681;
    wire N__48680;
    wire N__48677;
    wire N__48672;
    wire N__48671;
    wire N__48670;
    wire N__48667;
    wire N__48666;
    wire N__48663;
    wire N__48660;
    wire N__48657;
    wire N__48654;
    wire N__48651;
    wire N__48648;
    wire N__48647;
    wire N__48646;
    wire N__48645;
    wire N__48642;
    wire N__48637;
    wire N__48628;
    wire N__48625;
    wire N__48620;
    wire N__48613;
    wire N__48610;
    wire N__48607;
    wire N__48604;
    wire N__48597;
    wire N__48594;
    wire N__48589;
    wire N__48576;
    wire N__48573;
    wire N__48572;
    wire N__48569;
    wire N__48566;
    wire N__48563;
    wire N__48560;
    wire N__48559;
    wire N__48554;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48537;
    wire N__48534;
    wire N__48531;
    wire N__48528;
    wire N__48527;
    wire N__48526;
    wire N__48523;
    wire N__48520;
    wire N__48519;
    wire N__48516;
    wire N__48513;
    wire N__48510;
    wire N__48507;
    wire N__48498;
    wire N__48495;
    wire N__48492;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48482;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48474;
    wire N__48471;
    wire N__48468;
    wire N__48465;
    wire N__48462;
    wire N__48453;
    wire N__48452;
    wire N__48451;
    wire N__48450;
    wire N__48449;
    wire N__48448;
    wire N__48447;
    wire N__48446;
    wire N__48445;
    wire N__48444;
    wire N__48443;
    wire N__48442;
    wire N__48441;
    wire N__48440;
    wire N__48439;
    wire N__48438;
    wire N__48437;
    wire N__48436;
    wire N__48435;
    wire N__48434;
    wire N__48433;
    wire N__48432;
    wire N__48431;
    wire N__48430;
    wire N__48429;
    wire N__48428;
    wire N__48427;
    wire N__48426;
    wire N__48425;
    wire N__48424;
    wire N__48423;
    wire N__48422;
    wire N__48421;
    wire N__48420;
    wire N__48419;
    wire N__48418;
    wire N__48417;
    wire N__48416;
    wire N__48415;
    wire N__48414;
    wire N__48413;
    wire N__48412;
    wire N__48411;
    wire N__48410;
    wire N__48409;
    wire N__48408;
    wire N__48407;
    wire N__48406;
    wire N__48405;
    wire N__48404;
    wire N__48403;
    wire N__48402;
    wire N__48401;
    wire N__48400;
    wire N__48399;
    wire N__48398;
    wire N__48397;
    wire N__48396;
    wire N__48395;
    wire N__48394;
    wire N__48393;
    wire N__48392;
    wire N__48391;
    wire N__48390;
    wire N__48389;
    wire N__48388;
    wire N__48387;
    wire N__48386;
    wire N__48385;
    wire N__48384;
    wire N__48383;
    wire N__48240;
    wire N__48237;
    wire N__48234;
    wire N__48233;
    wire N__48230;
    wire N__48227;
    wire N__48222;
    wire N__48219;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48204;
    wire N__48201;
    wire N__48198;
    wire N__48197;
    wire N__48194;
    wire N__48191;
    wire N__48188;
    wire N__48185;
    wire N__48182;
    wire N__48177;
    wire N__48176;
    wire N__48173;
    wire N__48170;
    wire N__48165;
    wire N__48162;
    wire N__48161;
    wire N__48158;
    wire N__48155;
    wire N__48150;
    wire N__48149;
    wire N__48148;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48137;
    wire N__48134;
    wire N__48133;
    wire N__48132;
    wire N__48129;
    wire N__48124;
    wire N__48121;
    wire N__48116;
    wire N__48113;
    wire N__48108;
    wire N__48103;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48087;
    wire N__48084;
    wire N__48081;
    wire N__48078;
    wire N__48077;
    wire N__48074;
    wire N__48073;
    wire N__48070;
    wire N__48067;
    wire N__48064;
    wire N__48061;
    wire N__48058;
    wire N__48055;
    wire N__48052;
    wire N__48045;
    wire N__48042;
    wire N__48039;
    wire N__48038;
    wire N__48035;
    wire N__48032;
    wire N__48029;
    wire N__48028;
    wire N__48025;
    wire N__48022;
    wire N__48019;
    wire N__48016;
    wire N__48009;
    wire N__48006;
    wire N__48003;
    wire N__48000;
    wire N__47997;
    wire N__47996;
    wire N__47995;
    wire N__47994;
    wire N__47993;
    wire N__47992;
    wire N__47991;
    wire N__47988;
    wire N__47985;
    wire N__47982;
    wire N__47981;
    wire N__47978;
    wire N__47975;
    wire N__47970;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47950;
    wire N__47945;
    wire N__47940;
    wire N__47935;
    wire N__47928;
    wire N__47927;
    wire N__47924;
    wire N__47921;
    wire N__47918;
    wire N__47915;
    wire N__47912;
    wire N__47909;
    wire N__47906;
    wire N__47903;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47891;
    wire N__47886;
    wire N__47883;
    wire N__47882;
    wire N__47879;
    wire N__47876;
    wire N__47873;
    wire N__47870;
    wire N__47869;
    wire N__47866;
    wire N__47863;
    wire N__47860;
    wire N__47857;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47843;
    wire N__47840;
    wire N__47839;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47827;
    wire N__47820;
    wire N__47817;
    wire N__47814;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47802;
    wire N__47799;
    wire N__47798;
    wire N__47797;
    wire N__47796;
    wire N__47795;
    wire N__47792;
    wire N__47789;
    wire N__47784;
    wire N__47781;
    wire N__47780;
    wire N__47779;
    wire N__47778;
    wire N__47775;
    wire N__47770;
    wire N__47767;
    wire N__47760;
    wire N__47757;
    wire N__47754;
    wire N__47749;
    wire N__47742;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47732;
    wire N__47727;
    wire N__47724;
    wire N__47721;
    wire N__47718;
    wire N__47715;
    wire N__47712;
    wire N__47711;
    wire N__47708;
    wire N__47707;
    wire N__47704;
    wire N__47701;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47685;
    wire N__47682;
    wire N__47679;
    wire N__47678;
    wire N__47675;
    wire N__47672;
    wire N__47669;
    wire N__47664;
    wire N__47661;
    wire N__47658;
    wire N__47655;
    wire N__47654;
    wire N__47651;
    wire N__47648;
    wire N__47643;
    wire N__47640;
    wire N__47637;
    wire N__47634;
    wire N__47631;
    wire N__47630;
    wire N__47627;
    wire N__47624;
    wire N__47621;
    wire N__47618;
    wire N__47617;
    wire N__47612;
    wire N__47609;
    wire N__47604;
    wire N__47601;
    wire N__47598;
    wire N__47597;
    wire N__47594;
    wire N__47591;
    wire N__47586;
    wire N__47583;
    wire N__47582;
    wire N__47579;
    wire N__47576;
    wire N__47571;
    wire N__47570;
    wire N__47567;
    wire N__47564;
    wire N__47561;
    wire N__47556;
    wire N__47553;
    wire N__47550;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47538;
    wire N__47535;
    wire N__47534;
    wire N__47531;
    wire N__47530;
    wire N__47529;
    wire N__47528;
    wire N__47527;
    wire N__47526;
    wire N__47525;
    wire N__47524;
    wire N__47523;
    wire N__47520;
    wire N__47519;
    wire N__47518;
    wire N__47515;
    wire N__47512;
    wire N__47507;
    wire N__47506;
    wire N__47505;
    wire N__47504;
    wire N__47503;
    wire N__47502;
    wire N__47501;
    wire N__47498;
    wire N__47497;
    wire N__47496;
    wire N__47495;
    wire N__47494;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47477;
    wire N__47476;
    wire N__47473;
    wire N__47468;
    wire N__47465;
    wire N__47462;
    wire N__47459;
    wire N__47458;
    wire N__47455;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47437;
    wire N__47432;
    wire N__47423;
    wire N__47422;
    wire N__47419;
    wire N__47416;
    wire N__47409;
    wire N__47406;
    wire N__47403;
    wire N__47398;
    wire N__47395;
    wire N__47390;
    wire N__47385;
    wire N__47382;
    wire N__47379;
    wire N__47374;
    wire N__47369;
    wire N__47366;
    wire N__47359;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47328;
    wire N__47325;
    wire N__47324;
    wire N__47323;
    wire N__47320;
    wire N__47317;
    wire N__47314;
    wire N__47311;
    wire N__47308;
    wire N__47305;
    wire N__47298;
    wire N__47295;
    wire N__47294;
    wire N__47291;
    wire N__47290;
    wire N__47287;
    wire N__47284;
    wire N__47281;
    wire N__47278;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47264;
    wire N__47263;
    wire N__47260;
    wire N__47255;
    wire N__47252;
    wire N__47249;
    wire N__47246;
    wire N__47241;
    wire N__47238;
    wire N__47237;
    wire N__47236;
    wire N__47235;
    wire N__47232;
    wire N__47231;
    wire N__47230;
    wire N__47229;
    wire N__47226;
    wire N__47225;
    wire N__47220;
    wire N__47217;
    wire N__47212;
    wire N__47209;
    wire N__47206;
    wire N__47203;
    wire N__47200;
    wire N__47197;
    wire N__47194;
    wire N__47181;
    wire N__47180;
    wire N__47177;
    wire N__47176;
    wire N__47173;
    wire N__47172;
    wire N__47169;
    wire N__47168;
    wire N__47165;
    wire N__47164;
    wire N__47163;
    wire N__47160;
    wire N__47157;
    wire N__47156;
    wire N__47153;
    wire N__47148;
    wire N__47143;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47129;
    wire N__47126;
    wire N__47115;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47105;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47088;
    wire N__47085;
    wire N__47084;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47066;
    wire N__47063;
    wire N__47060;
    wire N__47057;
    wire N__47054;
    wire N__47051;
    wire N__47048;
    wire N__47043;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47028;
    wire N__47025;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47015;
    wire N__47012;
    wire N__47009;
    wire N__47006;
    wire N__47003;
    wire N__46998;
    wire N__46995;
    wire N__46992;
    wire N__46989;
    wire N__46986;
    wire N__46983;
    wire N__46980;
    wire N__46979;
    wire N__46978;
    wire N__46977;
    wire N__46974;
    wire N__46971;
    wire N__46970;
    wire N__46969;
    wire N__46966;
    wire N__46965;
    wire N__46964;
    wire N__46963;
    wire N__46960;
    wire N__46959;
    wire N__46958;
    wire N__46955;
    wire N__46950;
    wire N__46945;
    wire N__46944;
    wire N__46943;
    wire N__46942;
    wire N__46941;
    wire N__46940;
    wire N__46937;
    wire N__46932;
    wire N__46931;
    wire N__46930;
    wire N__46929;
    wire N__46928;
    wire N__46927;
    wire N__46924;
    wire N__46923;
    wire N__46920;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46908;
    wire N__46905;
    wire N__46898;
    wire N__46895;
    wire N__46890;
    wire N__46887;
    wire N__46886;
    wire N__46883;
    wire N__46882;
    wire N__46879;
    wire N__46878;
    wire N__46875;
    wire N__46872;
    wire N__46871;
    wire N__46868;
    wire N__46865;
    wire N__46862;
    wire N__46859;
    wire N__46856;
    wire N__46853;
    wire N__46850;
    wire N__46841;
    wire N__46826;
    wire N__46821;
    wire N__46818;
    wire N__46807;
    wire N__46804;
    wire N__46801;
    wire N__46788;
    wire N__46787;
    wire N__46786;
    wire N__46783;
    wire N__46778;
    wire N__46777;
    wire N__46776;
    wire N__46775;
    wire N__46774;
    wire N__46769;
    wire N__46766;
    wire N__46763;
    wire N__46758;
    wire N__46755;
    wire N__46746;
    wire N__46745;
    wire N__46744;
    wire N__46743;
    wire N__46740;
    wire N__46737;
    wire N__46734;
    wire N__46729;
    wire N__46726;
    wire N__46723;
    wire N__46722;
    wire N__46719;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46705;
    wire N__46702;
    wire N__46695;
    wire N__46692;
    wire N__46689;
    wire N__46688;
    wire N__46687;
    wire N__46684;
    wire N__46683;
    wire N__46680;
    wire N__46679;
    wire N__46678;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46670;
    wire N__46669;
    wire N__46666;
    wire N__46663;
    wire N__46658;
    wire N__46657;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46643;
    wire N__46642;
    wire N__46639;
    wire N__46634;
    wire N__46631;
    wire N__46626;
    wire N__46621;
    wire N__46618;
    wire N__46613;
    wire N__46602;
    wire N__46599;
    wire N__46596;
    wire N__46593;
    wire N__46592;
    wire N__46589;
    wire N__46586;
    wire N__46581;
    wire N__46580;
    wire N__46579;
    wire N__46578;
    wire N__46571;
    wire N__46570;
    wire N__46569;
    wire N__46568;
    wire N__46567;
    wire N__46564;
    wire N__46561;
    wire N__46552;
    wire N__46549;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46535;
    wire N__46534;
    wire N__46531;
    wire N__46530;
    wire N__46529;
    wire N__46528;
    wire N__46525;
    wire N__46524;
    wire N__46523;
    wire N__46520;
    wire N__46519;
    wire N__46518;
    wire N__46517;
    wire N__46516;
    wire N__46515;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46495;
    wire N__46492;
    wire N__46489;
    wire N__46488;
    wire N__46487;
    wire N__46484;
    wire N__46483;
    wire N__46482;
    wire N__46481;
    wire N__46476;
    wire N__46475;
    wire N__46472;
    wire N__46467;
    wire N__46464;
    wire N__46457;
    wire N__46452;
    wire N__46451;
    wire N__46450;
    wire N__46449;
    wire N__46448;
    wire N__46445;
    wire N__46442;
    wire N__46439;
    wire N__46436;
    wire N__46431;
    wire N__46428;
    wire N__46425;
    wire N__46422;
    wire N__46417;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46401;
    wire N__46396;
    wire N__46393;
    wire N__46384;
    wire N__46381;
    wire N__46376;
    wire N__46371;
    wire N__46356;
    wire N__46353;
    wire N__46352;
    wire N__46349;
    wire N__46346;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46317;
    wire N__46314;
    wire N__46311;
    wire N__46308;
    wire N__46305;
    wire N__46302;
    wire N__46299;
    wire N__46296;
    wire N__46293;
    wire N__46290;
    wire N__46287;
    wire N__46284;
    wire N__46281;
    wire N__46278;
    wire N__46275;
    wire N__46274;
    wire N__46273;
    wire N__46268;
    wire N__46265;
    wire N__46260;
    wire N__46257;
    wire N__46256;
    wire N__46255;
    wire N__46250;
    wire N__46247;
    wire N__46242;
    wire N__46239;
    wire N__46238;
    wire N__46235;
    wire N__46234;
    wire N__46229;
    wire N__46226;
    wire N__46221;
    wire N__46218;
    wire N__46217;
    wire N__46216;
    wire N__46211;
    wire N__46208;
    wire N__46203;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46107;
    wire N__46104;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46068;
    wire N__46065;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46046;
    wire N__46043;
    wire N__46040;
    wire N__46039;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46007;
    wire N__46004;
    wire N__46001;
    wire N__45998;
    wire N__45995;
    wire N__45990;
    wire N__45987;
    wire N__45984;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45972;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45939;
    wire N__45938;
    wire N__45935;
    wire N__45934;
    wire N__45931;
    wire N__45928;
    wire N__45925;
    wire N__45918;
    wire N__45915;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45891;
    wire N__45890;
    wire N__45887;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45877;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45855;
    wire N__45852;
    wire N__45849;
    wire N__45848;
    wire N__45845;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45833;
    wire N__45828;
    wire N__45825;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45806;
    wire N__45805;
    wire N__45802;
    wire N__45799;
    wire N__45796;
    wire N__45793;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45764;
    wire N__45763;
    wire N__45762;
    wire N__45761;
    wire N__45760;
    wire N__45759;
    wire N__45758;
    wire N__45757;
    wire N__45756;
    wire N__45755;
    wire N__45754;
    wire N__45753;
    wire N__45752;
    wire N__45751;
    wire N__45750;
    wire N__45749;
    wire N__45748;
    wire N__45747;
    wire N__45746;
    wire N__45745;
    wire N__45744;
    wire N__45743;
    wire N__45742;
    wire N__45741;
    wire N__45740;
    wire N__45739;
    wire N__45738;
    wire N__45737;
    wire N__45734;
    wire N__45733;
    wire N__45732;
    wire N__45731;
    wire N__45730;
    wire N__45729;
    wire N__45728;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45720;
    wire N__45717;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45704;
    wire N__45701;
    wire N__45700;
    wire N__45699;
    wire N__45698;
    wire N__45697;
    wire N__45696;
    wire N__45695;
    wire N__45694;
    wire N__45693;
    wire N__45692;
    wire N__45691;
    wire N__45690;
    wire N__45689;
    wire N__45688;
    wire N__45687;
    wire N__45686;
    wire N__45685;
    wire N__45684;
    wire N__45681;
    wire N__45680;
    wire N__45679;
    wire N__45678;
    wire N__45677;
    wire N__45676;
    wire N__45673;
    wire N__45672;
    wire N__45671;
    wire N__45670;
    wire N__45667;
    wire N__45666;
    wire N__45665;
    wire N__45662;
    wire N__45661;
    wire N__45660;
    wire N__45659;
    wire N__45658;
    wire N__45657;
    wire N__45656;
    wire N__45655;
    wire N__45654;
    wire N__45651;
    wire N__45650;
    wire N__45649;
    wire N__45648;
    wire N__45647;
    wire N__45646;
    wire N__45645;
    wire N__45644;
    wire N__45643;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45635;
    wire N__45634;
    wire N__45633;
    wire N__45632;
    wire N__45631;
    wire N__45630;
    wire N__45629;
    wire N__45628;
    wire N__45627;
    wire N__45626;
    wire N__45625;
    wire N__45616;
    wire N__45607;
    wire N__45600;
    wire N__45591;
    wire N__45590;
    wire N__45589;
    wire N__45588;
    wire N__45587;
    wire N__45586;
    wire N__45585;
    wire N__45584;
    wire N__45581;
    wire N__45580;
    wire N__45579;
    wire N__45578;
    wire N__45577;
    wire N__45576;
    wire N__45573;
    wire N__45572;
    wire N__45571;
    wire N__45570;
    wire N__45569;
    wire N__45568;
    wire N__45567;
    wire N__45566;
    wire N__45565;
    wire N__45564;
    wire N__45563;
    wire N__45562;
    wire N__45559;
    wire N__45558;
    wire N__45557;
    wire N__45556;
    wire N__45555;
    wire N__45554;
    wire N__45553;
    wire N__45552;
    wire N__45551;
    wire N__45550;
    wire N__45549;
    wire N__45548;
    wire N__45547;
    wire N__45544;
    wire N__45543;
    wire N__45542;
    wire N__45541;
    wire N__45540;
    wire N__45539;
    wire N__45536;
    wire N__45535;
    wire N__45534;
    wire N__45533;
    wire N__45532;
    wire N__45531;
    wire N__45530;
    wire N__45527;
    wire N__45526;
    wire N__45525;
    wire N__45514;
    wire N__45507;
    wire N__45506;
    wire N__45505;
    wire N__45504;
    wire N__45503;
    wire N__45502;
    wire N__45501;
    wire N__45498;
    wire N__45497;
    wire N__45496;
    wire N__45493;
    wire N__45486;
    wire N__45479;
    wire N__45470;
    wire N__45463;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45452;
    wire N__45451;
    wire N__45450;
    wire N__45449;
    wire N__45448;
    wire N__45447;
    wire N__45446;
    wire N__45445;
    wire N__45444;
    wire N__45443;
    wire N__45442;
    wire N__45441;
    wire N__45440;
    wire N__45439;
    wire N__45438;
    wire N__45437;
    wire N__45436;
    wire N__45435;
    wire N__45434;
    wire N__45433;
    wire N__45432;
    wire N__45423;
    wire N__45418;
    wire N__45417;
    wire N__45416;
    wire N__45415;
    wire N__45414;
    wire N__45413;
    wire N__45412;
    wire N__45411;
    wire N__45402;
    wire N__45401;
    wire N__45400;
    wire N__45399;
    wire N__45396;
    wire N__45395;
    wire N__45394;
    wire N__45393;
    wire N__45392;
    wire N__45391;
    wire N__45386;
    wire N__45375;
    wire N__45368;
    wire N__45357;
    wire N__45348;
    wire N__45339;
    wire N__45338;
    wire N__45333;
    wire N__45326;
    wire N__45325;
    wire N__45324;
    wire N__45323;
    wire N__45322;
    wire N__45319;
    wire N__45318;
    wire N__45317;
    wire N__45314;
    wire N__45313;
    wire N__45312;
    wire N__45311;
    wire N__45310;
    wire N__45309;
    wire N__45308;
    wire N__45307;
    wire N__45304;
    wire N__45303;
    wire N__45302;
    wire N__45299;
    wire N__45298;
    wire N__45297;
    wire N__45296;
    wire N__45293;
    wire N__45292;
    wire N__45289;
    wire N__45286;
    wire N__45285;
    wire N__45284;
    wire N__45283;
    wire N__45282;
    wire N__45281;
    wire N__45280;
    wire N__45279;
    wire N__45276;
    wire N__45269;
    wire N__45262;
    wire N__45251;
    wire N__45244;
    wire N__45239;
    wire N__45232;
    wire N__45231;
    wire N__45228;
    wire N__45227;
    wire N__45224;
    wire N__45223;
    wire N__45220;
    wire N__45219;
    wire N__45218;
    wire N__45211;
    wire N__45206;
    wire N__45197;
    wire N__45190;
    wire N__45183;
    wire N__45174;
    wire N__45163;
    wire N__45152;
    wire N__45145;
    wire N__45142;
    wire N__45141;
    wire N__45140;
    wire N__45139;
    wire N__45138;
    wire N__45137;
    wire N__45136;
    wire N__45135;
    wire N__45134;
    wire N__45131;
    wire N__45128;
    wire N__45123;
    wire N__45116;
    wire N__45105;
    wire N__45104;
    wire N__45101;
    wire N__45100;
    wire N__45099;
    wire N__45098;
    wire N__45097;
    wire N__45096;
    wire N__45095;
    wire N__45094;
    wire N__45093;
    wire N__45092;
    wire N__45091;
    wire N__45090;
    wire N__45087;
    wire N__45082;
    wire N__45079;
    wire N__45074;
    wire N__45067;
    wire N__45060;
    wire N__45053;
    wire N__45046;
    wire N__45037;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45029;
    wire N__45028;
    wire N__45027;
    wire N__45026;
    wire N__45025;
    wire N__45024;
    wire N__45023;
    wire N__45020;
    wire N__45019;
    wire N__45018;
    wire N__45017;
    wire N__45016;
    wire N__45007;
    wire N__45004;
    wire N__44999;
    wire N__44990;
    wire N__44983;
    wire N__44980;
    wire N__44973;
    wire N__44962;
    wire N__44959;
    wire N__44958;
    wire N__44957;
    wire N__44956;
    wire N__44955;
    wire N__44950;
    wire N__44941;
    wire N__44938;
    wire N__44937;
    wire N__44936;
    wire N__44935;
    wire N__44934;
    wire N__44933;
    wire N__44932;
    wire N__44931;
    wire N__44930;
    wire N__44929;
    wire N__44928;
    wire N__44927;
    wire N__44926;
    wire N__44925;
    wire N__44924;
    wire N__44923;
    wire N__44918;
    wire N__44907;
    wire N__44900;
    wire N__44893;
    wire N__44886;
    wire N__44879;
    wire N__44872;
    wire N__44871;
    wire N__44870;
    wire N__44869;
    wire N__44864;
    wire N__44863;
    wire N__44862;
    wire N__44861;
    wire N__44860;
    wire N__44859;
    wire N__44856;
    wire N__44849;
    wire N__44844;
    wire N__44835;
    wire N__44834;
    wire N__44833;
    wire N__44832;
    wire N__44829;
    wire N__44828;
    wire N__44823;
    wire N__44812;
    wire N__44805;
    wire N__44794;
    wire N__44791;
    wire N__44774;
    wire N__44771;
    wire N__44762;
    wire N__44753;
    wire N__44748;
    wire N__44743;
    wire N__44740;
    wire N__44737;
    wire N__44730;
    wire N__44723;
    wire N__44722;
    wire N__44719;
    wire N__44718;
    wire N__44717;
    wire N__44716;
    wire N__44715;
    wire N__44714;
    wire N__44711;
    wire N__44710;
    wire N__44707;
    wire N__44706;
    wire N__44699;
    wire N__44692;
    wire N__44685;
    wire N__44678;
    wire N__44671;
    wire N__44670;
    wire N__44667;
    wire N__44666;
    wire N__44665;
    wire N__44656;
    wire N__44649;
    wire N__44646;
    wire N__44645;
    wire N__44644;
    wire N__44637;
    wire N__44636;
    wire N__44635;
    wire N__44634;
    wire N__44633;
    wire N__44632;
    wire N__44631;
    wire N__44630;
    wire N__44625;
    wire N__44618;
    wire N__44611;
    wire N__44602;
    wire N__44601;
    wire N__44600;
    wire N__44597;
    wire N__44596;
    wire N__44589;
    wire N__44582;
    wire N__44575;
    wire N__44568;
    wire N__44561;
    wire N__44554;
    wire N__44547;
    wire N__44538;
    wire N__44531;
    wire N__44528;
    wire N__44523;
    wire N__44522;
    wire N__44521;
    wire N__44520;
    wire N__44519;
    wire N__44518;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44500;
    wire N__44495;
    wire N__44492;
    wire N__44487;
    wire N__44486;
    wire N__44485;
    wire N__44484;
    wire N__44483;
    wire N__44474;
    wire N__44463;
    wire N__44450;
    wire N__44441;
    wire N__44440;
    wire N__44437;
    wire N__44436;
    wire N__44435;
    wire N__44434;
    wire N__44433;
    wire N__44426;
    wire N__44419;
    wire N__44416;
    wire N__44407;
    wire N__44398;
    wire N__44393;
    wire N__44386;
    wire N__44385;
    wire N__44382;
    wire N__44375;
    wire N__44368;
    wire N__44365;
    wire N__44360;
    wire N__44355;
    wire N__44346;
    wire N__44339;
    wire N__44332;
    wire N__44325;
    wire N__44320;
    wire N__44313;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44291;
    wire N__44288;
    wire N__44281;
    wire N__44272;
    wire N__44265;
    wire N__44258;
    wire N__44251;
    wire N__44248;
    wire N__44245;
    wire N__44240;
    wire N__44237;
    wire N__44228;
    wire N__44221;
    wire N__44208;
    wire N__44203;
    wire N__44196;
    wire N__44189;
    wire N__44186;
    wire N__44183;
    wire N__44176;
    wire N__44173;
    wire N__44168;
    wire N__44161;
    wire N__44148;
    wire N__44147;
    wire N__44144;
    wire N__44141;
    wire N__44138;
    wire N__44135;
    wire N__44130;
    wire N__44129;
    wire N__44128;
    wire N__44127;
    wire N__44124;
    wire N__44123;
    wire N__44122;
    wire N__44119;
    wire N__44118;
    wire N__44117;
    wire N__44116;
    wire N__44115;
    wire N__44114;
    wire N__44113;
    wire N__44110;
    wire N__44109;
    wire N__44106;
    wire N__44103;
    wire N__44100;
    wire N__44099;
    wire N__44098;
    wire N__44091;
    wire N__44090;
    wire N__44087;
    wire N__44086;
    wire N__44083;
    wire N__44082;
    wire N__44081;
    wire N__44070;
    wire N__44067;
    wire N__44064;
    wire N__44061;
    wire N__44058;
    wire N__44055;
    wire N__44052;
    wire N__44045;
    wire N__44038;
    wire N__44035;
    wire N__44026;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43997;
    wire N__43992;
    wire N__43989;
    wire N__43986;
    wire N__43985;
    wire N__43982;
    wire N__43979;
    wire N__43976;
    wire N__43975;
    wire N__43972;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43956;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43940;
    wire N__43937;
    wire N__43936;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43917;
    wire N__43914;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43898;
    wire N__43895;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43860;
    wire N__43857;
    wire N__43854;
    wire N__43853;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43843;
    wire N__43840;
    wire N__43833;
    wire N__43830;
    wire N__43827;
    wire N__43824;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43811;
    wire N__43810;
    wire N__43807;
    wire N__43804;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43785;
    wire N__43782;
    wire N__43779;
    wire N__43776;
    wire N__43773;
    wire N__43770;
    wire N__43767;
    wire N__43766;
    wire N__43763;
    wire N__43760;
    wire N__43757;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43743;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43733;
    wire N__43730;
    wire N__43727;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43695;
    wire N__43692;
    wire N__43689;
    wire N__43688;
    wire N__43685;
    wire N__43682;
    wire N__43679;
    wire N__43676;
    wire N__43671;
    wire N__43668;
    wire N__43667;
    wire N__43664;
    wire N__43663;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43648;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43616;
    wire N__43615;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43599;
    wire N__43596;
    wire N__43595;
    wire N__43592;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43572;
    wire N__43571;
    wire N__43568;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43548;
    wire N__43545;
    wire N__43540;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43500;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43490;
    wire N__43487;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43477;
    wire N__43470;
    wire N__43467;
    wire N__43464;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43451;
    wire N__43448;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43425;
    wire N__43422;
    wire N__43419;
    wire N__43416;
    wire N__43413;
    wire N__43410;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43399;
    wire N__43396;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43380;
    wire N__43377;
    wire N__43374;
    wire N__43371;
    wire N__43370;
    wire N__43369;
    wire N__43366;
    wire N__43361;
    wire N__43358;
    wire N__43353;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43335;
    wire N__43332;
    wire N__43329;
    wire N__43326;
    wire N__43323;
    wire N__43320;
    wire N__43319;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43304;
    wire N__43299;
    wire N__43296;
    wire N__43295;
    wire N__43294;
    wire N__43293;
    wire N__43290;
    wire N__43289;
    wire N__43286;
    wire N__43283;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43269;
    wire N__43266;
    wire N__43259;
    wire N__43256;
    wire N__43251;
    wire N__43250;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43232;
    wire N__43229;
    wire N__43228;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43200;
    wire N__43199;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43175;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43160;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43137;
    wire N__43132;
    wire N__43125;
    wire N__43122;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43110;
    wire N__43107;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43089;
    wire N__43086;
    wire N__43085;
    wire N__43084;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43068;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43052;
    wire N__43049;
    wire N__43048;
    wire N__43045;
    wire N__43042;
    wire N__43039;
    wire N__43036;
    wire N__43029;
    wire N__43026;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43008;
    wire N__43005;
    wire N__43002;
    wire N__42999;
    wire N__42998;
    wire N__42995;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42983;
    wire N__42978;
    wire N__42975;
    wire N__42974;
    wire N__42973;
    wire N__42972;
    wire N__42969;
    wire N__42966;
    wire N__42963;
    wire N__42960;
    wire N__42955;
    wire N__42948;
    wire N__42947;
    wire N__42942;
    wire N__42939;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42906;
    wire N__42903;
    wire N__42900;
    wire N__42899;
    wire N__42898;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42880;
    wire N__42877;
    wire N__42872;
    wire N__42867;
    wire N__42864;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42844;
    wire N__42841;
    wire N__42838;
    wire N__42831;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42807;
    wire N__42804;
    wire N__42801;
    wire N__42800;
    wire N__42797;
    wire N__42794;
    wire N__42791;
    wire N__42788;
    wire N__42785;
    wire N__42782;
    wire N__42779;
    wire N__42776;
    wire N__42771;
    wire N__42768;
    wire N__42767;
    wire N__42766;
    wire N__42765;
    wire N__42762;
    wire N__42759;
    wire N__42756;
    wire N__42753;
    wire N__42750;
    wire N__42747;
    wire N__42742;
    wire N__42735;
    wire N__42732;
    wire N__42729;
    wire N__42726;
    wire N__42725;
    wire N__42722;
    wire N__42719;
    wire N__42716;
    wire N__42715;
    wire N__42712;
    wire N__42709;
    wire N__42706;
    wire N__42703;
    wire N__42702;
    wire N__42701;
    wire N__42696;
    wire N__42693;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42676;
    wire N__42673;
    wire N__42666;
    wire N__42665;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42641;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42633;
    wire N__42630;
    wire N__42627;
    wire N__42626;
    wire N__42625;
    wire N__42622;
    wire N__42619;
    wire N__42614;
    wire N__42611;
    wire N__42610;
    wire N__42609;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42594;
    wire N__42589;
    wire N__42576;
    wire N__42575;
    wire N__42572;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42542;
    wire N__42539;
    wire N__42538;
    wire N__42535;
    wire N__42532;
    wire N__42529;
    wire N__42526;
    wire N__42519;
    wire N__42518;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42494;
    wire N__42491;
    wire N__42488;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42455;
    wire N__42454;
    wire N__42451;
    wire N__42448;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42426;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42401;
    wire N__42400;
    wire N__42397;
    wire N__42392;
    wire N__42387;
    wire N__42386;
    wire N__42383;
    wire N__42380;
    wire N__42377;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42326;
    wire N__42325;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42275;
    wire N__42270;
    wire N__42267;
    wire N__42264;
    wire N__42263;
    wire N__42262;
    wire N__42261;
    wire N__42260;
    wire N__42257;
    wire N__42256;
    wire N__42253;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42241;
    wire N__42236;
    wire N__42233;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42213;
    wire N__42210;
    wire N__42209;
    wire N__42208;
    wire N__42205;
    wire N__42202;
    wire N__42199;
    wire N__42194;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42170;
    wire N__42169;
    wire N__42164;
    wire N__42161;
    wire N__42156;
    wire N__42153;
    wire N__42150;
    wire N__42147;
    wire N__42144;
    wire N__42141;
    wire N__42138;
    wire N__42135;
    wire N__42132;
    wire N__42129;
    wire N__42128;
    wire N__42125;
    wire N__42124;
    wire N__42121;
    wire N__42118;
    wire N__42115;
    wire N__42110;
    wire N__42107;
    wire N__42104;
    wire N__42099;
    wire N__42096;
    wire N__42093;
    wire N__42090;
    wire N__42089;
    wire N__42086;
    wire N__42083;
    wire N__42080;
    wire N__42077;
    wire N__42076;
    wire N__42071;
    wire N__42068;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42056;
    wire N__42053;
    wire N__42052;
    wire N__42049;
    wire N__42046;
    wire N__42043;
    wire N__42040;
    wire N__42035;
    wire N__42030;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42020;
    wire N__42017;
    wire N__42014;
    wire N__42013;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__41999;
    wire N__41996;
    wire N__41991;
    wire N__41990;
    wire N__41989;
    wire N__41988;
    wire N__41985;
    wire N__41982;
    wire N__41981;
    wire N__41978;
    wire N__41977;
    wire N__41976;
    wire N__41975;
    wire N__41974;
    wire N__41973;
    wire N__41972;
    wire N__41969;
    wire N__41958;
    wire N__41957;
    wire N__41954;
    wire N__41953;
    wire N__41950;
    wire N__41949;
    wire N__41948;
    wire N__41945;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41933;
    wire N__41932;
    wire N__41929;
    wire N__41928;
    wire N__41923;
    wire N__41920;
    wire N__41913;
    wire N__41910;
    wire N__41905;
    wire N__41896;
    wire N__41883;
    wire N__41882;
    wire N__41881;
    wire N__41878;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41857;
    wire N__41852;
    wire N__41847;
    wire N__41844;
    wire N__41843;
    wire N__41840;
    wire N__41837;
    wire N__41834;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41804;
    wire N__41801;
    wire N__41798;
    wire N__41795;
    wire N__41790;
    wire N__41787;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41765;
    wire N__41764;
    wire N__41761;
    wire N__41756;
    wire N__41753;
    wire N__41748;
    wire N__41745;
    wire N__41742;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41723;
    wire N__41722;
    wire N__41719;
    wire N__41714;
    wire N__41711;
    wire N__41708;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41673;
    wire N__41670;
    wire N__41669;
    wire N__41666;
    wire N__41665;
    wire N__41664;
    wire N__41663;
    wire N__41662;
    wire N__41661;
    wire N__41660;
    wire N__41657;
    wire N__41654;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41644;
    wire N__41641;
    wire N__41640;
    wire N__41637;
    wire N__41636;
    wire N__41635;
    wire N__41632;
    wire N__41631;
    wire N__41626;
    wire N__41613;
    wire N__41612;
    wire N__41611;
    wire N__41604;
    wire N__41601;
    wire N__41600;
    wire N__41599;
    wire N__41598;
    wire N__41595;
    wire N__41594;
    wire N__41593;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41577;
    wire N__41574;
    wire N__41567;
    wire N__41564;
    wire N__41561;
    wire N__41558;
    wire N__41541;
    wire N__41538;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41528;
    wire N__41525;
    wire N__41522;
    wire N__41519;
    wire N__41514;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41492;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41477;
    wire N__41474;
    wire N__41473;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41459;
    wire N__41456;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41436;
    wire N__41433;
    wire N__41430;
    wire N__41427;
    wire N__41424;
    wire N__41423;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41366;
    wire N__41363;
    wire N__41362;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41346;
    wire N__41343;
    wire N__41340;
    wire N__41337;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41280;
    wire N__41279;
    wire N__41276;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41247;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41204;
    wire N__41203;
    wire N__41200;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41173;
    wire N__41170;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41154;
    wire N__41153;
    wire N__41150;
    wire N__41147;
    wire N__41146;
    wire N__41143;
    wire N__41140;
    wire N__41137;
    wire N__41132;
    wire N__41129;
    wire N__41124;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41108;
    wire N__41105;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41060;
    wire N__41059;
    wire N__41056;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41044;
    wire N__41041;
    wire N__41036;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__40998;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40986;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40956;
    wire N__40953;
    wire N__40952;
    wire N__40947;
    wire N__40944;
    wire N__40941;
    wire N__40938;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40928;
    wire N__40923;
    wire N__40920;
    wire N__40917;
    wire N__40914;
    wire N__40911;
    wire N__40908;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40893;
    wire N__40890;
    wire N__40889;
    wire N__40888;
    wire N__40887;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40852;
    wire N__40849;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40813;
    wire N__40812;
    wire N__40807;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40797;
    wire N__40794;
    wire N__40789;
    wire N__40784;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40757;
    wire N__40756;
    wire N__40755;
    wire N__40750;
    wire N__40747;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40734;
    wire N__40729;
    wire N__40726;
    wire N__40719;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40691;
    wire N__40688;
    wire N__40685;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40657;
    wire N__40656;
    wire N__40655;
    wire N__40652;
    wire N__40649;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40614;
    wire N__40611;
    wire N__40610;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40583;
    wire N__40580;
    wire N__40577;
    wire N__40572;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40560;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40544;
    wire N__40541;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40529;
    wire N__40526;
    wire N__40521;
    wire N__40518;
    wire N__40517;
    wire N__40514;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40502;
    wire N__40499;
    wire N__40494;
    wire N__40491;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40478;
    wire N__40475;
    wire N__40472;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40454;
    wire N__40449;
    wire N__40448;
    wire N__40445;
    wire N__40444;
    wire N__40443;
    wire N__40442;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40432;
    wire N__40429;
    wire N__40426;
    wire N__40423;
    wire N__40420;
    wire N__40417;
    wire N__40404;
    wire N__40401;
    wire N__40398;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40386;
    wire N__40383;
    wire N__40380;
    wire N__40377;
    wire N__40376;
    wire N__40373;
    wire N__40370;
    wire N__40365;
    wire N__40362;
    wire N__40361;
    wire N__40358;
    wire N__40355;
    wire N__40354;
    wire N__40353;
    wire N__40352;
    wire N__40351;
    wire N__40348;
    wire N__40347;
    wire N__40346;
    wire N__40343;
    wire N__40338;
    wire N__40335;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40314;
    wire N__40311;
    wire N__40296;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40277;
    wire N__40274;
    wire N__40273;
    wire N__40270;
    wire N__40267;
    wire N__40264;
    wire N__40261;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40230;
    wire N__40229;
    wire N__40228;
    wire N__40225;
    wire N__40222;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40190;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40180;
    wire N__40177;
    wire N__40172;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40152;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40106;
    wire N__40103;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40090;
    wire N__40085;
    wire N__40082;
    wire N__40077;
    wire N__40074;
    wire N__40071;
    wire N__40068;
    wire N__40065;
    wire N__40062;
    wire N__40059;
    wire N__40058;
    wire N__40057;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40045;
    wire N__40042;
    wire N__40035;
    wire N__40032;
    wire N__40029;
    wire N__40026;
    wire N__40023;
    wire N__40022;
    wire N__40019;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40004;
    wire N__39999;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39983;
    wire N__39982;
    wire N__39979;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39950;
    wire N__39949;
    wire N__39946;
    wire N__39941;
    wire N__39938;
    wire N__39933;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39911;
    wire N__39910;
    wire N__39907;
    wire N__39904;
    wire N__39901;
    wire N__39896;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39857;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39847;
    wire N__39846;
    wire N__39843;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39828;
    wire N__39825;
    wire N__39820;
    wire N__39817;
    wire N__39814;
    wire N__39811;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39795;
    wire N__39794;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39784;
    wire N__39779;
    wire N__39778;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39760;
    wire N__39757;
    wire N__39752;
    wire N__39749;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39729;
    wire N__39728;
    wire N__39725;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39705;
    wire N__39702;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39686;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39670;
    wire N__39663;
    wire N__39660;
    wire N__39659;
    wire N__39656;
    wire N__39653;
    wire N__39650;
    wire N__39647;
    wire N__39642;
    wire N__39639;
    wire N__39638;
    wire N__39637;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39606;
    wire N__39603;
    wire N__39600;
    wire N__39597;
    wire N__39594;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39586;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39570;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39552;
    wire N__39549;
    wire N__39548;
    wire N__39545;
    wire N__39544;
    wire N__39541;
    wire N__39540;
    wire N__39539;
    wire N__39538;
    wire N__39537;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39526;
    wire N__39525;
    wire N__39524;
    wire N__39523;
    wire N__39520;
    wire N__39519;
    wire N__39518;
    wire N__39517;
    wire N__39514;
    wire N__39513;
    wire N__39510;
    wire N__39509;
    wire N__39508;
    wire N__39507;
    wire N__39504;
    wire N__39503;
    wire N__39500;
    wire N__39499;
    wire N__39496;
    wire N__39491;
    wire N__39488;
    wire N__39483;
    wire N__39474;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39448;
    wire N__39443;
    wire N__39440;
    wire N__39423;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39412;
    wire N__39409;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39395;
    wire N__39392;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39380;
    wire N__39377;
    wire N__39376;
    wire N__39373;
    wire N__39370;
    wire N__39367;
    wire N__39364;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39341;
    wire N__39338;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39320;
    wire N__39317;
    wire N__39316;
    wire N__39313;
    wire N__39310;
    wire N__39307;
    wire N__39304;
    wire N__39297;
    wire N__39296;
    wire N__39293;
    wire N__39292;
    wire N__39289;
    wire N__39286;
    wire N__39283;
    wire N__39280;
    wire N__39273;
    wire N__39272;
    wire N__39269;
    wire N__39268;
    wire N__39265;
    wire N__39262;
    wire N__39259;
    wire N__39256;
    wire N__39249;
    wire N__39248;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39194;
    wire N__39191;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39176;
    wire N__39173;
    wire N__39170;
    wire N__39167;
    wire N__39164;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39125;
    wire N__39122;
    wire N__39119;
    wire N__39116;
    wire N__39113;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39075;
    wire N__39072;
    wire N__39069;
    wire N__39066;
    wire N__39063;
    wire N__39062;
    wire N__39057;
    wire N__39054;
    wire N__39053;
    wire N__39050;
    wire N__39047;
    wire N__39042;
    wire N__39041;
    wire N__39038;
    wire N__39035;
    wire N__39030;
    wire N__39027;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39015;
    wire N__39012;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38993;
    wire N__38990;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38927;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38910;
    wire N__38907;
    wire N__38906;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38889;
    wire N__38888;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38874;
    wire N__38871;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38859;
    wire N__38856;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38846;
    wire N__38841;
    wire N__38838;
    wire N__38837;
    wire N__38834;
    wire N__38831;
    wire N__38826;
    wire N__38823;
    wire N__38822;
    wire N__38819;
    wire N__38816;
    wire N__38811;
    wire N__38808;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38796;
    wire N__38793;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38781;
    wire N__38778;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38763;
    wire N__38760;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38748;
    wire N__38745;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38733;
    wire N__38730;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38708;
    wire N__38705;
    wire N__38702;
    wire N__38699;
    wire N__38694;
    wire N__38691;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38669;
    wire N__38666;
    wire N__38663;
    wire N__38660;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38648;
    wire N__38645;
    wire N__38642;
    wire N__38639;
    wire N__38634;
    wire N__38631;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38616;
    wire N__38613;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38601;
    wire N__38598;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38586;
    wire N__38583;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38571;
    wire N__38568;
    wire N__38567;
    wire N__38564;
    wire N__38561;
    wire N__38556;
    wire N__38553;
    wire N__38552;
    wire N__38549;
    wire N__38546;
    wire N__38541;
    wire N__38538;
    wire N__38537;
    wire N__38534;
    wire N__38531;
    wire N__38526;
    wire N__38523;
    wire N__38522;
    wire N__38519;
    wire N__38516;
    wire N__38513;
    wire N__38508;
    wire N__38505;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38493;
    wire N__38490;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38446;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38434;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38396;
    wire N__38393;
    wire N__38390;
    wire N__38387;
    wire N__38382;
    wire N__38379;
    wire N__38378;
    wire N__38375;
    wire N__38372;
    wire N__38367;
    wire N__38364;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38337;
    wire N__38334;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38315;
    wire N__38312;
    wire N__38309;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38284;
    wire N__38279;
    wire N__38276;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38259;
    wire N__38256;
    wire N__38253;
    wire N__38252;
    wire N__38249;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38232;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38204;
    wire N__38199;
    wire N__38196;
    wire N__38193;
    wire N__38190;
    wire N__38187;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38172;
    wire N__38169;
    wire N__38168;
    wire N__38165;
    wire N__38162;
    wire N__38159;
    wire N__38156;
    wire N__38153;
    wire N__38150;
    wire N__38145;
    wire N__38142;
    wire N__38139;
    wire N__38136;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38121;
    wire N__38120;
    wire N__38115;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38102;
    wire N__38097;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38066;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38039;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38022;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38003;
    wire N__38000;
    wire N__37997;
    wire N__37994;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37973;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37892;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37859;
    wire N__37854;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37820;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37793;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37764;
    wire N__37761;
    wire N__37758;
    wire N__37755;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37745;
    wire N__37744;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37701;
    wire N__37698;
    wire N__37695;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37681;
    wire N__37676;
    wire N__37673;
    wire N__37668;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37646;
    wire N__37641;
    wire N__37638;
    wire N__37635;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37616;
    wire N__37615;
    wire N__37612;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37587;
    wire N__37584;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37544;
    wire N__37541;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37521;
    wire N__37518;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37502;
    wire N__37499;
    wire N__37494;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37482;
    wire N__37481;
    wire N__37480;
    wire N__37477;
    wire N__37474;
    wire N__37471;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37446;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37423;
    wire N__37420;
    wire N__37417;
    wire N__37416;
    wire N__37413;
    wire N__37408;
    wire N__37405;
    wire N__37402;
    wire N__37399;
    wire N__37396;
    wire N__37395;
    wire N__37390;
    wire N__37387;
    wire N__37384;
    wire N__37381;
    wire N__37378;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37317;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37305;
    wire N__37302;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37294;
    wire N__37289;
    wire N__37286;
    wire N__37281;
    wire N__37278;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37270;
    wire N__37265;
    wire N__37262;
    wire N__37257;
    wire N__37256;
    wire N__37255;
    wire N__37254;
    wire N__37253;
    wire N__37252;
    wire N__37251;
    wire N__37250;
    wire N__37249;
    wire N__37248;
    wire N__37247;
    wire N__37246;
    wire N__37245;
    wire N__37244;
    wire N__37243;
    wire N__37242;
    wire N__37239;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37178;
    wire N__37169;
    wire N__37162;
    wire N__37155;
    wire N__37152;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37098;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37086;
    wire N__37083;
    wire N__37082;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37065;
    wire N__37062;
    wire N__37061;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37044;
    wire N__37041;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37027;
    wire N__37022;
    wire N__37019;
    wire N__37014;
    wire N__37011;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36976;
    wire N__36971;
    wire N__36968;
    wire N__36963;
    wire N__36960;
    wire N__36957;
    wire N__36956;
    wire N__36953;
    wire N__36950;
    wire N__36945;
    wire N__36942;
    wire N__36941;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36910;
    wire N__36905;
    wire N__36902;
    wire N__36901;
    wire N__36896;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36881;
    wire N__36876;
    wire N__36873;
    wire N__36870;
    wire N__36869;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36849;
    wire N__36848;
    wire N__36845;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36831;
    wire N__36828;
    wire N__36827;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36817;
    wire N__36810;
    wire N__36807;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36795;
    wire N__36792;
    wire N__36791;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36774;
    wire N__36771;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36738;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36713;
    wire N__36712;
    wire N__36709;
    wire N__36706;
    wire N__36703;
    wire N__36700;
    wire N__36697;
    wire N__36690;
    wire N__36687;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36677;
    wire N__36676;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36657;
    wire N__36656;
    wire N__36653;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36641;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36629;
    wire N__36626;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36609;
    wire N__36606;
    wire N__36605;
    wire N__36602;
    wire N__36601;
    wire N__36600;
    wire N__36597;
    wire N__36596;
    wire N__36595;
    wire N__36594;
    wire N__36593;
    wire N__36592;
    wire N__36591;
    wire N__36590;
    wire N__36587;
    wire N__36586;
    wire N__36583;
    wire N__36576;
    wire N__36575;
    wire N__36570;
    wire N__36569;
    wire N__36566;
    wire N__36565;
    wire N__36564;
    wire N__36561;
    wire N__36560;
    wire N__36557;
    wire N__36556;
    wire N__36555;
    wire N__36554;
    wire N__36551;
    wire N__36550;
    wire N__36549;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36528;
    wire N__36523;
    wire N__36508;
    wire N__36499;
    wire N__36494;
    wire N__36477;
    wire N__36474;
    wire N__36471;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36458;
    wire N__36457;
    wire N__36454;
    wire N__36449;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36427;
    wire N__36424;
    wire N__36421;
    wire N__36418;
    wire N__36411;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36403;
    wire N__36400;
    wire N__36397;
    wire N__36394;
    wire N__36387;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36369;
    wire N__36366;
    wire N__36365;
    wire N__36362;
    wire N__36361;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36335;
    wire N__36332;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36302;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36263;
    wire N__36260;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36240;
    wire N__36237;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36209;
    wire N__36208;
    wire N__36207;
    wire N__36206;
    wire N__36203;
    wire N__36200;
    wire N__36199;
    wire N__36198;
    wire N__36197;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36193;
    wire N__36192;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36176;
    wire N__36173;
    wire N__36172;
    wire N__36171;
    wire N__36170;
    wire N__36167;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36159;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36144;
    wire N__36141;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36121;
    wire N__36114;
    wire N__36099;
    wire N__36094;
    wire N__36081;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36048;
    wire N__36047;
    wire N__36044;
    wire N__36043;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36008;
    wire N__36005;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35989;
    wire N__35982;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35951;
    wire N__35948;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35928;
    wire N__35925;
    wire N__35924;
    wire N__35921;
    wire N__35918;
    wire N__35915;
    wire N__35912;
    wire N__35907;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35887;
    wire N__35882;
    wire N__35881;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35853;
    wire N__35850;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35835;
    wire N__35832;
    wire N__35829;
    wire N__35826;
    wire N__35825;
    wire N__35822;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35812;
    wire N__35809;
    wire N__35802;
    wire N__35801;
    wire N__35800;
    wire N__35797;
    wire N__35796;
    wire N__35795;
    wire N__35794;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35784;
    wire N__35783;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35772;
    wire N__35769;
    wire N__35768;
    wire N__35761;
    wire N__35758;
    wire N__35755;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35737;
    wire N__35736;
    wire N__35735;
    wire N__35734;
    wire N__35733;
    wire N__35726;
    wire N__35725;
    wire N__35724;
    wire N__35723;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35704;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35679;
    wire N__35676;
    wire N__35671;
    wire N__35670;
    wire N__35669;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35657;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35636;
    wire N__35633;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35603;
    wire N__35598;
    wire N__35595;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35575;
    wire N__35572;
    wire N__35569;
    wire N__35566;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35548;
    wire N__35545;
    wire N__35538;
    wire N__35535;
    wire N__35526;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35504;
    wire N__35503;
    wire N__35502;
    wire N__35499;
    wire N__35494;
    wire N__35491;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35475;
    wire N__35472;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35460;
    wire N__35457;
    wire N__35454;
    wire N__35451;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35425;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35411;
    wire N__35408;
    wire N__35403;
    wire N__35400;
    wire N__35397;
    wire N__35394;
    wire N__35393;
    wire N__35392;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35373;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35361;
    wire N__35358;
    wire N__35357;
    wire N__35356;
    wire N__35353;
    wire N__35348;
    wire N__35343;
    wire N__35340;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35301;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35283;
    wire N__35280;
    wire N__35279;
    wire N__35278;
    wire N__35275;
    wire N__35272;
    wire N__35269;
    wire N__35262;
    wire N__35259;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35249;
    wire N__35246;
    wire N__35243;
    wire N__35242;
    wire N__35239;
    wire N__35234;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35150;
    wire N__35149;
    wire N__35148;
    wire N__35147;
    wire N__35146;
    wire N__35145;
    wire N__35142;
    wire N__35137;
    wire N__35134;
    wire N__35129;
    wire N__35128;
    wire N__35127;
    wire N__35126;
    wire N__35125;
    wire N__35122;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35108;
    wire N__35107;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35084;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35016;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35006;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34982;
    wire N__34977;
    wire N__34976;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34952;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34916;
    wire N__34913;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34868;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34815;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34787;
    wire N__34784;
    wire N__34781;
    wire N__34780;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34742;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34723;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34691;
    wire N__34688;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34667;
    wire N__34662;
    wire N__34659;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34645;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34613;
    wire N__34612;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34598;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34577;
    wire N__34574;
    wire N__34571;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34554;
    wire N__34551;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34518;
    wire N__34517;
    wire N__34516;
    wire N__34515;
    wire N__34512;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34504;
    wire N__34501;
    wire N__34500;
    wire N__34499;
    wire N__34496;
    wire N__34491;
    wire N__34488;
    wire N__34483;
    wire N__34482;
    wire N__34481;
    wire N__34480;
    wire N__34477;
    wire N__34476;
    wire N__34473;
    wire N__34468;
    wire N__34463;
    wire N__34458;
    wire N__34455;
    wire N__34450;
    wire N__34437;
    wire N__34434;
    wire N__34433;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34375;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34289;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34276;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34257;
    wire N__34254;
    wire N__34251;
    wire N__34248;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34232;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34205;
    wire N__34200;
    wire N__34197;
    wire N__34196;
    wire N__34195;
    wire N__34194;
    wire N__34193;
    wire N__34192;
    wire N__34191;
    wire N__34190;
    wire N__34189;
    wire N__34186;
    wire N__34185;
    wire N__34184;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34172;
    wire N__34169;
    wire N__34168;
    wire N__34165;
    wire N__34164;
    wire N__34161;
    wire N__34160;
    wire N__34159;
    wire N__34156;
    wire N__34143;
    wire N__34138;
    wire N__34131;
    wire N__34124;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34076;
    wire N__34075;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34065;
    wire N__34064;
    wire N__34061;
    wire N__34054;
    wire N__34051;
    wire N__34046;
    wire N__34041;
    wire N__34040;
    wire N__34039;
    wire N__34036;
    wire N__34031;
    wire N__34028;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34016;
    wire N__34015;
    wire N__34012;
    wire N__34009;
    wire N__34004;
    wire N__34001;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33885;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33873;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33857;
    wire N__33854;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33830;
    wire N__33827;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33312;
    wire N__33309;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33275;
    wire N__33274;
    wire N__33273;
    wire N__33272;
    wire N__33271;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33263;
    wire N__33262;
    wire N__33259;
    wire N__33256;
    wire N__33255;
    wire N__33252;
    wire N__33251;
    wire N__33246;
    wire N__33243;
    wire N__33236;
    wire N__33231;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33207;
    wire N__33204;
    wire N__33203;
    wire N__33200;
    wire N__33197;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33177;
    wire N__33176;
    wire N__33173;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33153;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33066;
    wire N__33063;
    wire N__33062;
    wire N__33059;
    wire N__33056;
    wire N__33053;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33020;
    wire N__33017;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32903;
    wire N__32902;
    wire N__32901;
    wire N__32900;
    wire N__32899;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32893;
    wire N__32888;
    wire N__32887;
    wire N__32884;
    wire N__32883;
    wire N__32882;
    wire N__32879;
    wire N__32878;
    wire N__32875;
    wire N__32874;
    wire N__32867;
    wire N__32862;
    wire N__32859;
    wire N__32854;
    wire N__32851;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32823;
    wire N__32820;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32812;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32793;
    wire N__32792;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32782;
    wire N__32777;
    wire N__32774;
    wire N__32769;
    wire N__32766;
    wire N__32765;
    wire N__32764;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32746;
    wire N__32745;
    wire N__32740;
    wire N__32737;
    wire N__32734;
    wire N__32731;
    wire N__32728;
    wire N__32721;
    wire N__32718;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32710;
    wire N__32709;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32694;
    wire N__32689;
    wire N__32682;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32666;
    wire N__32663;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32648;
    wire N__32643;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32624;
    wire N__32623;
    wire N__32620;
    wire N__32615;
    wire N__32612;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32589;
    wire N__32588;
    wire N__32587;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32568;
    wire N__32565;
    wire N__32562;
    wire N__32559;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32530;
    wire N__32527;
    wire N__32524;
    wire N__32521;
    wire N__32516;
    wire N__32511;
    wire N__32508;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32486;
    wire N__32483;
    wire N__32480;
    wire N__32477;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32449;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32430;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32422;
    wire N__32417;
    wire N__32414;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32387;
    wire N__32384;
    wire N__32381;
    wire N__32380;
    wire N__32375;
    wire N__32372;
    wire N__32367;
    wire N__32364;
    wire N__32363;
    wire N__32360;
    wire N__32357;
    wire N__32356;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32337;
    wire N__32334;
    wire N__32333;
    wire N__32332;
    wire N__32329;
    wire N__32324;
    wire N__32321;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32304;
    wire N__32301;
    wire N__32298;
    wire N__32295;
    wire N__32292;
    wire N__32291;
    wire N__32288;
    wire N__32287;
    wire N__32284;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32250;
    wire N__32247;
    wire N__32246;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32182;
    wire N__32179;
    wire N__32176;
    wire N__32173;
    wire N__32170;
    wire N__32167;
    wire N__32164;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32077;
    wire N__32074;
    wire N__32071;
    wire N__32066;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32048;
    wire N__32045;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31972;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31913;
    wire N__31910;
    wire N__31907;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31877;
    wire N__31876;
    wire N__31875;
    wire N__31874;
    wire N__31871;
    wire N__31868;
    wire N__31867;
    wire N__31866;
    wire N__31865;
    wire N__31864;
    wire N__31863;
    wire N__31860;
    wire N__31859;
    wire N__31858;
    wire N__31855;
    wire N__31854;
    wire N__31853;
    wire N__31852;
    wire N__31851;
    wire N__31848;
    wire N__31845;
    wire N__31840;
    wire N__31839;
    wire N__31838;
    wire N__31837;
    wire N__31836;
    wire N__31835;
    wire N__31834;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31826;
    wire N__31823;
    wire N__31822;
    wire N__31819;
    wire N__31814;
    wire N__31807;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31784;
    wire N__31775;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31749;
    wire N__31734;
    wire N__31733;
    wire N__31732;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31692;
    wire N__31689;
    wire N__31688;
    wire N__31685;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31668;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31632;
    wire N__31629;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31611;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31599;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31585;
    wire N__31580;
    wire N__31577;
    wire N__31572;
    wire N__31569;
    wire N__31568;
    wire N__31565;
    wire N__31564;
    wire N__31561;
    wire N__31558;
    wire N__31555;
    wire N__31552;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31538;
    wire N__31537;
    wire N__31534;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31460;
    wire N__31455;
    wire N__31454;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31441;
    wire N__31438;
    wire N__31435;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31388;
    wire N__31387;
    wire N__31384;
    wire N__31379;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31361;
    wire N__31360;
    wire N__31357;
    wire N__31354;
    wire N__31351;
    wire N__31346;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31316;
    wire N__31313;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31295;
    wire N__31290;
    wire N__31287;
    wire N__31286;
    wire N__31283;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31214;
    wire N__31213;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31187;
    wire N__31186;
    wire N__31183;
    wire N__31178;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31160;
    wire N__31157;
    wire N__31156;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31144;
    wire N__31141;
    wire N__31138;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31074;
    wire N__31071;
    wire N__31070;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31058;
    wire N__31055;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31017;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31005;
    wire N__31004;
    wire N__31003;
    wire N__31000;
    wire N__30999;
    wire N__30996;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30977;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30914;
    wire N__30911;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30845;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30837;
    wire N__30836;
    wire N__30833;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30785;
    wire N__30784;
    wire N__30783;
    wire N__30782;
    wire N__30781;
    wire N__30780;
    wire N__30779;
    wire N__30778;
    wire N__30777;
    wire N__30776;
    wire N__30775;
    wire N__30774;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30722;
    wire N__30713;
    wire N__30706;
    wire N__30699;
    wire N__30690;
    wire N__30687;
    wire N__30686;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30666;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30658;
    wire N__30653;
    wire N__30650;
    wire N__30645;
    wire N__30644;
    wire N__30643;
    wire N__30640;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30628;
    wire N__30627;
    wire N__30626;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30609;
    wire N__30606;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30572;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30552;
    wire N__30549;
    wire N__30548;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30518;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30446;
    wire N__30443;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30414;
    wire N__30411;
    wire N__30410;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30330;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30306;
    wire N__30305;
    wire N__30304;
    wire N__30303;
    wire N__30302;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30294;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30286;
    wire N__30285;
    wire N__30284;
    wire N__30283;
    wire N__30278;
    wire N__30277;
    wire N__30276;
    wire N__30275;
    wire N__30274;
    wire N__30263;
    wire N__30258;
    wire N__30257;
    wire N__30256;
    wire N__30255;
    wire N__30252;
    wire N__30251;
    wire N__30250;
    wire N__30247;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30227;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30211;
    wire N__30206;
    wire N__30197;
    wire N__30194;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30167;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30130;
    wire N__30125;
    wire N__30122;
    wire N__30117;
    wire N__30116;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30108;
    wire N__30105;
    wire N__30100;
    wire N__30097;
    wire N__30096;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30066;
    wire N__30063;
    wire N__30062;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30045;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30027;
    wire N__30024;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30012;
    wire N__30009;
    wire N__30008;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29939;
    wire N__29934;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29904;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29849;
    wire N__29846;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29828;
    wire N__29827;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29809;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29791;
    wire N__29788;
    wire N__29781;
    wire N__29778;
    wire N__29777;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29715;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29652;
    wire N__29651;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29632;
    wire N__29627;
    wire N__29624;
    wire N__29619;
    wire N__29618;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29586;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29574;
    wire N__29571;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29474;
    wire N__29471;
    wire N__29470;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29451;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29443;
    wire N__29438;
    wire N__29435;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29412;
    wire N__29409;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29397;
    wire N__29396;
    wire N__29395;
    wire N__29392;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29370;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29276;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29171;
    wire N__29168;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29158;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29105;
    wire N__29102;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29082;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29069;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29033;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28977;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28969;
    wire N__28966;
    wire N__28961;
    wire N__28958;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28916;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28901;
    wire N__28898;
    wire N__28897;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28878;
    wire N__28877;
    wire N__28876;
    wire N__28875;
    wire N__28874;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28866;
    wire N__28865;
    wire N__28864;
    wire N__28863;
    wire N__28862;
    wire N__28859;
    wire N__28858;
    wire N__28857;
    wire N__28856;
    wire N__28855;
    wire N__28852;
    wire N__28851;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28843;
    wire N__28842;
    wire N__28841;
    wire N__28840;
    wire N__28839;
    wire N__28838;
    wire N__28837;
    wire N__28836;
    wire N__28835;
    wire N__28834;
    wire N__28833;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28815;
    wire N__28812;
    wire N__28807;
    wire N__28802;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28786;
    wire N__28783;
    wire N__28778;
    wire N__28777;
    wire N__28776;
    wire N__28775;
    wire N__28774;
    wire N__28769;
    wire N__28764;
    wire N__28757;
    wire N__28750;
    wire N__28745;
    wire N__28742;
    wire N__28735;
    wire N__28732;
    wire N__28725;
    wire N__28722;
    wire N__28717;
    wire N__28714;
    wire N__28709;
    wire N__28704;
    wire N__28701;
    wire N__28692;
    wire N__28677;
    wire N__28674;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28647;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28613;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28587;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28548;
    wire N__28545;
    wire N__28544;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28475;
    wire N__28474;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28433;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28418;
    wire N__28415;
    wire N__28410;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28397;
    wire N__28394;
    wire N__28393;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28355;
    wire N__28352;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28247;
    wire N__28244;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28208;
    wire N__28207;
    wire N__28204;
    wire N__28203;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28188;
    wire N__28187;
    wire N__28186;
    wire N__28183;
    wire N__28182;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28162;
    wire N__28157;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28070;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28056;
    wire N__28053;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28032;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27972;
    wire N__27971;
    wire N__27968;
    wire N__27963;
    wire N__27960;
    wire N__27957;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27942;
    wire N__27939;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27873;
    wire N__27872;
    wire N__27871;
    wire N__27866;
    wire N__27863;
    wire N__27860;
    wire N__27855;
    wire N__27854;
    wire N__27853;
    wire N__27850;
    wire N__27845;
    wire N__27842;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27825;
    wire N__27824;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27816;
    wire N__27815;
    wire N__27812;
    wire N__27803;
    wire N__27798;
    wire N__27795;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27783;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27750;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27737;
    wire N__27736;
    wire N__27733;
    wire N__27732;
    wire N__27729;
    wire N__27728;
    wire N__27725;
    wire N__27724;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27704;
    wire N__27701;
    wire N__27690;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27682;
    wire N__27679;
    wire N__27678;
    wire N__27675;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27667;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27655;
    wire N__27652;
    wire N__27647;
    wire N__27636;
    wire N__27635;
    wire N__27632;
    wire N__27631;
    wire N__27628;
    wire N__27627;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27542;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27464;
    wire N__27463;
    wire N__27460;
    wire N__27459;
    wire N__27458;
    wire N__27457;
    wire N__27456;
    wire N__27453;
    wire N__27452;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27441;
    wire N__27440;
    wire N__27439;
    wire N__27438;
    wire N__27437;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27423;
    wire N__27422;
    wire N__27421;
    wire N__27420;
    wire N__27419;
    wire N__27416;
    wire N__27415;
    wire N__27412;
    wire N__27407;
    wire N__27402;
    wire N__27401;
    wire N__27400;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27389;
    wire N__27388;
    wire N__27387;
    wire N__27384;
    wire N__27377;
    wire N__27372;
    wire N__27363;
    wire N__27360;
    wire N__27355;
    wire N__27350;
    wire N__27339;
    wire N__27332;
    wire N__27329;
    wire N__27312;
    wire N__27311;
    wire N__27308;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27293;
    wire N__27290;
    wire N__27285;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27271;
    wire N__27266;
    wire N__27263;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27121;
    wire N__27116;
    wire N__27113;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27095;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27045;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26987;
    wire N__26986;
    wire N__26983;
    wire N__26978;
    wire N__26975;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26957;
    wire N__26954;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26939;
    wire N__26936;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26897;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26849;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26792;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26766;
    wire N__26765;
    wire N__26762;
    wire N__26761;
    wire N__26758;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26720;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26707;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26652;
    wire N__26651;
    wire N__26648;
    wire N__26647;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26629;
    wire N__26626;
    wire N__26621;
    wire N__26618;
    wire N__26613;
    wire N__26610;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26595;
    wire N__26592;
    wire N__26591;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26573;
    wire N__26572;
    wire N__26567;
    wire N__26564;
    wire N__26559;
    wire N__26558;
    wire N__26557;
    wire N__26554;
    wire N__26553;
    wire N__26552;
    wire N__26549;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26537;
    wire N__26532;
    wire N__26523;
    wire N__26522;
    wire N__26519;
    wire N__26518;
    wire N__26515;
    wire N__26510;
    wire N__26505;
    wire N__26504;
    wire N__26501;
    wire N__26500;
    wire N__26499;
    wire N__26498;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26482;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26439;
    wire N__26438;
    wire N__26437;
    wire N__26434;
    wire N__26433;
    wire N__26432;
    wire N__26429;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26413;
    wire N__26406;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26390;
    wire N__26389;
    wire N__26386;
    wire N__26381;
    wire N__26378;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26351;
    wire N__26348;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26332;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26316;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26301;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26258;
    wire N__26253;
    wire N__26250;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26235;
    wire N__26232;
    wire N__26231;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26223;
    wire N__26220;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26171;
    wire N__26170;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26136;
    wire N__26135;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26120;
    wire N__26119;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26106;
    wire N__26103;
    wire N__26100;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26048;
    wire N__26047;
    wire N__26046;
    wire N__26045;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26033;
    wire N__26028;
    wire N__26025;
    wire N__26016;
    wire N__26013;
    wire N__26012;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25931;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25916;
    wire N__25913;
    wire N__25908;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25896;
    wire N__25895;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25842;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25794;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25733;
    wire N__25730;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25492;
    wire N__25487;
    wire N__25484;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25372;
    wire N__25369;
    wire N__25366;
    wire N__25363;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25346;
    wire N__25343;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25258;
    wire N__25253;
    wire N__25250;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25197;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25149;
    wire N__25148;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25124;
    wire N__25121;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24971;
    wire N__24970;
    wire N__24969;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24946;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24902;
    wire N__24899;
    wire N__24898;
    wire N__24895;
    wire N__24890;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24872;
    wire N__24869;
    wire N__24868;
    wire N__24865;
    wire N__24862;
    wire N__24859;
    wire N__24856;
    wire N__24849;
    wire N__24846;
    wire N__24845;
    wire N__24844;
    wire N__24841;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24783;
    wire N__24780;
    wire N__24779;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24760;
    wire N__24757;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24734;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24653;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24636;
    wire N__24635;
    wire N__24632;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24603;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24590;
    wire N__24589;
    wire N__24588;
    wire N__24587;
    wire N__24586;
    wire N__24585;
    wire N__24582;
    wire N__24581;
    wire N__24580;
    wire N__24577;
    wire N__24572;
    wire N__24567;
    wire N__24558;
    wire N__24553;
    wire N__24546;
    wire N__24543;
    wire N__24542;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24534;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24513;
    wire N__24510;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24461;
    wire N__24460;
    wire N__24457;
    wire N__24456;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24444;
    wire N__24441;
    wire N__24436;
    wire N__24433;
    wire N__24428;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24374;
    wire N__24371;
    wire N__24370;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24345;
    wire N__24342;
    wire N__24335;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24281;
    wire N__24278;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24242;
    wire N__24241;
    wire N__24240;
    wire N__24239;
    wire N__24238;
    wire N__24237;
    wire N__24236;
    wire N__24235;
    wire N__24234;
    wire N__24231;
    wire N__24218;
    wire N__24215;
    wire N__24214;
    wire N__24213;
    wire N__24210;
    wire N__24209;
    wire N__24208;
    wire N__24207;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24190;
    wire N__24185;
    wire N__24182;
    wire N__24181;
    wire N__24178;
    wire N__24177;
    wire N__24176;
    wire N__24175;
    wire N__24174;
    wire N__24173;
    wire N__24172;
    wire N__24171;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24167;
    wire N__24164;
    wire N__24157;
    wire N__24152;
    wire N__24137;
    wire N__24132;
    wire N__24127;
    wire N__24120;
    wire N__24105;
    wire N__24102;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24034;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24004;
    wire N__23999;
    wire N__23996;
    wire N__23991;
    wire N__23990;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23979;
    wire N__23976;
    wire N__23971;
    wire N__23968;
    wire N__23963;
    wire N__23960;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23943;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23904;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23892;
    wire N__23889;
    wire N__23888;
    wire N__23887;
    wire N__23882;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23858;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23829;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23817;
    wire N__23814;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23777;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23695;
    wire N__23690;
    wire N__23687;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23600;
    wire N__23599;
    wire N__23596;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23577;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23471;
    wire N__23468;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23390;
    wire N__23387;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23319;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23283;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23247;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23214;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23168;
    wire N__23163;
    wire N__23160;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23143;
    wire N__23138;
    wire N__23135;
    wire N__23130;
    wire N__23127;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23075;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23054;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23030;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23010;
    wire N__23007;
    wire N__23006;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22970;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22943;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22923;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22898;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22877;
    wire N__22874;
    wire N__22871;
    wire N__22870;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22835;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22808;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22788;
    wire N__22785;
    wire N__22784;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22710;
    wire N__22707;
    wire N__22706;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22694;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22674;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22662;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22635;
    wire N__22632;
    wire N__22631;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22611;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22583;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22553;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22517;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22481;
    wire N__22476;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22425;
    wire N__22424;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22380;
    wire N__22379;
    wire N__22378;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22367;
    wire N__22366;
    wire N__22365;
    wire N__22364;
    wire N__22355;
    wire N__22350;
    wire N__22345;
    wire N__22342;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22085;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22031;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21941;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21743;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21710;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21675;
    wire N__21674;
    wire N__21671;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21656;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21533;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21481;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21440;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21337;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21281;
    wire N__21278;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21245;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21168;
    wire N__21167;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21138;
    wire N__21135;
    wire N__21134;
    wire N__21131;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21099;
    wire N__21096;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21082;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21066;
    wire N__21065;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21038;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21020;
    wire N__21017;
    wire N__21016;
    wire N__21013;
    wire N__21010;
    wire N__21007;
    wire N__21004;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20951;
    wire N__20948;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20933;
    wire N__20928;
    wire N__20925;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20910;
    wire N__20907;
    wire N__20906;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20850;
    wire N__20849;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20803;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20787;
    wire N__20786;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20624;
    wire N__20621;
    wire N__20616;
    wire N__20613;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20603;
    wire N__20598;
    wire N__20595;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20583;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20556;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20541;
    wire N__20538;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20426;
    wire N__20425;
    wire N__20424;
    wire N__20423;
    wire N__20420;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20412;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20394;
    wire N__20385;
    wire N__20382;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20336;
    wire N__20335;
    wire N__20332;
    wire N__20327;
    wire N__20324;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20222;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20209;
    wire N__20204;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20164;
    wire N__20163;
    wire N__20158;
    wire N__20153;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20138;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20102;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20003;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19966;
    wire N__19961;
    wire N__19958;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19916;
    wire N__19915;
    wire N__19912;
    wire N__19907;
    wire N__19904;
    wire N__19899;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19881;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19850;
    wire N__19847;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19823;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19728;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19694;
    wire N__19691;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19616;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19604;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19596;
    wire N__19595;
    wire N__19594;
    wire N__19587;
    wire N__19586;
    wire N__19583;
    wire N__19582;
    wire N__19581;
    wire N__19580;
    wire N__19575;
    wire N__19574;
    wire N__19571;
    wire N__19566;
    wire N__19565;
    wire N__19564;
    wire N__19561;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19545;
    wire N__19540;
    wire N__19527;
    wire N__19524;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19516;
    wire N__19515;
    wire N__19514;
    wire N__19513;
    wire N__19512;
    wire N__19511;
    wire N__19510;
    wire N__19505;
    wire N__19504;
    wire N__19501;
    wire N__19500;
    wire N__19497;
    wire N__19496;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19484;
    wire N__19481;
    wire N__19480;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19461;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19431;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19419;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19388;
    wire N__19387;
    wire N__19382;
    wire N__19379;
    wire N__19378;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19366;
    wire N__19363;
    wire N__19358;
    wire N__19353;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19341;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19313;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19287;
    wire N__19286;
    wire N__19283;
    wire N__19282;
    wire N__19281;
    wire N__19278;
    wire N__19273;
    wire N__19272;
    wire N__19271;
    wire N__19268;
    wire N__19267;
    wire N__19266;
    wire N__19265;
    wire N__19264;
    wire N__19263;
    wire N__19262;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19232;
    wire N__19227;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19174;
    wire N__19173;
    wire N__19170;
    wire N__19165;
    wire N__19162;
    wire N__19155;
    wire N__19154;
    wire N__19151;
    wire N__19150;
    wire N__19149;
    wire N__19146;
    wire N__19145;
    wire N__19144;
    wire N__19143;
    wire N__19142;
    wire N__19139;
    wire N__19134;
    wire N__19131;
    wire N__19126;
    wire N__19123;
    wire N__19122;
    wire N__19119;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19082;
    wire N__19077;
    wire N__19074;
    wire N__19073;
    wire N__19068;
    wire N__19065;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19050;
    wire N__19049;
    wire N__19044;
    wire N__19041;
    wire N__19038;
    wire N__19037;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18987;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18971;
    wire N__18968;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18815;
    wire N__18812;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18797;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18557;
    wire N__18552;
    wire N__18549;
    wire N__18548;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18521;
    wire N__18520;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18504;
    wire N__18503;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18489;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18474;
    wire N__18471;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18440;
    wire N__18435;
    wire N__18434;
    wire N__18433;
    wire N__18432;
    wire N__18429;
    wire N__18424;
    wire N__18421;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire NEOPXL_c;
    wire \nx.n13325_cascade_ ;
    wire \nx.n11535_cascade_ ;
    wire \nx.n11672_cascade_ ;
    wire \nx.n13326 ;
    wire \nx.n11692 ;
    wire \nx.n12204 ;
    wire \nx.n11696_cascade_ ;
    wire \nx.n7131_cascade_ ;
    wire \nx.n13263_cascade_ ;
    wire \nx.n7120_cascade_ ;
    wire \nx.n13262_cascade_ ;
    wire \nx.n3739 ;
    wire \nx.n3739_cascade_ ;
    wire \nx.n7120 ;
    wire \nx.n9700_cascade_ ;
    wire \nx.n7131 ;
    wire \nx.n12117_cascade_ ;
    wire n7239_cascade_;
    wire \nx.n9700 ;
    wire \nx.n9702 ;
    wire \nx.n11606 ;
    wire update_color;
    wire \nx.n10_adj_653 ;
    wire \nx.n13271 ;
    wire \nx.n12369_cascade_ ;
    wire neo_pixel_transmitter_t0_15;
    wire neo_pixel_transmitter_t0_8;
    wire \nx.n2908_cascade_ ;
    wire \nx.n3007_cascade_ ;
    wire \nx.n3106_cascade_ ;
    wire \nx.n19_adj_698 ;
    wire \nx.n3105_cascade_ ;
    wire \nx.n3100_cascade_ ;
    wire \nx.n29_adj_697_cascade_ ;
    wire \nx.n12331_cascade_ ;
    wire \nx.n12335 ;
    wire \nx.n37_adj_695_cascade_ ;
    wire \nx.n12333 ;
    wire \nx.n31_adj_691_cascade_ ;
    wire \nx.n49_adj_693_cascade_ ;
    wire \nx.n48_adj_692 ;
    wire \nx.n3116_cascade_ ;
    wire bfn_1_26_0_;
    wire \nx.n3176 ;
    wire \nx.n10888 ;
    wire \nx.n10889 ;
    wire \nx.n10890 ;
    wire \nx.n3106 ;
    wire \nx.n3173 ;
    wire \nx.n10891 ;
    wire \nx.n3105 ;
    wire \nx.n3172 ;
    wire \nx.n10892 ;
    wire \nx.n10893 ;
    wire \nx.n3170 ;
    wire \nx.n10894 ;
    wire \nx.n10895 ;
    wire \nx.n3102 ;
    wire \nx.n3169 ;
    wire bfn_1_27_0_;
    wire \nx.n10896 ;
    wire \nx.n3100 ;
    wire \nx.n3167 ;
    wire \nx.n10897 ;
    wire \nx.n10898 ;
    wire \nx.n10899 ;
    wire \nx.n10900 ;
    wire \nx.n3163 ;
    wire \nx.n10901 ;
    wire \nx.n10902 ;
    wire \nx.n10903 ;
    wire bfn_1_28_0_;
    wire \nx.n10904 ;
    wire \nx.n10905 ;
    wire \nx.n10906 ;
    wire \nx.n10907 ;
    wire \nx.n10908 ;
    wire \nx.n10909 ;
    wire \nx.n3154 ;
    wire \nx.n10910 ;
    wire \nx.n10911 ;
    wire \nx.n3153 ;
    wire bfn_1_29_0_;
    wire \nx.n3152 ;
    wire \nx.n10912 ;
    wire \nx.n10913 ;
    wire \nx.n10914 ;
    wire \nx.n10_adj_619_cascade_ ;
    wire \nx.n12_adj_621_cascade_ ;
    wire \nx.n1136_cascade_ ;
    wire \nx.n1203_cascade_ ;
    wire \nx.n1208_cascade_ ;
    wire bfn_1_31_0_;
    wire \nx.n10453 ;
    wire \nx.n10454 ;
    wire \nx.n10455 ;
    wire \nx.n10456 ;
    wire \nx.n10457 ;
    wire \nx.n10458 ;
    wire \nx.n10459 ;
    wire \nx.n10460 ;
    wire bfn_1_32_0_;
    wire \nx.n1203 ;
    wire \nx.n1270 ;
    wire \nx.n1302_cascade_ ;
    wire \nx.n1276 ;
    wire \nx.n1209 ;
    wire \nx.n1206_cascade_ ;
    wire \nx.n1273 ;
    wire \nx.n7 ;
    wire neo_pixel_transmitter_t0_23;
    wire neo_pixel_transmitter_t0_24;
    wire \nx.n7_adj_713_cascade_ ;
    wire \nx.n13491 ;
    wire \nx.n12933_cascade_ ;
    wire \nx.n12939 ;
    wire \nx.n10918 ;
    wire \nx.start ;
    wire \nx.n18_adj_711_cascade_ ;
    wire \nx.n20_adj_712 ;
    wire neo_pixel_transmitter_t0_6;
    wire neo_pixel_transmitter_t0_14;
    wire neo_pixel_transmitter_t0_5;
    wire neopxl_color_prev_5;
    wire n10_adj_776;
    wire neo_pixel_transmitter_t0_3;
    wire n12_adj_774;
    wire neo_pixel_transmitter_t0_12;
    wire \nx.neo_pixel_transmitter_done ;
    wire \nx.n11487_cascade_ ;
    wire \nx.n103 ;
    wire n9_adj_777;
    wire neopxl_color_prev_4;
    wire state_0_adj_727;
    wire state_1_adj_726;
    wire n7239;
    wire \nx.n7392 ;
    wire \nx.n13155 ;
    wire \nx.n13456_cascade_ ;
    wire \nx.n13156 ;
    wire \nx.n13459 ;
    wire \nx.n4_adj_642 ;
    wire neo_pixel_transmitter_t0_26;
    wire neo_pixel_transmitter_t0_16;
    wire \nx.color_bit_N_571_4 ;
    wire \nx.n13158 ;
    wire \nx.n59 ;
    wire \nx.n12371 ;
    wire \nx.n13042 ;
    wire \nx.n10947 ;
    wire \nx.n10947_cascade_ ;
    wire \nx.n10975 ;
    wire \nx.n3008_cascade_ ;
    wire \nx.n3096 ;
    wire \nx.n3096_cascade_ ;
    wire \nx.n47_adj_694 ;
    wire \nx.n45 ;
    wire \nx.n49_cascade_ ;
    wire \nx.n3017_cascade_ ;
    wire \nx.n3086 ;
    wire \nx.n3087 ;
    wire \nx.n3086_cascade_ ;
    wire \nx.n3085 ;
    wire \nx.n42_adj_689 ;
    wire \nx.n3103 ;
    wire \nx.n3097 ;
    wire \nx.n3164 ;
    wire \nx.n3097_cascade_ ;
    wire \nx.n3168 ;
    wire \nx.n35_adj_699_cascade_ ;
    wire \nx.n3101 ;
    wire \nx.n12337 ;
    wire \nx.n3109 ;
    wire \nx.n12349 ;
    wire \nx.n3174 ;
    wire \nx.n23_adj_700 ;
    wire \nx.n3107 ;
    wire \nx.n3162 ;
    wire \nx.n12327_cascade_ ;
    wire \nx.n3095 ;
    wire \nx.n3166 ;
    wire \nx.n3177 ;
    wire \nx.n3209 ;
    wire \nx.n3171 ;
    wire \nx.n3175 ;
    wire \nx.n3108 ;
    wire \nx.n3165 ;
    wire \nx.n3098 ;
    wire \nx.n13_adj_696_cascade_ ;
    wire \nx.n31_adj_702 ;
    wire \nx.n21_adj_701 ;
    wire \nx.n12325_cascade_ ;
    wire \nx.n12339 ;
    wire \nx.n12347 ;
    wire \nx.n3151 ;
    wire \nx.n61 ;
    wire \nx.n3099 ;
    wire neopxl_color_prev_7;
    wire \nx.n54 ;
    wire \nx.n43_adj_709_cascade_ ;
    wire \nx.n49_adj_710 ;
    wire state_3_N_377_1;
    wire \nx.n3084 ;
    wire \nx.n1177 ;
    wire bfn_2_29_0_;
    wire \nx.n1109 ;
    wire \nx.n1176 ;
    wire \nx.n10461 ;
    wire \nx.n10462 ;
    wire \nx.n1174 ;
    wire \nx.n10463 ;
    wire \nx.n10464 ;
    wire \nx.n10465 ;
    wire \nx.n1171 ;
    wire \nx.n10466 ;
    wire \nx.n10467 ;
    wire \nx.n1202 ;
    wire \nx.n1173 ;
    wire \nx.n1172 ;
    wire \nx.n1204 ;
    wire \nx.n1271 ;
    wire \nx.n1204_cascade_ ;
    wire \nx.n11_adj_624 ;
    wire \nx.n13 ;
    wire \nx.n1206 ;
    wire \nx.n1275 ;
    wire \nx.n1235_cascade_ ;
    wire \nx.n1208 ;
    wire \nx.n1175 ;
    wire \nx.n1136 ;
    wire \nx.n1207 ;
    wire \nx.n1274 ;
    wire \nx.n1207_cascade_ ;
    wire \nx.n1306_cascade_ ;
    wire \nx.n10_adj_626 ;
    wire bfn_2_31_0_;
    wire \nx.n10573 ;
    wire \nx.n10574 ;
    wire \nx.n10575 ;
    wire \nx.n10576 ;
    wire \nx.n10577 ;
    wire \nx.n10578 ;
    wire \nx.n10579 ;
    wire \nx.n10580 ;
    wire bfn_2_32_0_;
    wire \nx.n1301 ;
    wire \nx.n10581 ;
    wire \nx.n1302 ;
    wire \nx.n1369 ;
    wire neo_pixel_transmitter_t0_1;
    wire neo_pixel_transmitter_t0_31;
    wire neo_pixel_transmitter_t0_4;
    wire bfn_3_17_0_;
    wire \nx.n10479 ;
    wire \nx.n10480 ;
    wire \nx.n10481 ;
    wire \nx.n10482 ;
    wire \nx.n10483 ;
    wire \nx.n10484 ;
    wire \nx.n10485 ;
    wire \nx.n10486 ;
    wire bfn_3_18_0_;
    wire \nx.n10487 ;
    wire \nx.n10488 ;
    wire \nx.n10489 ;
    wire \nx.n10490 ;
    wire \nx.n10491 ;
    wire \nx.n10492 ;
    wire \nx.n10493 ;
    wire \nx.n10494 ;
    wire bfn_3_19_0_;
    wire \nx.n10495 ;
    wire \nx.n10496 ;
    wire \nx.n10497 ;
    wire \nx.n10498 ;
    wire \nx.n10499 ;
    wire \nx.n10500 ;
    wire \nx.n10501 ;
    wire \nx.n10502 ;
    wire bfn_3_20_0_;
    wire \nx.n10503 ;
    wire \nx.n10504 ;
    wire \nx.n10505 ;
    wire \nx.n10506 ;
    wire \nx.n10507 ;
    wire \nx.n10508 ;
    wire \nx.n10509 ;
    wire bfn_3_21_0_;
    wire \nx.n32_adj_651 ;
    wire timer_1;
    wire \nx.n11533 ;
    wire \nx.n10422 ;
    wire \nx.one_wire_N_528_2 ;
    wire \nx.n10423 ;
    wire \nx.n30_adj_598 ;
    wire timer_3;
    wire \nx.one_wire_N_528_3 ;
    wire \nx.n10424 ;
    wire \nx.n29 ;
    wire timer_4;
    wire \nx.one_wire_N_528_4 ;
    wire \nx.n10425 ;
    wire timer_5;
    wire \nx.n28 ;
    wire \nx.one_wire_N_528_5 ;
    wire \nx.n10426 ;
    wire timer_6;
    wire \nx.n27 ;
    wire \nx.one_wire_N_528_6 ;
    wire \nx.n10427 ;
    wire \nx.one_wire_N_528_7 ;
    wire \nx.n10428 ;
    wire \nx.n10429 ;
    wire \nx.n25 ;
    wire timer_8;
    wire \nx.one_wire_N_528_8 ;
    wire bfn_3_22_0_;
    wire \nx.one_wire_N_528_9 ;
    wire \nx.n10430 ;
    wire timer_10;
    wire \nx.one_wire_N_528_10 ;
    wire \nx.n10431 ;
    wire \nx.n10432 ;
    wire \nx.one_wire_N_528_11 ;
    wire timer_12;
    wire \nx.n21_adj_620 ;
    wire \nx.n10433 ;
    wire \nx.n12945 ;
    wire \nx.n10434 ;
    wire \nx.n12947 ;
    wire \nx.n19_adj_622 ;
    wire timer_14;
    wire \nx.n10435 ;
    wire \nx.n10436 ;
    wire \nx.n10436_THRU_CRY_0_THRU_CO ;
    wire \nx.n12949 ;
    wire \nx.n18_adj_623 ;
    wire timer_15;
    wire bfn_3_23_0_;
    wire \nx.n12951 ;
    wire \nx.n17 ;
    wire timer_16;
    wire \nx.n10437 ;
    wire \nx.n12953 ;
    wire \nx.n10438 ;
    wire \nx.n12955 ;
    wire \nx.n10439 ;
    wire \nx.n12957 ;
    wire \nx.n10440 ;
    wire \nx.n12959 ;
    wire \nx.n10441 ;
    wire \nx.n10442 ;
    wire \nx.n10442_THRU_CRY_0_THRU_CO ;
    wire \nx.n10442_THRU_CRY_1_THRU_CO ;
    wire \nx.n12961 ;
    wire bfn_3_24_0_;
    wire \nx.n12963 ;
    wire \nx.n10443 ;
    wire \nx.n12965 ;
    wire \nx.n10 ;
    wire timer_23;
    wire \nx.n10444 ;
    wire \nx.n12967 ;
    wire \nx.n9 ;
    wire timer_24;
    wire \nx.n10445 ;
    wire \nx.n12969 ;
    wire \nx.n10446 ;
    wire \nx.n12971 ;
    wire \nx.n7_adj_597 ;
    wire timer_26;
    wire \nx.n10447 ;
    wire \nx.n10448 ;
    wire GNDG0;
    wire \nx.n10448_THRU_CRY_0_THRU_CO ;
    wire \nx.n10448_THRU_CRY_1_THRU_CO ;
    wire \nx.n12973 ;
    wire bfn_3_25_0_;
    wire \nx.n12975 ;
    wire \nx.n10449 ;
    wire \nx.n12977 ;
    wire \nx.n10450 ;
    wire \nx.n12979 ;
    wire \nx.n10451 ;
    wire timer_31;
    wire \nx.n2 ;
    wire \nx.n12981 ;
    wire \nx.n10452 ;
    wire \nx.n7181 ;
    wire timer_27;
    wire neo_pixel_transmitter_t0_27;
    wire \nx.n6 ;
    wire \nx.n3077 ;
    wire bfn_3_26_0_;
    wire \nx.n3076 ;
    wire \nx.n10862 ;
    wire \nx.n3008 ;
    wire \nx.n3075 ;
    wire \nx.n10863 ;
    wire \nx.n3007 ;
    wire \nx.n3074 ;
    wire \nx.n10864 ;
    wire \nx.n3073 ;
    wire \nx.n10865 ;
    wire \nx.n3072 ;
    wire \nx.n10866 ;
    wire \nx.n3071 ;
    wire \nx.n10867 ;
    wire \nx.n3070 ;
    wire \nx.n10868 ;
    wire \nx.n10869 ;
    wire \nx.n3069 ;
    wire bfn_3_27_0_;
    wire \nx.n3001 ;
    wire \nx.n3068 ;
    wire \nx.n10870 ;
    wire \nx.n3067 ;
    wire \nx.n10871 ;
    wire \nx.n2999 ;
    wire \nx.n3066 ;
    wire \nx.n10872 ;
    wire \nx.n3065 ;
    wire \nx.n10873 ;
    wire \nx.n3064 ;
    wire \nx.n10874 ;
    wire \nx.n3063 ;
    wire \nx.n10875 ;
    wire \nx.n10876 ;
    wire \nx.n10877 ;
    wire bfn_3_28_0_;
    wire \nx.n10878 ;
    wire \nx.n3059 ;
    wire \nx.n10879 ;
    wire \nx.n10880 ;
    wire \nx.n10881 ;
    wire \nx.n10882 ;
    wire \nx.n3055 ;
    wire \nx.n10883 ;
    wire \nx.n3054 ;
    wire \nx.n10884 ;
    wire \nx.n10885 ;
    wire \nx.n3053 ;
    wire bfn_3_29_0_;
    wire \nx.n3052 ;
    wire \nx.n10886 ;
    wire \nx.n10887 ;
    wire \nx.n3083 ;
    wire \nx.n45_adj_707 ;
    wire \nx.n11_adj_628_cascade_ ;
    wire \nx.n16_adj_627 ;
    wire \nx.n1307 ;
    wire \nx.n1334_cascade_ ;
    wire \nx.n1374 ;
    wire \nx.n1277 ;
    wire \nx.n1309 ;
    wire \nx.n1376 ;
    wire \nx.n1309_cascade_ ;
    wire \nx.n1272 ;
    wire \nx.n1205 ;
    wire \nx.n1235 ;
    wire \nx.n1377 ;
    wire bfn_3_31_0_;
    wire \nx.n10582 ;
    wire \nx.n10583 ;
    wire \nx.n10584 ;
    wire \nx.n10585 ;
    wire \nx.n10586 ;
    wire \nx.n10587 ;
    wire \nx.n10588 ;
    wire \nx.n10589 ;
    wire bfn_3_32_0_;
    wire \nx.n10590 ;
    wire \nx.n10591 ;
    wire \nx.n1303 ;
    wire \nx.n1370 ;
    wire \nx.n1400 ;
    wire \nx.n3 ;
    wire timer_30;
    wire neo_pixel_transmitter_t0_30;
    wire \nx.n31_adj_650 ;
    wire \nx.n16_adj_661 ;
    wire timer_17;
    wire neo_pixel_transmitter_t0_17;
    wire timer_2;
    wire neo_pixel_transmitter_t0_2;
    wire timer_29;
    wire timer_9;
    wire neo_pixel_transmitter_t0_10;
    wire \nx.n23_adj_617 ;
    wire neo_pixel_transmitter_t0_29;
    wire \nx.n4 ;
    wire timer_11;
    wire timer_21;
    wire timer_13;
    wire neo_pixel_transmitter_t0_11;
    wire \nx.n22_adj_618 ;
    wire neo_pixel_transmitter_t0_13;
    wire \nx.n20 ;
    wire timer_7;
    wire \nx.n13159 ;
    wire neo_pixel_transmitter_t0_21;
    wire \nx.n12 ;
    wire timer_25;
    wire timer_18;
    wire \nx.n5 ;
    wire neo_pixel_transmitter_t0_25;
    wire \nx.n8 ;
    wire neo_pixel_transmitter_t0_18;
    wire \nx.n15 ;
    wire timer_28;
    wire neo_pixel_transmitter_t0_28;
    wire \nx.n2995_cascade_ ;
    wire \nx.n44_adj_681 ;
    wire \nx.n33_adj_682_cascade_ ;
    wire \nx.n48 ;
    wire \nx.n3005 ;
    wire neo_pixel_transmitter_t0_7;
    wire \nx.n26 ;
    wire \nx.n3006 ;
    wire \nx.n2899_cascade_ ;
    wire \nx.n2998 ;
    wire \nx.n2894_cascade_ ;
    wire \nx.n2985 ;
    wire \nx.n2985_cascade_ ;
    wire \nx.n2986 ;
    wire \nx.n40_adj_683 ;
    wire \nx.n43_adj_677 ;
    wire \nx.n40_adj_678 ;
    wire \nx.n47_cascade_ ;
    wire \nx.n2918_cascade_ ;
    wire \nx.n3000 ;
    wire \nx.n38_adj_676 ;
    wire \nx.n2996 ;
    wire \nx.n2997 ;
    wire \nx.n2987 ;
    wire \nx.n3004 ;
    wire \nx.n2988 ;
    wire \nx.n2988_cascade_ ;
    wire \nx.n41_adj_686 ;
    wire \nx.n2994_cascade_ ;
    wire \nx.n3002 ;
    wire \nx.n42_adj_684 ;
    wire \nx.n3009 ;
    wire \nx.n2992 ;
    wire \nx.n2989 ;
    wire \nx.n3056 ;
    wire \nx.n3104 ;
    wire \nx.n3088_cascade_ ;
    wire \nx.n44_adj_690 ;
    wire \nx.n3061 ;
    wire \nx.n2994 ;
    wire \nx.n2991 ;
    wire \nx.n3058 ;
    wire \nx.n3161 ;
    wire \nx.n12353 ;
    wire \nx.n3160 ;
    wire \nx.n12355 ;
    wire \nx.n12357_cascade_ ;
    wire \nx.n3159 ;
    wire \nx.n3158 ;
    wire \nx.n12359_cascade_ ;
    wire \nx.n3157 ;
    wire \nx.n12361_cascade_ ;
    wire \nx.n3090 ;
    wire \nx.n3156 ;
    wire \nx.n12363_cascade_ ;
    wire \nx.n3116 ;
    wire \nx.n3088 ;
    wire \nx.n12365_cascade_ ;
    wire \nx.n3155 ;
    wire \nx.n12367 ;
    wire \nx.n2990 ;
    wire \nx.n3057 ;
    wire \nx.n3089 ;
    wire \nx.bit_ctr_0 ;
    wire bfn_4_27_0_;
    wire \nx.bit_ctr_1 ;
    wire \nx.n10391 ;
    wire \nx.bit_ctr_2 ;
    wire \nx.n10392 ;
    wire \nx.bit_ctr_3 ;
    wire \nx.n10393 ;
    wire \nx.bit_ctr_4 ;
    wire \nx.n10394 ;
    wire \nx.n10395 ;
    wire \nx.n10396 ;
    wire \nx.n10397 ;
    wire \nx.n10398 ;
    wire bfn_4_28_0_;
    wire \nx.n10399 ;
    wire \nx.n10400 ;
    wire \nx.n10401 ;
    wire \nx.n10402 ;
    wire \nx.n10403 ;
    wire \nx.n10404 ;
    wire \nx.n10405 ;
    wire \nx.n10406 ;
    wire bfn_4_29_0_;
    wire \nx.n10407 ;
    wire \nx.n10408 ;
    wire \nx.n10409 ;
    wire \nx.n10410 ;
    wire \nx.n10411 ;
    wire \nx.n10412 ;
    wire \nx.n10413 ;
    wire \nx.n10414 ;
    wire \nx.bit_ctr_24 ;
    wire bfn_4_30_0_;
    wire \nx.n10415 ;
    wire \nx.n10416 ;
    wire \nx.n10417 ;
    wire \nx.n10418 ;
    wire \nx.n10419 ;
    wire \nx.n10420 ;
    wire \nx.n10421 ;
    wire \nx.n7230 ;
    wire \nx.n7411 ;
    wire \nx.n1308 ;
    wire \nx.n1375 ;
    wire \nx.n1373 ;
    wire \nx.n1306 ;
    wire \nx.n1371 ;
    wire \nx.n1304 ;
    wire \nx.n1305 ;
    wire \nx.n1372 ;
    wire \nx.n1334 ;
    wire \nx.n1404_cascade_ ;
    wire \nx.bit_ctr_23 ;
    wire \nx.n47_adj_706 ;
    wire \nx.n1404 ;
    wire \nx.n1471 ;
    wire \nx.bit_ctr_21 ;
    wire \nx.n1477 ;
    wire \nx.n1509_cascade_ ;
    wire \nx.n16_adj_629 ;
    wire \nx.n18_adj_630_cascade_ ;
    wire \nx.n13_adj_631 ;
    wire \nx.n1469 ;
    wire \nx.n1433_cascade_ ;
    wire \nx.n1402 ;
    wire \nx.n1501_cascade_ ;
    wire \nx.n9672 ;
    wire timer_22;
    wire timer_19;
    wire n13171;
    wire n13170;
    wire neo_pixel_transmitter_t0_9;
    wire \nx.n24 ;
    wire neo_pixel_transmitter_t0_19;
    wire \nx.n14 ;
    wire neopxl_color_prev_6;
    wire neopxl_color_prev_15;
    wire n11_adj_775;
    wire neopxl_color_prev_13;
    wire \nx.n13_adj_649 ;
    wire timer_20;
    wire neo_pixel_transmitter_t0_20;
    wire \nx.n2809_cascade_ ;
    wire \nx.n31_adj_613_cascade_ ;
    wire \nx.n39_adj_614 ;
    wire \nx.n2896_cascade_ ;
    wire \nx.n2898_cascade_ ;
    wire \nx.n42_adj_675_cascade_ ;
    wire \nx.n32_adj_674 ;
    wire \nx.n46 ;
    wire \nx.n2977 ;
    wire bfn_5_22_0_;
    wire \nx.n2976 ;
    wire \nx.n10837 ;
    wire \nx.n2908 ;
    wire \nx.n2975 ;
    wire \nx.n10838 ;
    wire \nx.n2907 ;
    wire \nx.n2974 ;
    wire \nx.n10839 ;
    wire \nx.n2906 ;
    wire \nx.n2973 ;
    wire \nx.n10840 ;
    wire \nx.n2972 ;
    wire \nx.n10841 ;
    wire \nx.n10842 ;
    wire \nx.n2970 ;
    wire \nx.n10843 ;
    wire \nx.n10844 ;
    wire \nx.n2969 ;
    wire bfn_5_23_0_;
    wire \nx.n2901 ;
    wire \nx.n2968 ;
    wire \nx.n10845 ;
    wire \nx.n2967 ;
    wire \nx.n10846 ;
    wire \nx.n2899 ;
    wire \nx.n2966 ;
    wire \nx.n10847 ;
    wire \nx.n2898 ;
    wire \nx.n2965 ;
    wire \nx.n10848 ;
    wire \nx.n2897 ;
    wire \nx.n2964 ;
    wire \nx.n10849 ;
    wire \nx.n2896 ;
    wire \nx.n2963 ;
    wire \nx.n10850 ;
    wire \nx.n2962 ;
    wire \nx.n10851 ;
    wire \nx.n10852 ;
    wire bfn_5_24_0_;
    wire \nx.n2960 ;
    wire \nx.n10853 ;
    wire \nx.n2959 ;
    wire \nx.n10854 ;
    wire \nx.n2958 ;
    wire \nx.n10855 ;
    wire \nx.n2957 ;
    wire \nx.n10856 ;
    wire \nx.n2956 ;
    wire \nx.n10857 ;
    wire \nx.n2955 ;
    wire \nx.n10858 ;
    wire \nx.n2954 ;
    wire \nx.n10859 ;
    wire \nx.n10860 ;
    wire \nx.n2953 ;
    wire bfn_5_25_0_;
    wire \nx.n10861 ;
    wire \nx.n2984 ;
    wire \nx.n2961 ;
    wire \nx.n2894 ;
    wire \nx.n2993 ;
    wire \nx.n3060 ;
    wire \nx.n2993_cascade_ ;
    wire \nx.n3092 ;
    wire \nx.n3091 ;
    wire \nx.n3092_cascade_ ;
    wire \nx.n46_adj_688 ;
    wire \nx.n50 ;
    wire \nx.n3093 ;
    wire \nx.n36_adj_687 ;
    wire \nx.n1077 ;
    wire bfn_5_26_0_;
    wire \nx.n10468 ;
    wire \nx.n10469 ;
    wire \nx.n10470 ;
    wire \nx.n10471 ;
    wire \nx.n10472 ;
    wire \nx.n10473 ;
    wire \nx.n1103 ;
    wire \nx.n46_adj_705 ;
    wire \nx.n1075 ;
    wire \nx.n1107 ;
    wire \nx.n1073 ;
    wire \nx.n1105 ;
    wire \nx.n11617_cascade_ ;
    wire \nx.n1076 ;
    wire \nx.n1037_cascade_ ;
    wire \nx.n1108 ;
    wire \nx.n1007 ;
    wire \nx.n1074 ;
    wire \nx.n1106 ;
    wire \nx.n1009 ;
    wire \nx.bit_ctr_25 ;
    wire \nx.n1009_cascade_ ;
    wire \nx.n7_adj_616 ;
    wire \nx.bit_ctr_5 ;
    wire \nx.bit_ctr_6 ;
    wire \nx.n44_adj_708 ;
    wire \nx.n1005 ;
    wire \nx.n1072 ;
    wire \nx.n1005_cascade_ ;
    wire \nx.n1037 ;
    wire \nx.n1104 ;
    wire \nx.n1008 ;
    wire \nx.n7084_cascade_ ;
    wire \nx.n838_cascade_ ;
    wire \nx.n12595_cascade_ ;
    wire \nx.n9618_cascade_ ;
    wire \nx.n608 ;
    wire \nx.n11738_cascade_ ;
    wire \nx.n708 ;
    wire \nx.n739_cascade_ ;
    wire \nx.n11738 ;
    wire \nx.n807 ;
    wire \nx.bit_ctr_31 ;
    wire \nx.n9618 ;
    wire \nx.bit_ctr_29 ;
    wire \nx.n11771_cascade_ ;
    wire \nx.n1470 ;
    wire \nx.n1403 ;
    wire \nx.bit_ctr_30 ;
    wire \nx.n48_adj_704 ;
    wire \nx.n1407 ;
    wire \nx.n1474 ;
    wire \nx.n1506_cascade_ ;
    wire \nx.n18_adj_632 ;
    wire \nx.n1475 ;
    wire \nx.n1408 ;
    wire \nx.n1401 ;
    wire \nx.n1468 ;
    wire \nx.n1472 ;
    wire \nx.n1405 ;
    wire \nx.n1473 ;
    wire \nx.n1406 ;
    wire neopxl_color_15;
    wire \nx.n2700_cascade_ ;
    wire \nx.n2801_cascade_ ;
    wire \nx.n29_adj_607 ;
    wire \nx.n37_adj_608_cascade_ ;
    wire \nx.n40_adj_609 ;
    wire \nx.n42_cascade_ ;
    wire \nx.n2720_cascade_ ;
    wire \nx.n2797_cascade_ ;
    wire bfn_6_21_0_;
    wire \nx.n2809 ;
    wire \nx.n2876 ;
    wire \nx.n10813 ;
    wire \nx.n2808 ;
    wire \nx.n2875 ;
    wire \nx.n10814 ;
    wire \nx.n2807 ;
    wire \nx.n2874 ;
    wire \nx.n10815 ;
    wire \nx.n10816 ;
    wire \nx.n2805 ;
    wire \nx.n2872 ;
    wire \nx.n10817 ;
    wire \nx.n10818 ;
    wire \nx.n10819 ;
    wire \nx.n10820 ;
    wire \nx.n2802 ;
    wire \nx.n2869 ;
    wire bfn_6_22_0_;
    wire \nx.n10821 ;
    wire \nx.n2800 ;
    wire \nx.n2867 ;
    wire \nx.n10822 ;
    wire \nx.n2799 ;
    wire \nx.n2866 ;
    wire \nx.n10823 ;
    wire \nx.n2798 ;
    wire \nx.n2865 ;
    wire \nx.n10824 ;
    wire \nx.n2797 ;
    wire \nx.n2864 ;
    wire \nx.n10825 ;
    wire \nx.n10826 ;
    wire \nx.n2795 ;
    wire \nx.n2862 ;
    wire \nx.n10827 ;
    wire \nx.n10828 ;
    wire bfn_6_23_0_;
    wire \nx.n10829 ;
    wire \nx.n10830 ;
    wire \nx.n10831 ;
    wire \nx.n10832 ;
    wire \nx.n10833 ;
    wire \nx.n10834 ;
    wire \nx.n10835 ;
    wire \nx.n10836 ;
    wire bfn_6_24_0_;
    wire \nx.n2885 ;
    wire \nx.n2858 ;
    wire \nx.n2791_cascade_ ;
    wire \nx.n2859 ;
    wire \nx.n2891 ;
    wire \nx.n2856 ;
    wire \nx.n2789_cascade_ ;
    wire \nx.n2995 ;
    wire \nx.n3062 ;
    wire \nx.n3017 ;
    wire \nx.n3094 ;
    wire \nx.n28_adj_660_cascade_ ;
    wire \nx.n16 ;
    wire \nx.n1928_cascade_ ;
    wire \nx.n1908_cascade_ ;
    wire \nx.n24_adj_648 ;
    wire \nx.n1877 ;
    wire \nx.n1829_cascade_ ;
    wire \nx.n1906_cascade_ ;
    wire \nx.n22_adj_605 ;
    wire \nx.n1006 ;
    wire \nx.n1804_cascade_ ;
    wire \nx.n19_cascade_ ;
    wire \nx.n26_adj_600 ;
    wire \nx.bit_ctr_27 ;
    wire \nx.bit_ctr_28 ;
    wire \nx.n739 ;
    wire \nx.bit_ctr_26 ;
    wire \nx.n977 ;
    wire bfn_6_28_0_;
    wire \nx.n7082 ;
    wire \nx.n976 ;
    wire \nx.n10474 ;
    wire \nx.n7342 ;
    wire \nx.n975 ;
    wire \nx.n10475 ;
    wire \nx.n974 ;
    wire \nx.n10476 ;
    wire \nx.n906 ;
    wire \nx.n973 ;
    wire \nx.n10477 ;
    wire \nx.n13064 ;
    wire \nx.n10478 ;
    wire \nx.n4_adj_596 ;
    wire \nx.n5260 ;
    wire \nx.n11559 ;
    wire \nx.n838 ;
    wire \nx.n11674 ;
    wire \nx.n20_adj_634 ;
    wire \nx.n1532_cascade_ ;
    wire \nx.n1606_cascade_ ;
    wire \nx.n22_adj_647_cascade_ ;
    wire \nx.n1631_cascade_ ;
    wire \nx.n19_adj_602 ;
    wire \nx.n1409 ;
    wire \nx.n1476 ;
    wire \nx.n1433 ;
    wire \nx.n1508_cascade_ ;
    wire \nx.n16_adj_633 ;
    wire \nx.n1599_cascade_ ;
    wire bfn_6_31_0_;
    wire \nx.n10592 ;
    wire \nx.n1508 ;
    wire \nx.n1575 ;
    wire \nx.n10593 ;
    wire \nx.n1507 ;
    wire \nx.n1574 ;
    wire \nx.n10594 ;
    wire \nx.n10595 ;
    wire \nx.n1505 ;
    wire \nx.n1572 ;
    wire \nx.n10596 ;
    wire \nx.n1504 ;
    wire \nx.n1571 ;
    wire \nx.n10597 ;
    wire \nx.n10598 ;
    wire \nx.n10599 ;
    wire \nx.n1502 ;
    wire \nx.n1569 ;
    wire bfn_6_32_0_;
    wire \nx.n1501 ;
    wire \nx.n1568 ;
    wire \nx.n10600 ;
    wire \nx.n1500 ;
    wire \nx.n1567 ;
    wire \nx.n10601 ;
    wire \nx.n1499 ;
    wire \nx.n10602 ;
    wire neopxl_color_13;
    wire n11683;
    wire timer_0;
    wire neo_pixel_transmitter_t0_0;
    wire \nx.n33_adj_652 ;
    wire pin_out_0;
    wire pin_out_1;
    wire \nx.bit_ctr_8 ;
    wire \nx.n2777 ;
    wire bfn_7_19_0_;
    wire \nx.n2776 ;
    wire \nx.n10790 ;
    wire \nx.n2708 ;
    wire \nx.n2775 ;
    wire \nx.n10791 ;
    wire \nx.n2707 ;
    wire \nx.n2774 ;
    wire \nx.n10792 ;
    wire \nx.n2706 ;
    wire \nx.n2773 ;
    wire \nx.n10793 ;
    wire \nx.n10794 ;
    wire \nx.n2771 ;
    wire \nx.n10795 ;
    wire \nx.n2770 ;
    wire \nx.n10796 ;
    wire \nx.n10797 ;
    wire \nx.n2702 ;
    wire \nx.n2769 ;
    wire bfn_7_20_0_;
    wire \nx.n2768 ;
    wire \nx.n10798 ;
    wire \nx.n2700 ;
    wire \nx.n2767 ;
    wire \nx.n10799 ;
    wire \nx.n2766 ;
    wire \nx.n10800 ;
    wire \nx.n2765 ;
    wire \nx.n10801 ;
    wire \nx.n2764 ;
    wire \nx.n10802 ;
    wire \nx.n2696 ;
    wire \nx.n2763 ;
    wire \nx.n10803 ;
    wire \nx.n2762 ;
    wire \nx.n10804 ;
    wire \nx.n10805 ;
    wire bfn_7_21_0_;
    wire \nx.n10806 ;
    wire \nx.n2759 ;
    wire \nx.n10807 ;
    wire \nx.n10808 ;
    wire \nx.n2757 ;
    wire \nx.n10809 ;
    wire \nx.n2756 ;
    wire \nx.n10810 ;
    wire \nx.n10811 ;
    wire \nx.n10812 ;
    wire neo_pixel_transmitter_t0_22;
    wire \nx.n11 ;
    wire \nx.n2761 ;
    wire \nx.n2860 ;
    wire \nx.n2793_cascade_ ;
    wire \nx.n2892 ;
    wire \nx.n2758 ;
    wire \nx.n2760 ;
    wire \nx.n2873 ;
    wire \nx.n2806 ;
    wire \nx.n2905 ;
    wire \nx.n2793 ;
    wire \nx.n2791 ;
    wire \nx.n2792 ;
    wire \nx.n2786 ;
    wire \nx.n38_adj_625_cascade_ ;
    wire \nx.n42_adj_635 ;
    wire \nx.n41_adj_643 ;
    wire \nx.n43_cascade_ ;
    wire \nx.n44 ;
    wire \nx.n2854 ;
    wire \nx.n2819_cascade_ ;
    wire \nx.n2886 ;
    wire \nx.n2789 ;
    wire \nx.n26_adj_615 ;
    wire \nx.n2863 ;
    wire \nx.n2796 ;
    wire \nx.n2895 ;
    wire \nx.n2877 ;
    wire \nx.bit_ctr_7 ;
    wire \nx.n2909 ;
    wire \nx.n2868 ;
    wire \nx.n2801 ;
    wire \nx.n2900 ;
    wire \nx.n2861 ;
    wire \nx.n2794 ;
    wire \nx.n2893 ;
    wire \nx.n2788 ;
    wire \nx.n2855 ;
    wire \nx.n2887 ;
    wire \nx.n2890 ;
    wire \nx.n2888 ;
    wire \nx.n2887_cascade_ ;
    wire \nx.n39_adj_679 ;
    wire \nx.n2803 ;
    wire \nx.n2870 ;
    wire \nx.n2902 ;
    wire \nx.n2871 ;
    wire \nx.n2903 ;
    wire \nx.n2790 ;
    wire \nx.n2819 ;
    wire \nx.n2857 ;
    wire \nx.n2889 ;
    wire \nx.bit_ctr_16 ;
    wire bfn_7_25_0_;
    wire \nx.n1909 ;
    wire \nx.n13435 ;
    wire \nx.n10642 ;
    wire \nx.n1908 ;
    wire \nx.n10643 ;
    wire \nx.n1907 ;
    wire \nx.n10644 ;
    wire \nx.n1906 ;
    wire \nx.n10645 ;
    wire \nx.n10646 ;
    wire \nx.n1904 ;
    wire \nx.n10647 ;
    wire \nx.n1903 ;
    wire \nx.n10648 ;
    wire \nx.n10649 ;
    wire bfn_7_26_0_;
    wire \nx.n10650 ;
    wire \nx.n10651 ;
    wire \nx.n1899 ;
    wire \nx.n10652 ;
    wire \nx.n10653 ;
    wire \nx.n10654 ;
    wire \nx.n10655 ;
    wire \nx.n1928 ;
    wire \nx.n10656 ;
    wire \nx.n1897 ;
    wire \nx.n1902 ;
    wire \nx.n10994 ;
    wire \nx.n13425 ;
    wire \nx.n1701_cascade_ ;
    wire \nx.n1801_cascade_ ;
    wire \nx.n23 ;
    wire \nx.n1577 ;
    wire \nx.bit_ctr_20 ;
    wire \nx.n1609_cascade_ ;
    wire \nx.n16_adj_646 ;
    wire \nx.n1570 ;
    wire \nx.n1503 ;
    wire \nx.bit_ctr_19 ;
    wire \nx.n1677 ;
    wire bfn_7_30_0_;
    wire \nx.n1609 ;
    wire \nx.n1676 ;
    wire \nx.n10603 ;
    wire \nx.n10604 ;
    wire \nx.n1607 ;
    wire \nx.n1674 ;
    wire \nx.n10605 ;
    wire \nx.n10606 ;
    wire \nx.n1672 ;
    wire \nx.n10607 ;
    wire \nx.n10608 ;
    wire \nx.n1603 ;
    wire \nx.n1670 ;
    wire \nx.n10609 ;
    wire \nx.n10610 ;
    wire \nx.n1602 ;
    wire \nx.n1669 ;
    wire bfn_7_31_0_;
    wire \nx.n10611 ;
    wire \nx.n10612 ;
    wire \nx.n1599 ;
    wire \nx.n1666 ;
    wire \nx.n10613 ;
    wire \nx.n1598 ;
    wire \nx.n10614 ;
    wire \nx.n1600 ;
    wire \nx.n1667 ;
    wire n7258_cascade_;
    wire n7236;
    wire n7270_cascade_;
    wire n7254;
    wire pin_out_5;
    wire n13152_cascade_;
    wire n13146;
    wire n13462_cascade_;
    wire n13153;
    wire pin_out_3;
    wire pin_out_2;
    wire n13147;
    wire n13168;
    wire n13167_cascade_;
    wire n13450;
    wire \nx.n2694 ;
    wire \nx.n2697 ;
    wire \nx.n2704 ;
    wire \nx.n2695 ;
    wire \nx.n2698 ;
    wire \nx.n2698_cascade_ ;
    wire \nx.n39_adj_610 ;
    wire \nx.n2703 ;
    wire \nx.n2709 ;
    wire \nx.n2592_cascade_ ;
    wire \nx.n2689 ;
    wire \nx.n2690 ;
    wire \nx.n2689_cascade_ ;
    wire \nx.n2691 ;
    wire \nx.n2701 ;
    wire \nx.n2105_cascade_ ;
    wire \nx.n2595_cascade_ ;
    wire \nx.n28_adj_663 ;
    wire \nx.n26_adj_664_cascade_ ;
    wire \nx.n25_adj_666 ;
    wire \nx.n2027_cascade_ ;
    wire \nx.n2099_cascade_ ;
    wire \nx.n2904 ;
    wire \nx.n2971 ;
    wire \nx.n2918 ;
    wire \nx.n3003 ;
    wire bfn_9_23_0_;
    wire \nx.n10657 ;
    wire \nx.n10658 ;
    wire \nx.n10659 ;
    wire \nx.n2006 ;
    wire \nx.n2073 ;
    wire \nx.n10660 ;
    wire \nx.n2005 ;
    wire \nx.n2072 ;
    wire \nx.n10661 ;
    wire \nx.n2004 ;
    wire \nx.n2071 ;
    wire \nx.n10662 ;
    wire \nx.n10663 ;
    wire \nx.n10664 ;
    wire bfn_9_24_0_;
    wire \nx.n2001 ;
    wire \nx.n2068 ;
    wire \nx.n10665 ;
    wire \nx.n2000 ;
    wire \nx.n2067 ;
    wire \nx.n10666 ;
    wire \nx.n1999 ;
    wire \nx.n2066 ;
    wire \nx.n10667 ;
    wire \nx.n10668 ;
    wire \nx.n10669 ;
    wire \nx.n1996 ;
    wire \nx.n2063 ;
    wire \nx.n10670 ;
    wire \nx.n10671 ;
    wire \nx.n10672 ;
    wire \nx.n1994 ;
    wire bfn_9_25_0_;
    wire \nx.n1901 ;
    wire \nx.n1905 ;
    wire \nx.n25_adj_606 ;
    wire \nx.n22 ;
    wire \nx.n1900 ;
    wire \nx.n1799_cascade_ ;
    wire \nx.n1898 ;
    wire \nx.n1797_cascade_ ;
    wire \nx.n1896 ;
    wire \nx.bit_ctr_17 ;
    wire \nx.bit_ctr_22 ;
    wire \nx.n30_adj_703 ;
    wire bfn_9_27_0_;
    wire \nx.n1809 ;
    wire \nx.n1876 ;
    wire \nx.n10628 ;
    wire \nx.n1808 ;
    wire \nx.n1875 ;
    wire \nx.n10629 ;
    wire \nx.n1807 ;
    wire \nx.n1874 ;
    wire \nx.n10630 ;
    wire \nx.n1873 ;
    wire \nx.n10631 ;
    wire \nx.n1805 ;
    wire \nx.n1872 ;
    wire \nx.n10632 ;
    wire \nx.n1804 ;
    wire \nx.n1871 ;
    wire \nx.n10633 ;
    wire \nx.n1870 ;
    wire \nx.n10634 ;
    wire \nx.n10635 ;
    wire \nx.n1869 ;
    wire bfn_9_28_0_;
    wire \nx.n1801 ;
    wire \nx.n1868 ;
    wire \nx.n10636 ;
    wire \nx.n1800 ;
    wire \nx.n1867 ;
    wire \nx.n10637 ;
    wire \nx.n1799 ;
    wire \nx.n1866 ;
    wire \nx.n10638 ;
    wire \nx.n1865 ;
    wire \nx.n10639 ;
    wire \nx.n1797 ;
    wire \nx.n1864 ;
    wire \nx.n10640 ;
    wire \nx.n1829 ;
    wire \nx.n10641 ;
    wire \nx.n1895 ;
    wire \nx.n1668 ;
    wire \nx.n1601 ;
    wire \nx.n1509 ;
    wire \nx.n1576 ;
    wire \nx.n1608_cascade_ ;
    wire \nx.n18 ;
    wire \nx.n1506 ;
    wire \nx.n1573 ;
    wire \nx.n1532 ;
    wire \nx.n1605 ;
    wire \nx.n1604 ;
    wire \nx.n1671 ;
    wire \nx.n1606 ;
    wire \nx.n1673 ;
    wire n21_cascade_;
    wire n6150;
    wire pin_out_6;
    wire n7262;
    wire pin_out_7;
    wire n8_adj_780;
    wire n8_adj_780_cascade_;
    wire n7274;
    wire \nx.n2677 ;
    wire bfn_10_17_0_;
    wire \nx.n2676 ;
    wire \nx.n10768 ;
    wire \nx.n2675 ;
    wire \nx.n10769 ;
    wire \nx.n2674 ;
    wire \nx.n10770 ;
    wire \nx.n10771 ;
    wire \nx.n2672 ;
    wire \nx.n10772 ;
    wire \nx.n2671 ;
    wire \nx.n10773 ;
    wire \nx.n2670 ;
    wire \nx.n10774 ;
    wire \nx.n10775 ;
    wire \nx.n2669 ;
    wire bfn_10_18_0_;
    wire \nx.n2668 ;
    wire \nx.n10776 ;
    wire \nx.n10777 ;
    wire \nx.n2666 ;
    wire \nx.n10778 ;
    wire \nx.n2665 ;
    wire \nx.n10779 ;
    wire \nx.n2664 ;
    wire \nx.n10780 ;
    wire \nx.n2663 ;
    wire \nx.n10781 ;
    wire \nx.n2595 ;
    wire \nx.n2662 ;
    wire \nx.n10782 ;
    wire \nx.n10783 ;
    wire bfn_10_19_0_;
    wire \nx.n10784 ;
    wire \nx.n2592 ;
    wire \nx.n2659 ;
    wire \nx.n10785 ;
    wire \nx.n2658 ;
    wire \nx.n10786 ;
    wire \nx.n2657 ;
    wire \nx.n10787 ;
    wire \nx.n10788 ;
    wire \nx.n10789 ;
    wire \nx.n2660 ;
    wire \nx.n2692 ;
    wire \nx.n34_adj_603_cascade_ ;
    wire \nx.n39_cascade_ ;
    wire \nx.n2621_cascade_ ;
    wire \nx.n2661 ;
    wire \nx.n2693 ;
    wire \nx.n2667 ;
    wire \nx.n2699 ;
    wire \nx.n2687 ;
    wire \nx.n2699_cascade_ ;
    wire \nx.n36 ;
    wire \nx.n41 ;
    wire \nx.n2656 ;
    wire \nx.n31_adj_655_cascade_ ;
    wire \nx.n24_adj_654 ;
    wire \nx.n36_adj_656_cascade_ ;
    wire \nx.n33_adj_659 ;
    wire \nx.n2423_cascade_ ;
    wire \nx.n2491_cascade_ ;
    wire \nx.n2394_cascade_ ;
    wire \nx.n2077 ;
    wire \nx.n2070 ;
    wire \nx.n2069 ;
    wire \nx.n2076 ;
    wire \nx.bit_ctr_15 ;
    wire \nx.n2003 ;
    wire \nx.n2009 ;
    wire \nx.n27_adj_665 ;
    wire \nx.n2074 ;
    wire \nx.n2064 ;
    wire \nx.n1997 ;
    wire \nx.n2062 ;
    wire \nx.n1995 ;
    wire \nx.n26_adj_667 ;
    wire \nx.n30_adj_668_cascade_ ;
    wire \nx.n28_adj_669 ;
    wire \nx.n2008 ;
    wire \nx.n2075 ;
    wire \nx.n2107_cascade_ ;
    wire \nx.n29_adj_670 ;
    wire \nx.n2065 ;
    wire \nx.n1998 ;
    wire \nx.n2027 ;
    wire \nx.n2097_cascade_ ;
    wire \nx.n27_adj_671 ;
    wire \nx.n2007 ;
    wire \nx.n2002 ;
    wire \nx.n22_adj_662 ;
    wire \nx.n1803 ;
    wire \nx.n22_adj_673_cascade_ ;
    wire \nx.n16_adj_672 ;
    wire \nx.n1798 ;
    wire \nx.n1608 ;
    wire \nx.n1675 ;
    wire \nx.n1631 ;
    wire \nx.n1707_cascade_ ;
    wire \nx.n1806 ;
    wire \nx.n20_adj_680 ;
    wire \nx.n24_adj_685 ;
    wire \nx.n1730_cascade_ ;
    wire \nx.n1802 ;
    wire \nx.bit_ctr_18 ;
    wire \nx.n1777 ;
    wire bfn_10_28_0_;
    wire \nx.n1709 ;
    wire \nx.n1776 ;
    wire \nx.n10615 ;
    wire \nx.n1708 ;
    wire \nx.n1775 ;
    wire \nx.n10616 ;
    wire \nx.n1707 ;
    wire \nx.n1774 ;
    wire \nx.n10617 ;
    wire \nx.n1706 ;
    wire \nx.n1773 ;
    wire \nx.n10618 ;
    wire \nx.n1705 ;
    wire \nx.n1772 ;
    wire \nx.n10619 ;
    wire \nx.n1704 ;
    wire \nx.n1771 ;
    wire \nx.n10620 ;
    wire \nx.n1703 ;
    wire \nx.n1770 ;
    wire \nx.n10621 ;
    wire \nx.n10622 ;
    wire \nx.n1702 ;
    wire \nx.n1769 ;
    wire bfn_10_29_0_;
    wire \nx.n1701 ;
    wire \nx.n1768 ;
    wire \nx.n10623 ;
    wire \nx.n1700 ;
    wire \nx.n1767 ;
    wire \nx.n10624 ;
    wire \nx.n1699 ;
    wire \nx.n1766 ;
    wire \nx.n10625 ;
    wire \nx.n1698 ;
    wire \nx.n1765 ;
    wire \nx.n10626 ;
    wire \nx.n1730 ;
    wire \nx.n1697 ;
    wire \nx.n10627 ;
    wire \nx.n1796 ;
    wire pin_oe_22;
    wire n6158;
    wire n8;
    wire n22_adj_740_cascade_;
    wire n5907;
    wire n6162;
    wire n6162_cascade_;
    wire n7278;
    wire n6156;
    wire n7266_cascade_;
    wire pin_out_4;
    wire \nx.n2609 ;
    wire \nx.bit_ctr_9 ;
    wire \nx.n2609_cascade_ ;
    wire \nx.n28_adj_599_cascade_ ;
    wire \nx.n35 ;
    wire \nx.n40 ;
    wire \nx.n2608 ;
    wire \nx.n2596 ;
    wire \nx.n2599 ;
    wire \nx.n2596_cascade_ ;
    wire \nx.n2604 ;
    wire \nx.n37 ;
    wire \nx.n2598 ;
    wire \nx.n38 ;
    wire \nx.n2602 ;
    wire \nx.n2606 ;
    wire \nx.n2673 ;
    wire \nx.n2606_cascade_ ;
    wire \nx.n2621 ;
    wire \nx.n2705 ;
    wire \nx.n2772 ;
    wire \nx.n2705_cascade_ ;
    wire \nx.n2804 ;
    wire \nx.n2594 ;
    wire \nx.n2504_cascade_ ;
    wire \nx.n2603 ;
    wire \nx.n2589 ;
    wire \nx.n2688 ;
    wire \nx.n2720 ;
    wire \nx.n2755 ;
    wire \nx.n2787 ;
    wire \nx.n2590 ;
    wire \nx.n2591 ;
    wire \nx.n2296_cascade_ ;
    wire \nx.n2395_cascade_ ;
    wire \nx.n2494_cascade_ ;
    wire \nx.n2593 ;
    wire \nx.n2293_cascade_ ;
    wire \nx.bit_ctr_14 ;
    wire bfn_11_23_0_;
    wire \nx.n2109 ;
    wire \nx.n13436 ;
    wire \nx.n10673 ;
    wire \nx.n2108 ;
    wire \nx.n10674 ;
    wire \nx.n2107 ;
    wire \nx.n10675 ;
    wire \nx.n2106 ;
    wire \nx.n10676 ;
    wire \nx.n2105 ;
    wire \nx.n10677 ;
    wire \nx.n2104 ;
    wire \nx.n10678 ;
    wire \nx.n2103 ;
    wire \nx.n10679 ;
    wire \nx.n10680 ;
    wire \nx.n2102 ;
    wire bfn_11_24_0_;
    wire \nx.n2101 ;
    wire \nx.n10681 ;
    wire \nx.n2100 ;
    wire \nx.n10682 ;
    wire \nx.n2099 ;
    wire \nx.n10683 ;
    wire \nx.n2098 ;
    wire \nx.n10684 ;
    wire \nx.n2097 ;
    wire \nx.n10685 ;
    wire \nx.n2096 ;
    wire \nx.n10686 ;
    wire \nx.n2095 ;
    wire \nx.n10687 ;
    wire \nx.n10688 ;
    wire \nx.n2094 ;
    wire bfn_11_25_0_;
    wire \nx.n2093 ;
    wire \nx.n2126 ;
    wire \nx.n10689 ;
    wire n12171;
    wire n6_adj_761;
    wire n15_cascade_;
    wire n14;
    wire n12091;
    wire n24_adj_720_cascade_;
    wire n11898;
    wire neopxl_color_7;
    wire n22_adj_724;
    wire n17_adj_765;
    wire n16_adj_764_cascade_;
    wire n10978;
    wire n36;
    wire n7166_cascade_;
    wire n6152;
    wire n8_adj_751_cascade_;
    wire n7294_cascade_;
    wire pin_out_11;
    wire n6154;
    wire n8_adj_744;
    wire n13048_cascade_;
    wire n13264;
    wire \nx.n2597 ;
    wire \nx.n2601 ;
    wire \nx.n2497_cascade_ ;
    wire \nx.n26_adj_611_cascade_ ;
    wire \nx.n33 ;
    wire \nx.n38_adj_612_cascade_ ;
    wire \nx.n2522_cascade_ ;
    wire \nx.n2600 ;
    wire \nx.n2605 ;
    wire \nx.n35_adj_639 ;
    wire \nx.bit_ctr_10 ;
    wire \nx.n2577 ;
    wire bfn_12_20_0_;
    wire \nx.n2509 ;
    wire \nx.n2576 ;
    wire \nx.n10747 ;
    wire \nx.n10748 ;
    wire \nx.n2574 ;
    wire \nx.n10749 ;
    wire \nx.n2573 ;
    wire \nx.n10750 ;
    wire \nx.n2505 ;
    wire \nx.n2572 ;
    wire \nx.n10751 ;
    wire \nx.n2571 ;
    wire \nx.n10752 ;
    wire \nx.n2570 ;
    wire \nx.n10753 ;
    wire \nx.n10754 ;
    wire \nx.n2569 ;
    wire bfn_12_21_0_;
    wire \nx.n2501 ;
    wire \nx.n2568 ;
    wire \nx.n10755 ;
    wire \nx.n2567 ;
    wire \nx.n10756 ;
    wire \nx.n2499 ;
    wire \nx.n2566 ;
    wire \nx.n10757 ;
    wire \nx.n2565 ;
    wire \nx.n10758 ;
    wire \nx.n2497 ;
    wire \nx.n2564 ;
    wire \nx.n10759 ;
    wire \nx.n2496 ;
    wire \nx.n2563 ;
    wire \nx.n10760 ;
    wire \nx.n2562 ;
    wire \nx.n10761 ;
    wire \nx.n10762 ;
    wire \nx.n2494 ;
    wire \nx.n2561 ;
    wire bfn_12_22_0_;
    wire \nx.n2493 ;
    wire \nx.n2560 ;
    wire \nx.n10763 ;
    wire \nx.n2492 ;
    wire \nx.n2559 ;
    wire \nx.n10764 ;
    wire \nx.n2491 ;
    wire \nx.n2558 ;
    wire \nx.n10765 ;
    wire \nx.n2557 ;
    wire \nx.n10766 ;
    wire \nx.n10767 ;
    wire \nx.n2588 ;
    wire \nx.n30_adj_640 ;
    wire \nx.n34_cascade_ ;
    wire \nx.n21 ;
    wire \nx.n2225_cascade_ ;
    wire \nx.n31 ;
    wire \nx.n28_adj_601 ;
    wire neopxl_color_12;
    wire neopxl_color_prev_12;
    wire \nx.n30 ;
    wire \nx.n22_adj_604 ;
    wire delay_counter_0;
    wire bfn_12_26_0_;
    wire delay_counter_1;
    wire n10517;
    wire delay_counter_2;
    wire n10518;
    wire delay_counter_3;
    wire n10519;
    wire delay_counter_4;
    wire n10520;
    wire delay_counter_5;
    wire n10521;
    wire delay_counter_6;
    wire n10522;
    wire delay_counter_7;
    wire n10523;
    wire n10524;
    wire delay_counter_8;
    wire bfn_12_27_0_;
    wire delay_counter_9;
    wire n10525;
    wire delay_counter_10;
    wire n10526;
    wire delay_counter_11;
    wire n10527;
    wire delay_counter_12;
    wire n10528;
    wire delay_counter_13;
    wire n10529;
    wire delay_counter_14;
    wire n10530;
    wire delay_counter_15;
    wire n10531;
    wire n10532;
    wire delay_counter_16;
    wire bfn_12_28_0_;
    wire delay_counter_17;
    wire n10533;
    wire delay_counter_18;
    wire n10534;
    wire delay_counter_19;
    wire n10535;
    wire delay_counter_20;
    wire n10536;
    wire delay_counter_21;
    wire n10537;
    wire delay_counter_22;
    wire n10538;
    wire delay_counter_23;
    wire n10539;
    wire n10540;
    wire delay_counter_24;
    wire bfn_12_29_0_;
    wire delay_counter_25;
    wire n10541;
    wire delay_counter_26;
    wire n10542;
    wire delay_counter_27;
    wire n10543;
    wire delay_counter_28;
    wire n10544;
    wire delay_counter_29;
    wire n10545;
    wire delay_counter_30;
    wire n10546;
    wire n10547;
    wire n7442;
    wire n10_adj_779_cascade_;
    wire n10_adj_779;
    wire n7290_cascade_;
    wire pin_out_10;
    wire n7135;
    wire n7155_cascade_;
    wire n6190;
    wire n6190_cascade_;
    wire n7334;
    wire n6170;
    wire n9415;
    wire pin_in_8;
    wire n13480_cascade_;
    wire current_pin_7__N_157_cascade_;
    wire pin_in_0;
    wire pin_in_10;
    wire n2289_cascade_;
    wire pin_in_6;
    wire n13453;
    wire n13364_cascade_;
    wire n150;
    wire n13483;
    wire n13360;
    wire \nx.n2575 ;
    wire \nx.n2522 ;
    wire \nx.n2607 ;
    wire \nx.n2495 ;
    wire \nx.n2503 ;
    wire \nx.n2503_cascade_ ;
    wire \nx.n36_adj_636 ;
    wire \nx.n2502 ;
    wire \nx.n2508 ;
    wire \nx.n2506 ;
    wire neopxl_color_5;
    wire n22_adj_730;
    wire \nx.n2498 ;
    wire \nx.n2404_cascade_ ;
    wire \nx.n34_adj_657 ;
    wire \nx.n2490 ;
    wire \nx.n2504 ;
    wire \nx.n22_adj_637_cascade_ ;
    wire \nx.n2507 ;
    wire \nx.n37_adj_638 ;
    wire \nx.n2500 ;
    wire \nx.n2300_cascade_ ;
    wire \nx.n33_adj_644 ;
    wire \nx.n34_adj_641 ;
    wire \nx.n32_cascade_ ;
    wire \nx.n2324_cascade_ ;
    wire \nx.bit_ctr_13 ;
    wire \nx.n2277 ;
    wire bfn_13_23_0_;
    wire \nx.n2209 ;
    wire \nx.n2276 ;
    wire \nx.n10690 ;
    wire \nx.n2208 ;
    wire \nx.n2275 ;
    wire \nx.n10691 ;
    wire \nx.n10692 ;
    wire \nx.n2206 ;
    wire \nx.n2273 ;
    wire \nx.n10693 ;
    wire \nx.n2205 ;
    wire \nx.n2272 ;
    wire \nx.n10694 ;
    wire \nx.n10695 ;
    wire \nx.n2203 ;
    wire \nx.n2270 ;
    wire \nx.n10696 ;
    wire \nx.n10697 ;
    wire bfn_13_24_0_;
    wire \nx.n2201 ;
    wire \nx.n2268 ;
    wire \nx.n10698 ;
    wire \nx.n10699 ;
    wire \nx.n10700 ;
    wire \nx.n10701 ;
    wire \nx.n2197 ;
    wire \nx.n2264 ;
    wire \nx.n10702 ;
    wire \nx.n2196 ;
    wire \nx.n2263 ;
    wire \nx.n10703 ;
    wire \nx.n2195 ;
    wire \nx.n2262 ;
    wire \nx.n10704 ;
    wire \nx.n10705 ;
    wire \nx.n2194 ;
    wire \nx.n2261 ;
    wire bfn_13_25_0_;
    wire \nx.n10706 ;
    wire \nx.n2192 ;
    wire \nx.n10707 ;
    wire n7155;
    wire n6166;
    wire n6166_cascade_;
    wire n7286;
    wire n7_adj_753_cascade_;
    wire pin_in_2;
    wire n22_adj_740;
    wire n21_adj_741_cascade_;
    wire n7128;
    wire n7150_cascade_;
    wire pin_in_11;
    wire n2355;
    wire n21_adj_714;
    wire n7_adj_719_cascade_;
    wire n7150;
    wire pin_in_9;
    wire n2337;
    wire n2343_cascade_;
    wire n2325;
    wire pin_in_3;
    wire pin_in_1;
    wire n2361;
    wire n13474_cascade_;
    wire pin_in_12;
    wire n13477;
    wire pin_in_13;
    wire pin_in_15;
    wire n2367;
    wire n33;
    wire n2379_cascade_;
    wire n45_adj_772;
    wire neopxl_color_4;
    wire n22_adj_732;
    wire n7232;
    wire n43;
    wire n52_adj_770;
    wire neopxl_color_6;
    wire n22_adj_728;
    wire \nx.bit_ctr_11 ;
    wire \nx.n2477 ;
    wire bfn_14_21_0_;
    wire \nx.n2409 ;
    wire \nx.n2476 ;
    wire \nx.n10727 ;
    wire \nx.n2408 ;
    wire \nx.n2475 ;
    wire \nx.n10728 ;
    wire \nx.n2407 ;
    wire \nx.n2474 ;
    wire \nx.n10729 ;
    wire \nx.n2473 ;
    wire \nx.n10730 ;
    wire \nx.n2405 ;
    wire \nx.n2472 ;
    wire \nx.n10731 ;
    wire \nx.n2404 ;
    wire \nx.n2471 ;
    wire \nx.n10732 ;
    wire \nx.n2470 ;
    wire \nx.n10733 ;
    wire \nx.n10734 ;
    wire \nx.n2469 ;
    wire bfn_14_22_0_;
    wire \nx.n2401 ;
    wire \nx.n2468 ;
    wire \nx.n10735 ;
    wire \nx.n2467 ;
    wire \nx.n10736 ;
    wire \nx.n2399 ;
    wire \nx.n2466 ;
    wire \nx.n10737 ;
    wire \nx.n2465 ;
    wire \nx.n10738 ;
    wire \nx.n2464 ;
    wire \nx.n10739 ;
    wire \nx.n2463 ;
    wire \nx.n10740 ;
    wire \nx.n2395 ;
    wire \nx.n2462 ;
    wire \nx.n10741 ;
    wire \nx.n10742 ;
    wire \nx.n2394 ;
    wire \nx.n2461 ;
    wire bfn_14_23_0_;
    wire \nx.n2393 ;
    wire \nx.n2460 ;
    wire \nx.n10743 ;
    wire \nx.n2392 ;
    wire \nx.n2459 ;
    wire \nx.n10744 ;
    wire \nx.n2458 ;
    wire \nx.n10745 ;
    wire \nx.n2423 ;
    wire \nx.n10746 ;
    wire \nx.n2489 ;
    wire \nx.n2207 ;
    wire \nx.n2274 ;
    wire \nx.n2391 ;
    wire \nx.n2271 ;
    wire \nx.n2204 ;
    wire \nx.n2265 ;
    wire \nx.n2198 ;
    wire \nx.n2297_cascade_ ;
    wire \nx.n9650 ;
    wire \nx.n31_adj_645 ;
    wire \nx.n2269 ;
    wire \nx.n2202 ;
    wire \nx.n2267 ;
    wire \nx.n2200 ;
    wire \nx.n2266 ;
    wire \nx.n2199 ;
    wire \nx.n2260 ;
    wire \nx.n2193 ;
    wire \nx.n2225 ;
    wire \nx.n2396 ;
    wire n13177_cascade_;
    wire LED_c;
    wire n13176;
    wire n21_adj_741;
    wire n6172;
    wire n7298;
    wire n6172_cascade_;
    wire n6174;
    wire n7302;
    wire n7_adj_753;
    wire n6176;
    wire n7306_cascade_;
    wire pin_out_9;
    wire n13162;
    wire n13161_cascade_;
    wire n8_adj_751;
    wire n6164;
    wire n7282_cascade_;
    wire pin_out_8;
    wire n6184;
    wire n7322_cascade_;
    wire n13471;
    wire n13465;
    wire n10_adj_736;
    wire pin_in_14;
    wire n7145;
    wire n7314;
    wire n6;
    wire n6182;
    wire n7318_cascade_;
    wire n9_adj_733;
    wire n6188;
    wire n7330;
    wire pin_out_18;
    wire pin_out_16;
    wire n13438_cascade_;
    wire pin_out_17;
    wire n13441_cascade_;
    wire n13142_cascade_;
    wire n13362;
    wire n149_cascade_;
    wire pin_out_19;
    wire n8_adj_746;
    wire n6186;
    wire n7326;
    wire n11_adj_734;
    wire n11_adj_734_cascade_;
    wire n36_adj_773;
    wire pin_out_21;
    wire pin_out_20;
    wire n19_adj_735_cascade_;
    wire n13141;
    wire n1;
    wire n8_adj_747;
    wire n9426;
    wire n6178;
    wire n7310_cascade_;
    wire \nx.n2398 ;
    wire \nx.n2397 ;
    wire neopxl_color_14;
    wire neopxl_color_prev_14;
    wire \nx.n2400 ;
    wire \nx.n2400_cascade_ ;
    wire \nx.n2403 ;
    wire \nx.n35_adj_658 ;
    wire \nx.n2402 ;
    wire \nx.n2406 ;
    wire \nx.bit_ctr_12 ;
    wire \nx.n2377 ;
    wire bfn_15_23_0_;
    wire \nx.n2309 ;
    wire \nx.n2376 ;
    wire \nx.n10708 ;
    wire \nx.n2308 ;
    wire \nx.n2375 ;
    wire \nx.n10709 ;
    wire \nx.n2307 ;
    wire \nx.n2374 ;
    wire \nx.n10710 ;
    wire \nx.n2306 ;
    wire \nx.n2373 ;
    wire \nx.n10711 ;
    wire \nx.n2305 ;
    wire \nx.n2372 ;
    wire \nx.n10712 ;
    wire \nx.n2304 ;
    wire \nx.n2371 ;
    wire \nx.n10713 ;
    wire \nx.n2303 ;
    wire \nx.n2370 ;
    wire \nx.n10714 ;
    wire \nx.n10715 ;
    wire \nx.n2302 ;
    wire \nx.n2369 ;
    wire bfn_15_24_0_;
    wire \nx.n2301 ;
    wire \nx.n2368 ;
    wire \nx.n10716 ;
    wire \nx.n2300 ;
    wire \nx.n2367 ;
    wire \nx.n10717 ;
    wire \nx.n2299 ;
    wire \nx.n2366 ;
    wire \nx.n10718 ;
    wire \nx.n2298 ;
    wire \nx.n2365 ;
    wire \nx.n10719 ;
    wire \nx.n2297 ;
    wire \nx.n2364 ;
    wire \nx.n10720 ;
    wire \nx.n2296 ;
    wire \nx.n2363 ;
    wire \nx.n10721 ;
    wire \nx.n2295 ;
    wire \nx.n2362 ;
    wire \nx.n10722 ;
    wire \nx.n10723 ;
    wire \nx.n2294 ;
    wire \nx.n2361 ;
    wire bfn_15_25_0_;
    wire \nx.n2293 ;
    wire \nx.n2360 ;
    wire \nx.n10724 ;
    wire \nx.n2292 ;
    wire \nx.n2359 ;
    wire \nx.n10725 ;
    wire CONSTANT_ONE_NET;
    wire \nx.n2291 ;
    wire \nx.n2324 ;
    wire \nx.n10726 ;
    wire \nx.n2390 ;
    wire n26;
    wire bfn_15_26_0_;
    wire n25;
    wire n10548;
    wire n24;
    wire n10549;
    wire n23;
    wire n10550;
    wire n22;
    wire n10551;
    wire n21_adj_737;
    wire n10552;
    wire n20;
    wire n10553;
    wire n19_adj_718;
    wire n10554;
    wire n10555;
    wire n18;
    wire bfn_15_27_0_;
    wire n17;
    wire n10556;
    wire n16;
    wire n10557;
    wire n15_adj_759;
    wire n10558;
    wire n14_adj_745;
    wire n10559;
    wire n13;
    wire n10560;
    wire n12;
    wire n10561;
    wire n11_adj_758;
    wire n10562;
    wire n10563;
    wire n10_adj_757;
    wire bfn_15_28_0_;
    wire n9;
    wire n10564;
    wire n8_adj_755;
    wire n10565;
    wire n7;
    wire n10566;
    wire n6_adj_756;
    wire n10567;
    wire blink_counter_21;
    wire n10568;
    wire blink_counter_22;
    wire n10569;
    wire blink_counter_23;
    wire n10570;
    wire n10571;
    wire blink_counter_24;
    wire bfn_15_29_0_;
    wire n10572;
    wire blink_counter_25;
    wire n45;
    wire bfn_16_15_0_;
    wire n10510;
    wire n10511;
    wire n10512;
    wire n10513;
    wire n10514;
    wire n10515;
    wire n10516;
    wire n8_adj_763_cascade_;
    wire current_pin_7__N_155;
    wire n7_adj_719;
    wire n21;
    wire current_pin_7__N_155_cascade_;
    wire n7166;
    wire n6180;
    wire n6971;
    wire n12135;
    wire n149;
    wire n7231;
    wire n12208;
    wire n7500_cascade_;
    wire pin_out_22;
    wire n8_adj_723;
    wire n4_adj_778;
    wire n7142;
    wire n7142_cascade_;
    wire counter_7;
    wire counter_6;
    wire n73;
    wire pin_in_7;
    wire n2385;
    wire n12123_cascade_;
    wire n48_adj_771;
    wire pin_in_4;
    wire n2313;
    wire n13144_cascade_;
    wire n13279;
    wire n14_adj_717;
    wire n11;
    wire n30;
    wire delay_counter_31;
    wire n11612;
    wire n11481;
    wire n13273;
    wire state_7_N_167_0;
    wire counter_3;
    wire counter_4;
    wire counter_0;
    wire counter_2;
    wire counter_1;
    wire n10_adj_762_cascade_;
    wire counter_5;
    wire n18_adj_742;
    wire n4;
    wire pin_out_13;
    wire pin_out_12;
    wire n13164_cascade_;
    wire n13468;
    wire n6_adj_748;
    wire pin_in_22;
    wire n6_adj_748_cascade_;
    wire pin_out_15;
    wire pin_out_14;
    wire n13165;
    wire bfn_17_17_0_;
    wire n10384;
    wire n10385;
    wire n10386;
    wire current_pin_4;
    wire n10387;
    wire current_pin_5;
    wire n10388;
    wire current_pin_6;
    wire n10389;
    wire n10390;
    wire current_pin_7;
    wire CLK_c;
    wire n7223;
    wire n7401;
    wire n7409;
    wire n11_adj_743;
    wire n2421;
    wire n2373;
    wire n11_adj_739;
    wire n39;
    wire n42;
    wire n40_cascade_;
    wire n41;
    wire pin_in_19;
    wire pin_in_18;
    wire pin_in_16;
    wire n13444_cascade_;
    wire pin_in_17;
    wire n13447;
    wire n14_adj_752;
    wire pin_in_5;
    wire n15_adj_749_cascade_;
    wire n15_adj_750;
    wire n37;
    wire current_pin_0;
    wire pin_in_21;
    wire pin_in_20;
    wire n19_adj_715;
    wire n6_adj_766;
    wire n54_adj_768;
    wire n53_adj_769;
    wire n13037_cascade_;
    wire n55_adj_767;
    wire n7249;
    wire n7249_cascade_;
    wire n7395;
    wire current_pin_3;
    wire n10;
    wire current_pin_2;
    wire current_pin_1;
    wire n9456;
    wire state_0;
    wire state_1;
    wire state_2;
    wire n15_adj_721;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__51103),
            .DIN(N__51102),
            .DOUT(N__51101),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__51103),
            .PADOUT(N__51102),
            .PADIN(N__51101),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__42351),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam NEOPXL_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam NEOPXL_pad_iopad.PULLUP=1'b0;
    IO_PAD NEOPXL_pad_iopad (
            .OE(N__51094),
            .DIN(N__51093),
            .DOUT(N__51092),
            .PACKAGEPIN(NEOPXL));
    defparam NEOPXL_pad_preio.PIN_TYPE=6'b011001;
    defparam NEOPXL_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO NEOPXL_pad_preio (
            .PADOEN(N__51094),
            .PADOUT(N__51093),
            .PADIN(N__51092),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__18414),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin0_iopad.PULLUP=1'b1;
    IO_PAD pin0_iopad (
            .OE(N__51085),
            .DIN(N__51084),
            .DOUT(N__51083),
            .PACKAGEPIN(USBPU));
    defparam pin0_preio.PIN_TYPE=6'b101001;
    defparam pin0_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin0_preio (
            .PADOEN(N__51085),
            .PADOUT(N__51084),
            .PADIN(N__51083),
            .CLOCKENABLE(),
            .DIN0(pin_in_0),
            .DIN1(),
            .DOUT0(N__28623),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35735));
    defparam pin1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin1_iopad.PULLUP=1'b1;
    IO_PAD pin1_iopad (
            .OE(N__51076),
            .DIN(N__51075),
            .DOUT(N__51074),
            .PACKAGEPIN(ENCODER0_A));
    defparam pin1_preio.PIN_TYPE=6'b101001;
    defparam pin1_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin1_preio (
            .PADOEN(N__51076),
            .PADOUT(N__51075),
            .PADIN(N__51074),
            .CLOCKENABLE(),
            .DIN0(pin_in_1),
            .DIN1(),
            .DOUT0(N__28587),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35801));
    defparam pin10_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin10_iopad.PULLUP=1'b1;
    IO_PAD pin10_iopad (
            .OE(N__51067),
            .DIN(N__51066),
            .DOUT(N__51065),
            .PACKAGEPIN(TX));
    defparam pin10_preio.PIN_TYPE=6'b101001;
    defparam pin10_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin10_preio (
            .PADOEN(N__51067),
            .PADOUT(N__51066),
            .PADIN(N__51065),
            .CLOCKENABLE(),
            .DIN0(pin_in_10),
            .DIN1(),
            .DOUT0(N__38943),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35670));
    defparam pin11_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin11_iopad.PULLUP=1'b1;
    IO_PAD pin11_iopad (
            .OE(N__51058),
            .DIN(N__51057),
            .DOUT(N__51056),
            .PACKAGEPIN(RX));
    defparam pin11_preio.PIN_TYPE=6'b101001;
    defparam pin11_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin11_preio (
            .PADOEN(N__51058),
            .PADOUT(N__51057),
            .PADIN(N__51056),
            .CLOCKENABLE(),
            .DIN0(pin_in_11),
            .DIN1(),
            .DOUT0(N__37560),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35734));
    defparam pin12_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin12_iopad.PULLUP=1'b1;
    IO_PAD pin12_iopad (
            .OE(N__51049),
            .DIN(N__51048),
            .DOUT(N__51047),
            .PACKAGEPIN(CS_CLK));
    defparam pin12_preio.PIN_TYPE=6'b101001;
    defparam pin12_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin12_preio (
            .PADOEN(N__51049),
            .PADOUT(N__51048),
            .PADIN(N__51047),
            .CLOCKENABLE(),
            .DIN0(pin_in_12),
            .DIN1(),
            .DOUT0(N__48045),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35723));
    defparam pin13_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin13_iopad.PULLUP=1'b1;
    IO_PAD pin13_iopad (
            .OE(N__51040),
            .DIN(N__51039),
            .DOUT(N__51038),
            .PACKAGEPIN(CS));
    defparam pin13_preio.PIN_TYPE=6'b101001;
    defparam pin13_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin13_preio (
            .PADOEN(N__51040),
            .PADOUT(N__51039),
            .PADIN(N__51038),
            .CLOCKENABLE(),
            .DIN0(pin_in_13),
            .DIN1(),
            .DOUT0(N__48084),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35737));
    defparam pin14_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin14_iopad.PULLUP=1'b1;
    IO_PAD pin14_iopad (
            .OE(N__51031),
            .DIN(N__51030),
            .DOUT(N__51029),
            .PACKAGEPIN(CS_MISO));
    defparam pin14_preio.PIN_TYPE=6'b101001;
    defparam pin14_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin14_preio (
            .PADOEN(N__51031),
            .PADOUT(N__51030),
            .PADIN(N__51029),
            .CLOCKENABLE(),
            .DIN0(pin_in_14),
            .DIN1(),
            .DOUT0(N__47850),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35668));
    defparam pin15_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin15_iopad.PULLUP=1'b1;
    IO_PAD pin15_iopad (
            .OE(N__51022),
            .DIN(N__51021),
            .DOUT(N__51020),
            .PACKAGEPIN(SCL));
    defparam pin15_preio.PIN_TYPE=6'b101001;
    defparam pin15_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin15_preio (
            .PADOEN(N__51022),
            .PADOUT(N__51021),
            .PADIN(N__51020),
            .CLOCKENABLE(),
            .DIN0(pin_in_15),
            .DIN1(),
            .DOUT0(N__47882),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35768));
    defparam pin16_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin16_iopad.PULLUP=1'b1;
    IO_PAD pin16_iopad (
            .OE(N__51013),
            .DIN(N__51012),
            .DOUT(N__51011),
            .PACKAGEPIN(SDA));
    defparam pin16_preio.PIN_TYPE=6'b101001;
    defparam pin16_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin16_preio (
            .PADOEN(N__51013),
            .PADOUT(N__51012),
            .PADIN(N__51011),
            .CLOCKENABLE(),
            .DIN0(pin_in_16),
            .DIN1(),
            .DOUT0(N__43101),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35793));
    defparam pin17_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin17_iopad.PULLUP=1'b1;
    IO_PAD pin17_iopad (
            .OE(N__51004),
            .DIN(N__51003),
            .DOUT(N__51002),
            .PACKAGEPIN(INLC));
    defparam pin17_preio.PIN_TYPE=6'b101001;
    defparam pin17_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin17_preio (
            .PADOEN(N__51004),
            .PADOUT(N__51003),
            .PADIN(N__51002),
            .CLOCKENABLE(),
            .DIN0(pin_in_17),
            .DIN1(),
            .DOUT0(N__43065),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35796));
    defparam pin18_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin18_iopad.PULLUP=1'b1;
    IO_PAD pin18_iopad (
            .OE(N__50995),
            .DIN(N__50994),
            .DOUT(N__50993),
            .PACKAGEPIN(INHC));
    defparam pin18_preio.PIN_TYPE=6'b101001;
    defparam pin18_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin18_preio (
            .PADOEN(N__50995),
            .PADOUT(N__50994),
            .PADIN(N__50993),
            .CLOCKENABLE(),
            .DIN0(pin_in_18),
            .DIN1(),
            .DOUT0(N__42555),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35795));
    defparam pin19_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin19_iopad.PULLUP=1'b1;
    IO_PAD pin19_iopad (
            .OE(N__50986),
            .DIN(N__50985),
            .DOUT(N__50984),
            .PACKAGEPIN(INLB));
    defparam pin19_preio.PIN_TYPE=6'b101001;
    defparam pin19_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin19_preio (
            .PADOEN(N__50986),
            .PADOUT(N__50985),
            .PADIN(N__50984),
            .CLOCKENABLE(),
            .DIN0(pin_in_19),
            .DIN1(),
            .DOUT0(N__43011),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35772));
    defparam pin2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin2_iopad.PULLUP=1'b1;
    IO_PAD pin2_iopad (
            .OE(N__50977),
            .DIN(N__50976),
            .DOUT(N__50975),
            .PACKAGEPIN(ENCODER0_B));
    defparam pin2_preio.PIN_TYPE=6'b101001;
    defparam pin2_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin2_preio (
            .PADOEN(N__50977),
            .PADOUT(N__50976),
            .PADIN(N__50975),
            .CLOCKENABLE(),
            .DIN0(pin_in_2),
            .DIN1(),
            .DOUT0(N__31374),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35725));
    defparam pin20_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin20_iopad.PULLUP=1'b1;
    IO_PAD pin20_iopad (
            .OE(N__50968),
            .DIN(N__50967),
            .DOUT(N__50966),
            .PACKAGEPIN(INHB));
    defparam pin20_preio.PIN_TYPE=6'b101001;
    defparam pin20_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin20_preio (
            .PADOEN(N__50968),
            .PADOUT(N__50967),
            .PADIN(N__50966),
            .CLOCKENABLE(),
            .DIN0(pin_in_20),
            .DIN1(),
            .DOUT0(N__42867),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35794));
    defparam pin21_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin21_iopad.PULLUP=1'b1;
    IO_PAD pin21_iopad (
            .OE(N__50959),
            .DIN(N__50958),
            .DOUT(N__50957),
            .PACKAGEPIN(INLA));
    defparam pin21_preio.PIN_TYPE=6'b101001;
    defparam pin21_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin21_preio (
            .PADOEN(N__50959),
            .PADOUT(N__50958),
            .PADIN(N__50957),
            .CLOCKENABLE(),
            .DIN0(pin_in_21),
            .DIN1(),
            .DOUT0(N__42909),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35736));
    defparam pin22_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin22_iopad.PULLUP=1'b1;
    IO_PAD pin22_iopad (
            .OE(N__50950),
            .DIN(N__50949),
            .DOUT(N__50948),
            .PACKAGEPIN(INHA));
    defparam pin22_preio.PIN_TYPE=6'b101001;
    defparam pin22_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin22_preio (
            .PADOEN(N__50950),
            .PADOUT(N__50949),
            .PADIN(N__50948),
            .CLOCKENABLE(),
            .DIN0(pin_in_22),
            .DIN1(),
            .DOUT0(N__47337),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35679));
    defparam pin3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin3_iopad.PULLUP=1'b1;
    IO_PAD pin3_iopad (
            .OE(N__50941),
            .DIN(N__50940),
            .DOUT(N__50939),
            .PACKAGEPIN(ENCODER1_A));
    defparam pin3_preio.PIN_TYPE=6'b101001;
    defparam pin3_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin3_preio (
            .PADOEN(N__50941),
            .PADOUT(N__50940),
            .PADIN(N__50939),
            .CLOCKENABLE(),
            .DIN0(pin_in_3),
            .DIN1(),
            .DOUT0(N__31401),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35724));
    defparam pin4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin4_iopad.PULLUP=1'b1;
    IO_PAD pin4_iopad (
            .OE(N__50932),
            .DIN(N__50931),
            .DOUT(N__50930),
            .PACKAGEPIN(ENCODER1_B));
    defparam pin4_preio.PIN_TYPE=6'b101001;
    defparam pin4_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin4_preio (
            .PADOEN(N__50932),
            .PADOUT(N__50931),
            .PADIN(N__50930),
            .CLOCKENABLE(),
            .DIN0(pin_in_4),
            .DIN1(),
            .DOUT0(N__35964),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35733));
    defparam pin5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin5_iopad.PULLUP=1'b1;
    IO_PAD pin5_iopad (
            .OE(N__50923),
            .DIN(N__50922),
            .DOUT(N__50921),
            .PACKAGEPIN(HALL1));
    defparam pin5_preio.PIN_TYPE=6'b101001;
    defparam pin5_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin5_preio (
            .PADOEN(N__50923),
            .PADOUT(N__50922),
            .PADIN(N__50921),
            .CLOCKENABLE(),
            .DIN0(pin_in_5),
            .DIN1(),
            .DOUT0(N__31230),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35800));
    defparam pin6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin6_iopad.PULLUP=1'b1;
    IO_PAD pin6_iopad (
            .OE(N__50914),
            .DIN(N__50913),
            .DOUT(N__50912),
            .PACKAGEPIN(HALL2));
    defparam pin6_preio.PIN_TYPE=6'b101001;
    defparam pin6_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin6_preio (
            .PADOEN(N__50914),
            .PADOUT(N__50913),
            .PADIN(N__50912),
            .CLOCKENABLE(),
            .DIN0(pin_in_6),
            .DIN1(),
            .DOUT0(N__33561),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35782));
    defparam pin7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin7_iopad.PULLUP=1'b1;
    IO_PAD pin7_iopad (
            .OE(N__50905),
            .DIN(N__50904),
            .DOUT(N__50903),
            .PACKAGEPIN(HALL3));
    defparam pin7_preio.PIN_TYPE=6'b101001;
    defparam pin7_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin7_preio (
            .PADOEN(N__50905),
            .PADOUT(N__50904),
            .PADIN(N__50903),
            .CLOCKENABLE(),
            .DIN0(pin_in_7),
            .DIN1(),
            .DOUT0(N__33516),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35783));
    defparam pin8_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin8_iopad.PULLUP=1'b1;
    IO_PAD pin8_iopad (
            .OE(N__50896),
            .DIN(N__50895),
            .DOUT(N__50894),
            .PACKAGEPIN(FAULT_N));
    defparam pin8_preio.PIN_TYPE=6'b101001;
    defparam pin8_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin8_preio (
            .PADOEN(N__50896),
            .PADOUT(N__50895),
            .PADIN(N__50894),
            .CLOCKENABLE(),
            .DIN0(pin_in_8),
            .DIN1(),
            .DOUT0(N__42411),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35802));
    defparam pin9_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin9_iopad.PULLUP=1'b1;
    IO_PAD pin9_iopad (
            .OE(N__50887),
            .DIN(N__50886),
            .DOUT(N__50885),
            .PACKAGEPIN(DE));
    defparam pin9_preio.PIN_TYPE=6'b101001;
    defparam pin9_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin9_preio (
            .PADOEN(N__50887),
            .PADOUT(N__50886),
            .PADIN(N__50885),
            .CLOCKENABLE(),
            .DIN0(pin_in_9),
            .DIN1(),
            .DOUT0(N__42507),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35669));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__50878),
            .DIN(N__50877),
            .DOUT(N__50876),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__50878),
            .PADOUT(N__50877),
            .PADIN(N__50876),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__12374 (
            .O(N__50859),
            .I(N__50856));
    LocalMux I__12373 (
            .O(N__50856),
            .I(n6_adj_766));
    InMux I__12372 (
            .O(N__50853),
            .I(N__50850));
    LocalMux I__12371 (
            .O(N__50850),
            .I(N__50847));
    Odrv4 I__12370 (
            .O(N__50847),
            .I(n54_adj_768));
    InMux I__12369 (
            .O(N__50844),
            .I(N__50841));
    LocalMux I__12368 (
            .O(N__50841),
            .I(N__50838));
    Span4Mux_h I__12367 (
            .O(N__50838),
            .I(N__50835));
    Odrv4 I__12366 (
            .O(N__50835),
            .I(n53_adj_769));
    CascadeMux I__12365 (
            .O(N__50832),
            .I(n13037_cascade_));
    InMux I__12364 (
            .O(N__50829),
            .I(N__50826));
    LocalMux I__12363 (
            .O(N__50826),
            .I(N__50823));
    Odrv4 I__12362 (
            .O(N__50823),
            .I(n55_adj_767));
    CEMux I__12361 (
            .O(N__50820),
            .I(N__50817));
    LocalMux I__12360 (
            .O(N__50817),
            .I(N__50812));
    CEMux I__12359 (
            .O(N__50816),
            .I(N__50809));
    InMux I__12358 (
            .O(N__50815),
            .I(N__50806));
    Span4Mux_h I__12357 (
            .O(N__50812),
            .I(N__50803));
    LocalMux I__12356 (
            .O(N__50809),
            .I(N__50800));
    LocalMux I__12355 (
            .O(N__50806),
            .I(N__50797));
    Odrv4 I__12354 (
            .O(N__50803),
            .I(n7249));
    Odrv12 I__12353 (
            .O(N__50800),
            .I(n7249));
    Odrv4 I__12352 (
            .O(N__50797),
            .I(n7249));
    CascadeMux I__12351 (
            .O(N__50790),
            .I(n7249_cascade_));
    SRMux I__12350 (
            .O(N__50787),
            .I(N__50784));
    LocalMux I__12349 (
            .O(N__50784),
            .I(N__50781));
    Odrv12 I__12348 (
            .O(N__50781),
            .I(n7395));
    CascadeMux I__12347 (
            .O(N__50778),
            .I(N__50774));
    InMux I__12346 (
            .O(N__50777),
            .I(N__50767));
    InMux I__12345 (
            .O(N__50774),
            .I(N__50762));
    InMux I__12344 (
            .O(N__50773),
            .I(N__50762));
    InMux I__12343 (
            .O(N__50772),
            .I(N__50749));
    InMux I__12342 (
            .O(N__50771),
            .I(N__50744));
    InMux I__12341 (
            .O(N__50770),
            .I(N__50744));
    LocalMux I__12340 (
            .O(N__50767),
            .I(N__50739));
    LocalMux I__12339 (
            .O(N__50762),
            .I(N__50739));
    InMux I__12338 (
            .O(N__50761),
            .I(N__50734));
    InMux I__12337 (
            .O(N__50760),
            .I(N__50734));
    InMux I__12336 (
            .O(N__50759),
            .I(N__50731));
    InMux I__12335 (
            .O(N__50758),
            .I(N__50727));
    CascadeMux I__12334 (
            .O(N__50757),
            .I(N__50723));
    InMux I__12333 (
            .O(N__50756),
            .I(N__50718));
    InMux I__12332 (
            .O(N__50755),
            .I(N__50715));
    CascadeMux I__12331 (
            .O(N__50754),
            .I(N__50709));
    InMux I__12330 (
            .O(N__50753),
            .I(N__50706));
    InMux I__12329 (
            .O(N__50752),
            .I(N__50703));
    LocalMux I__12328 (
            .O(N__50749),
            .I(N__50696));
    LocalMux I__12327 (
            .O(N__50744),
            .I(N__50696));
    Span4Mux_v I__12326 (
            .O(N__50739),
            .I(N__50696));
    LocalMux I__12325 (
            .O(N__50734),
            .I(N__50691));
    LocalMux I__12324 (
            .O(N__50731),
            .I(N__50691));
    InMux I__12323 (
            .O(N__50730),
            .I(N__50688));
    LocalMux I__12322 (
            .O(N__50727),
            .I(N__50684));
    InMux I__12321 (
            .O(N__50726),
            .I(N__50675));
    InMux I__12320 (
            .O(N__50723),
            .I(N__50675));
    InMux I__12319 (
            .O(N__50722),
            .I(N__50675));
    InMux I__12318 (
            .O(N__50721),
            .I(N__50675));
    LocalMux I__12317 (
            .O(N__50718),
            .I(N__50670));
    LocalMux I__12316 (
            .O(N__50715),
            .I(N__50670));
    InMux I__12315 (
            .O(N__50714),
            .I(N__50665));
    InMux I__12314 (
            .O(N__50713),
            .I(N__50665));
    InMux I__12313 (
            .O(N__50712),
            .I(N__50662));
    InMux I__12312 (
            .O(N__50709),
            .I(N__50659));
    LocalMux I__12311 (
            .O(N__50706),
            .I(N__50656));
    LocalMux I__12310 (
            .O(N__50703),
            .I(N__50653));
    Span4Mux_h I__12309 (
            .O(N__50696),
            .I(N__50648));
    Span4Mux_v I__12308 (
            .O(N__50691),
            .I(N__50648));
    LocalMux I__12307 (
            .O(N__50688),
            .I(N__50645));
    InMux I__12306 (
            .O(N__50687),
            .I(N__50642));
    Span4Mux_v I__12305 (
            .O(N__50684),
            .I(N__50633));
    LocalMux I__12304 (
            .O(N__50675),
            .I(N__50633));
    Span4Mux_v I__12303 (
            .O(N__50670),
            .I(N__50633));
    LocalMux I__12302 (
            .O(N__50665),
            .I(N__50633));
    LocalMux I__12301 (
            .O(N__50662),
            .I(current_pin_3));
    LocalMux I__12300 (
            .O(N__50659),
            .I(current_pin_3));
    Odrv4 I__12299 (
            .O(N__50656),
            .I(current_pin_3));
    Odrv4 I__12298 (
            .O(N__50653),
            .I(current_pin_3));
    Odrv4 I__12297 (
            .O(N__50648),
            .I(current_pin_3));
    Odrv12 I__12296 (
            .O(N__50645),
            .I(current_pin_3));
    LocalMux I__12295 (
            .O(N__50642),
            .I(current_pin_3));
    Odrv4 I__12294 (
            .O(N__50633),
            .I(current_pin_3));
    InMux I__12293 (
            .O(N__50616),
            .I(N__50612));
    CascadeMux I__12292 (
            .O(N__50615),
            .I(N__50608));
    LocalMux I__12291 (
            .O(N__50612),
            .I(N__50604));
    InMux I__12290 (
            .O(N__50611),
            .I(N__50599));
    InMux I__12289 (
            .O(N__50608),
            .I(N__50599));
    CascadeMux I__12288 (
            .O(N__50607),
            .I(N__50596));
    Span4Mux_v I__12287 (
            .O(N__50604),
            .I(N__50590));
    LocalMux I__12286 (
            .O(N__50599),
            .I(N__50590));
    InMux I__12285 (
            .O(N__50596),
            .I(N__50587));
    InMux I__12284 (
            .O(N__50595),
            .I(N__50584));
    Span4Mux_h I__12283 (
            .O(N__50590),
            .I(N__50579));
    LocalMux I__12282 (
            .O(N__50587),
            .I(N__50579));
    LocalMux I__12281 (
            .O(N__50584),
            .I(n10));
    Odrv4 I__12280 (
            .O(N__50579),
            .I(n10));
    CascadeMux I__12279 (
            .O(N__50574),
            .I(N__50570));
    InMux I__12278 (
            .O(N__50573),
            .I(N__50559));
    InMux I__12277 (
            .O(N__50570),
            .I(N__50551));
    InMux I__12276 (
            .O(N__50569),
            .I(N__50548));
    InMux I__12275 (
            .O(N__50568),
            .I(N__50545));
    CascadeMux I__12274 (
            .O(N__50567),
            .I(N__50541));
    CascadeMux I__12273 (
            .O(N__50566),
            .I(N__50538));
    InMux I__12272 (
            .O(N__50565),
            .I(N__50528));
    InMux I__12271 (
            .O(N__50564),
            .I(N__50525));
    InMux I__12270 (
            .O(N__50563),
            .I(N__50520));
    InMux I__12269 (
            .O(N__50562),
            .I(N__50520));
    LocalMux I__12268 (
            .O(N__50559),
            .I(N__50517));
    InMux I__12267 (
            .O(N__50558),
            .I(N__50512));
    InMux I__12266 (
            .O(N__50557),
            .I(N__50512));
    InMux I__12265 (
            .O(N__50556),
            .I(N__50509));
    InMux I__12264 (
            .O(N__50555),
            .I(N__50506));
    InMux I__12263 (
            .O(N__50554),
            .I(N__50503));
    LocalMux I__12262 (
            .O(N__50551),
            .I(N__50500));
    LocalMux I__12261 (
            .O(N__50548),
            .I(N__50496));
    LocalMux I__12260 (
            .O(N__50545),
            .I(N__50493));
    InMux I__12259 (
            .O(N__50544),
            .I(N__50487));
    InMux I__12258 (
            .O(N__50541),
            .I(N__50482));
    InMux I__12257 (
            .O(N__50538),
            .I(N__50482));
    InMux I__12256 (
            .O(N__50537),
            .I(N__50479));
    InMux I__12255 (
            .O(N__50536),
            .I(N__50476));
    InMux I__12254 (
            .O(N__50535),
            .I(N__50473));
    InMux I__12253 (
            .O(N__50534),
            .I(N__50470));
    InMux I__12252 (
            .O(N__50533),
            .I(N__50467));
    InMux I__12251 (
            .O(N__50532),
            .I(N__50462));
    InMux I__12250 (
            .O(N__50531),
            .I(N__50462));
    LocalMux I__12249 (
            .O(N__50528),
            .I(N__50459));
    LocalMux I__12248 (
            .O(N__50525),
            .I(N__50454));
    LocalMux I__12247 (
            .O(N__50520),
            .I(N__50454));
    Span4Mux_h I__12246 (
            .O(N__50517),
            .I(N__50449));
    LocalMux I__12245 (
            .O(N__50512),
            .I(N__50449));
    LocalMux I__12244 (
            .O(N__50509),
            .I(N__50446));
    LocalMux I__12243 (
            .O(N__50506),
            .I(N__50437));
    LocalMux I__12242 (
            .O(N__50503),
            .I(N__50437));
    Span12Mux_v I__12241 (
            .O(N__50500),
            .I(N__50437));
    InMux I__12240 (
            .O(N__50499),
            .I(N__50434));
    Span4Mux_v I__12239 (
            .O(N__50496),
            .I(N__50429));
    Span4Mux_h I__12238 (
            .O(N__50493),
            .I(N__50429));
    InMux I__12237 (
            .O(N__50492),
            .I(N__50424));
    InMux I__12236 (
            .O(N__50491),
            .I(N__50424));
    InMux I__12235 (
            .O(N__50490),
            .I(N__50421));
    LocalMux I__12234 (
            .O(N__50487),
            .I(N__50418));
    LocalMux I__12233 (
            .O(N__50482),
            .I(N__50411));
    LocalMux I__12232 (
            .O(N__50479),
            .I(N__50411));
    LocalMux I__12231 (
            .O(N__50476),
            .I(N__50411));
    LocalMux I__12230 (
            .O(N__50473),
            .I(N__50398));
    LocalMux I__12229 (
            .O(N__50470),
            .I(N__50398));
    LocalMux I__12228 (
            .O(N__50467),
            .I(N__50398));
    LocalMux I__12227 (
            .O(N__50462),
            .I(N__50398));
    Span4Mux_v I__12226 (
            .O(N__50459),
            .I(N__50398));
    Span4Mux_h I__12225 (
            .O(N__50454),
            .I(N__50398));
    Span4Mux_h I__12224 (
            .O(N__50449),
            .I(N__50393));
    Span4Mux_h I__12223 (
            .O(N__50446),
            .I(N__50393));
    InMux I__12222 (
            .O(N__50445),
            .I(N__50388));
    InMux I__12221 (
            .O(N__50444),
            .I(N__50388));
    Span12Mux_h I__12220 (
            .O(N__50437),
            .I(N__50385));
    LocalMux I__12219 (
            .O(N__50434),
            .I(N__50378));
    Span4Mux_h I__12218 (
            .O(N__50429),
            .I(N__50378));
    LocalMux I__12217 (
            .O(N__50424),
            .I(N__50378));
    LocalMux I__12216 (
            .O(N__50421),
            .I(N__50369));
    Span4Mux_h I__12215 (
            .O(N__50418),
            .I(N__50369));
    Span4Mux_v I__12214 (
            .O(N__50411),
            .I(N__50369));
    Span4Mux_h I__12213 (
            .O(N__50398),
            .I(N__50369));
    Odrv4 I__12212 (
            .O(N__50393),
            .I(current_pin_2));
    LocalMux I__12211 (
            .O(N__50388),
            .I(current_pin_2));
    Odrv12 I__12210 (
            .O(N__50385),
            .I(current_pin_2));
    Odrv4 I__12209 (
            .O(N__50378),
            .I(current_pin_2));
    Odrv4 I__12208 (
            .O(N__50369),
            .I(current_pin_2));
    CascadeMux I__12207 (
            .O(N__50358),
            .I(N__50349));
    InMux I__12206 (
            .O(N__50357),
            .I(N__50339));
    InMux I__12205 (
            .O(N__50356),
            .I(N__50329));
    InMux I__12204 (
            .O(N__50355),
            .I(N__50322));
    InMux I__12203 (
            .O(N__50354),
            .I(N__50322));
    InMux I__12202 (
            .O(N__50353),
            .I(N__50317));
    InMux I__12201 (
            .O(N__50352),
            .I(N__50317));
    InMux I__12200 (
            .O(N__50349),
            .I(N__50310));
    InMux I__12199 (
            .O(N__50348),
            .I(N__50310));
    InMux I__12198 (
            .O(N__50347),
            .I(N__50305));
    InMux I__12197 (
            .O(N__50346),
            .I(N__50305));
    InMux I__12196 (
            .O(N__50345),
            .I(N__50298));
    InMux I__12195 (
            .O(N__50344),
            .I(N__50298));
    InMux I__12194 (
            .O(N__50343),
            .I(N__50298));
    InMux I__12193 (
            .O(N__50342),
            .I(N__50295));
    LocalMux I__12192 (
            .O(N__50339),
            .I(N__50292));
    CascadeMux I__12191 (
            .O(N__50338),
            .I(N__50289));
    InMux I__12190 (
            .O(N__50337),
            .I(N__50281));
    InMux I__12189 (
            .O(N__50336),
            .I(N__50272));
    InMux I__12188 (
            .O(N__50335),
            .I(N__50272));
    InMux I__12187 (
            .O(N__50334),
            .I(N__50272));
    InMux I__12186 (
            .O(N__50333),
            .I(N__50272));
    CascadeMux I__12185 (
            .O(N__50332),
            .I(N__50269));
    LocalMux I__12184 (
            .O(N__50329),
            .I(N__50266));
    InMux I__12183 (
            .O(N__50328),
            .I(N__50257));
    InMux I__12182 (
            .O(N__50327),
            .I(N__50257));
    LocalMux I__12181 (
            .O(N__50322),
            .I(N__50253));
    LocalMux I__12180 (
            .O(N__50317),
            .I(N__50250));
    InMux I__12179 (
            .O(N__50316),
            .I(N__50247));
    InMux I__12178 (
            .O(N__50315),
            .I(N__50244));
    LocalMux I__12177 (
            .O(N__50310),
            .I(N__50241));
    LocalMux I__12176 (
            .O(N__50305),
            .I(N__50236));
    LocalMux I__12175 (
            .O(N__50298),
            .I(N__50236));
    LocalMux I__12174 (
            .O(N__50295),
            .I(N__50231));
    Span4Mux_h I__12173 (
            .O(N__50292),
            .I(N__50231));
    InMux I__12172 (
            .O(N__50289),
            .I(N__50224));
    InMux I__12171 (
            .O(N__50288),
            .I(N__50224));
    InMux I__12170 (
            .O(N__50287),
            .I(N__50224));
    InMux I__12169 (
            .O(N__50286),
            .I(N__50217));
    InMux I__12168 (
            .O(N__50285),
            .I(N__50217));
    InMux I__12167 (
            .O(N__50284),
            .I(N__50217));
    LocalMux I__12166 (
            .O(N__50281),
            .I(N__50212));
    LocalMux I__12165 (
            .O(N__50272),
            .I(N__50212));
    InMux I__12164 (
            .O(N__50269),
            .I(N__50209));
    Span12Mux_v I__12163 (
            .O(N__50266),
            .I(N__50206));
    InMux I__12162 (
            .O(N__50265),
            .I(N__50197));
    InMux I__12161 (
            .O(N__50264),
            .I(N__50197));
    InMux I__12160 (
            .O(N__50263),
            .I(N__50197));
    InMux I__12159 (
            .O(N__50262),
            .I(N__50194));
    LocalMux I__12158 (
            .O(N__50257),
            .I(N__50191));
    InMux I__12157 (
            .O(N__50256),
            .I(N__50188));
    Span4Mux_v I__12156 (
            .O(N__50253),
            .I(N__50185));
    Span4Mux_h I__12155 (
            .O(N__50250),
            .I(N__50182));
    LocalMux I__12154 (
            .O(N__50247),
            .I(N__50173));
    LocalMux I__12153 (
            .O(N__50244),
            .I(N__50173));
    Span4Mux_h I__12152 (
            .O(N__50241),
            .I(N__50173));
    Span4Mux_v I__12151 (
            .O(N__50236),
            .I(N__50173));
    Span4Mux_h I__12150 (
            .O(N__50231),
            .I(N__50164));
    LocalMux I__12149 (
            .O(N__50224),
            .I(N__50164));
    LocalMux I__12148 (
            .O(N__50217),
            .I(N__50164));
    Span4Mux_h I__12147 (
            .O(N__50212),
            .I(N__50164));
    LocalMux I__12146 (
            .O(N__50209),
            .I(N__50159));
    Span12Mux_h I__12145 (
            .O(N__50206),
            .I(N__50159));
    InMux I__12144 (
            .O(N__50205),
            .I(N__50154));
    InMux I__12143 (
            .O(N__50204),
            .I(N__50154));
    LocalMux I__12142 (
            .O(N__50197),
            .I(N__50147));
    LocalMux I__12141 (
            .O(N__50194),
            .I(N__50147));
    Span12Mux_s11_h I__12140 (
            .O(N__50191),
            .I(N__50147));
    LocalMux I__12139 (
            .O(N__50188),
            .I(current_pin_1));
    Odrv4 I__12138 (
            .O(N__50185),
            .I(current_pin_1));
    Odrv4 I__12137 (
            .O(N__50182),
            .I(current_pin_1));
    Odrv4 I__12136 (
            .O(N__50173),
            .I(current_pin_1));
    Odrv4 I__12135 (
            .O(N__50164),
            .I(current_pin_1));
    Odrv12 I__12134 (
            .O(N__50159),
            .I(current_pin_1));
    LocalMux I__12133 (
            .O(N__50154),
            .I(current_pin_1));
    Odrv12 I__12132 (
            .O(N__50147),
            .I(current_pin_1));
    InMux I__12131 (
            .O(N__50130),
            .I(N__50122));
    InMux I__12130 (
            .O(N__50129),
            .I(N__50119));
    InMux I__12129 (
            .O(N__50128),
            .I(N__50116));
    InMux I__12128 (
            .O(N__50127),
            .I(N__50113));
    InMux I__12127 (
            .O(N__50126),
            .I(N__50110));
    InMux I__12126 (
            .O(N__50125),
            .I(N__50107));
    LocalMux I__12125 (
            .O(N__50122),
            .I(N__50104));
    LocalMux I__12124 (
            .O(N__50119),
            .I(N__50099));
    LocalMux I__12123 (
            .O(N__50116),
            .I(N__50099));
    LocalMux I__12122 (
            .O(N__50113),
            .I(N__50094));
    LocalMux I__12121 (
            .O(N__50110),
            .I(N__50094));
    LocalMux I__12120 (
            .O(N__50107),
            .I(N__50089));
    Span4Mux_v I__12119 (
            .O(N__50104),
            .I(N__50089));
    Span4Mux_h I__12118 (
            .O(N__50099),
            .I(N__50086));
    Odrv12 I__12117 (
            .O(N__50094),
            .I(n9456));
    Odrv4 I__12116 (
            .O(N__50089),
            .I(n9456));
    Odrv4 I__12115 (
            .O(N__50086),
            .I(n9456));
    InMux I__12114 (
            .O(N__50079),
            .I(N__50072));
    InMux I__12113 (
            .O(N__50078),
            .I(N__50069));
    CascadeMux I__12112 (
            .O(N__50077),
            .I(N__50063));
    InMux I__12111 (
            .O(N__50076),
            .I(N__50060));
    InMux I__12110 (
            .O(N__50075),
            .I(N__50057));
    LocalMux I__12109 (
            .O(N__50072),
            .I(N__50054));
    LocalMux I__12108 (
            .O(N__50069),
            .I(N__50051));
    InMux I__12107 (
            .O(N__50068),
            .I(N__50048));
    InMux I__12106 (
            .O(N__50067),
            .I(N__50045));
    CascadeMux I__12105 (
            .O(N__50066),
            .I(N__50041));
    InMux I__12104 (
            .O(N__50063),
            .I(N__50038));
    LocalMux I__12103 (
            .O(N__50060),
            .I(N__50035));
    LocalMux I__12102 (
            .O(N__50057),
            .I(N__50031));
    Span4Mux_v I__12101 (
            .O(N__50054),
            .I(N__50028));
    Span4Mux_v I__12100 (
            .O(N__50051),
            .I(N__50023));
    LocalMux I__12099 (
            .O(N__50048),
            .I(N__50023));
    LocalMux I__12098 (
            .O(N__50045),
            .I(N__50020));
    InMux I__12097 (
            .O(N__50044),
            .I(N__50017));
    InMux I__12096 (
            .O(N__50041),
            .I(N__50011));
    LocalMux I__12095 (
            .O(N__50038),
            .I(N__50008));
    Span4Mux_v I__12094 (
            .O(N__50035),
            .I(N__50002));
    InMux I__12093 (
            .O(N__50034),
            .I(N__49996));
    Span4Mux_h I__12092 (
            .O(N__50031),
            .I(N__49993));
    Span4Mux_h I__12091 (
            .O(N__50028),
            .I(N__49990));
    Span4Mux_h I__12090 (
            .O(N__50023),
            .I(N__49987));
    Span4Mux_h I__12089 (
            .O(N__50020),
            .I(N__49979));
    LocalMux I__12088 (
            .O(N__50017),
            .I(N__49979));
    InMux I__12087 (
            .O(N__50016),
            .I(N__49974));
    InMux I__12086 (
            .O(N__50015),
            .I(N__49974));
    InMux I__12085 (
            .O(N__50014),
            .I(N__49971));
    LocalMux I__12084 (
            .O(N__50011),
            .I(N__49968));
    Span4Mux_v I__12083 (
            .O(N__50008),
            .I(N__49965));
    InMux I__12082 (
            .O(N__50007),
            .I(N__49962));
    InMux I__12081 (
            .O(N__50006),
            .I(N__49957));
    InMux I__12080 (
            .O(N__50005),
            .I(N__49957));
    Sp12to4 I__12079 (
            .O(N__50002),
            .I(N__49951));
    InMux I__12078 (
            .O(N__50001),
            .I(N__49948));
    InMux I__12077 (
            .O(N__50000),
            .I(N__49943));
    InMux I__12076 (
            .O(N__49999),
            .I(N__49943));
    LocalMux I__12075 (
            .O(N__49996),
            .I(N__49934));
    Span4Mux_v I__12074 (
            .O(N__49993),
            .I(N__49934));
    Span4Mux_h I__12073 (
            .O(N__49990),
            .I(N__49934));
    Span4Mux_v I__12072 (
            .O(N__49987),
            .I(N__49931));
    InMux I__12071 (
            .O(N__49986),
            .I(N__49924));
    InMux I__12070 (
            .O(N__49985),
            .I(N__49924));
    InMux I__12069 (
            .O(N__49984),
            .I(N__49924));
    Span4Mux_h I__12068 (
            .O(N__49979),
            .I(N__49920));
    LocalMux I__12067 (
            .O(N__49974),
            .I(N__49915));
    LocalMux I__12066 (
            .O(N__49971),
            .I(N__49915));
    Span4Mux_v I__12065 (
            .O(N__49968),
            .I(N__49906));
    Span4Mux_h I__12064 (
            .O(N__49965),
            .I(N__49906));
    LocalMux I__12063 (
            .O(N__49962),
            .I(N__49906));
    LocalMux I__12062 (
            .O(N__49957),
            .I(N__49906));
    InMux I__12061 (
            .O(N__49956),
            .I(N__49903));
    InMux I__12060 (
            .O(N__49955),
            .I(N__49898));
    InMux I__12059 (
            .O(N__49954),
            .I(N__49898));
    Span12Mux_v I__12058 (
            .O(N__49951),
            .I(N__49893));
    LocalMux I__12057 (
            .O(N__49948),
            .I(N__49893));
    LocalMux I__12056 (
            .O(N__49943),
            .I(N__49890));
    InMux I__12055 (
            .O(N__49942),
            .I(N__49885));
    InMux I__12054 (
            .O(N__49941),
            .I(N__49885));
    Span4Mux_h I__12053 (
            .O(N__49934),
            .I(N__49878));
    Span4Mux_v I__12052 (
            .O(N__49931),
            .I(N__49878));
    LocalMux I__12051 (
            .O(N__49924),
            .I(N__49878));
    InMux I__12050 (
            .O(N__49923),
            .I(N__49875));
    Span4Mux_v I__12049 (
            .O(N__49920),
            .I(N__49868));
    Span4Mux_h I__12048 (
            .O(N__49915),
            .I(N__49868));
    Span4Mux_h I__12047 (
            .O(N__49906),
            .I(N__49868));
    LocalMux I__12046 (
            .O(N__49903),
            .I(state_0));
    LocalMux I__12045 (
            .O(N__49898),
            .I(state_0));
    Odrv12 I__12044 (
            .O(N__49893),
            .I(state_0));
    Odrv12 I__12043 (
            .O(N__49890),
            .I(state_0));
    LocalMux I__12042 (
            .O(N__49885),
            .I(state_0));
    Odrv4 I__12041 (
            .O(N__49878),
            .I(state_0));
    LocalMux I__12040 (
            .O(N__49875),
            .I(state_0));
    Odrv4 I__12039 (
            .O(N__49868),
            .I(state_0));
    CascadeMux I__12038 (
            .O(N__49851),
            .I(N__49847));
    InMux I__12037 (
            .O(N__49850),
            .I(N__49844));
    InMux I__12036 (
            .O(N__49847),
            .I(N__49839));
    LocalMux I__12035 (
            .O(N__49844),
            .I(N__49835));
    InMux I__12034 (
            .O(N__49843),
            .I(N__49831));
    InMux I__12033 (
            .O(N__49842),
            .I(N__49825));
    LocalMux I__12032 (
            .O(N__49839),
            .I(N__49822));
    InMux I__12031 (
            .O(N__49838),
            .I(N__49819));
    Span4Mux_v I__12030 (
            .O(N__49835),
            .I(N__49815));
    InMux I__12029 (
            .O(N__49834),
            .I(N__49812));
    LocalMux I__12028 (
            .O(N__49831),
            .I(N__49808));
    InMux I__12027 (
            .O(N__49830),
            .I(N__49804));
    InMux I__12026 (
            .O(N__49829),
            .I(N__49800));
    CascadeMux I__12025 (
            .O(N__49828),
            .I(N__49797));
    LocalMux I__12024 (
            .O(N__49825),
            .I(N__49793));
    Span4Mux_v I__12023 (
            .O(N__49822),
            .I(N__49790));
    LocalMux I__12022 (
            .O(N__49819),
            .I(N__49787));
    InMux I__12021 (
            .O(N__49818),
            .I(N__49784));
    Span4Mux_h I__12020 (
            .O(N__49815),
            .I(N__49779));
    LocalMux I__12019 (
            .O(N__49812),
            .I(N__49779));
    CascadeMux I__12018 (
            .O(N__49811),
            .I(N__49776));
    Span4Mux_h I__12017 (
            .O(N__49808),
            .I(N__49768));
    InMux I__12016 (
            .O(N__49807),
            .I(N__49765));
    LocalMux I__12015 (
            .O(N__49804),
            .I(N__49762));
    InMux I__12014 (
            .O(N__49803),
            .I(N__49759));
    LocalMux I__12013 (
            .O(N__49800),
            .I(N__49754));
    InMux I__12012 (
            .O(N__49797),
            .I(N__49746));
    CascadeMux I__12011 (
            .O(N__49796),
            .I(N__49743));
    Span4Mux_v I__12010 (
            .O(N__49793),
            .I(N__49738));
    Span4Mux_h I__12009 (
            .O(N__49790),
            .I(N__49738));
    Span4Mux_v I__12008 (
            .O(N__49787),
            .I(N__49735));
    LocalMux I__12007 (
            .O(N__49784),
            .I(N__49730));
    Span4Mux_v I__12006 (
            .O(N__49779),
            .I(N__49730));
    InMux I__12005 (
            .O(N__49776),
            .I(N__49723));
    InMux I__12004 (
            .O(N__49775),
            .I(N__49723));
    InMux I__12003 (
            .O(N__49774),
            .I(N__49723));
    InMux I__12002 (
            .O(N__49773),
            .I(N__49719));
    CascadeMux I__12001 (
            .O(N__49772),
            .I(N__49716));
    InMux I__12000 (
            .O(N__49771),
            .I(N__49713));
    Span4Mux_h I__11999 (
            .O(N__49768),
            .I(N__49704));
    LocalMux I__11998 (
            .O(N__49765),
            .I(N__49704));
    Span4Mux_v I__11997 (
            .O(N__49762),
            .I(N__49704));
    LocalMux I__11996 (
            .O(N__49759),
            .I(N__49704));
    InMux I__11995 (
            .O(N__49758),
            .I(N__49701));
    CascadeMux I__11994 (
            .O(N__49757),
            .I(N__49698));
    Sp12to4 I__11993 (
            .O(N__49754),
            .I(N__49694));
    InMux I__11992 (
            .O(N__49753),
            .I(N__49691));
    InMux I__11991 (
            .O(N__49752),
            .I(N__49688));
    InMux I__11990 (
            .O(N__49751),
            .I(N__49685));
    InMux I__11989 (
            .O(N__49750),
            .I(N__49680));
    InMux I__11988 (
            .O(N__49749),
            .I(N__49680));
    LocalMux I__11987 (
            .O(N__49746),
            .I(N__49677));
    InMux I__11986 (
            .O(N__49743),
            .I(N__49674));
    Span4Mux_h I__11985 (
            .O(N__49738),
            .I(N__49665));
    Span4Mux_v I__11984 (
            .O(N__49735),
            .I(N__49665));
    Span4Mux_v I__11983 (
            .O(N__49730),
            .I(N__49665));
    LocalMux I__11982 (
            .O(N__49723),
            .I(N__49665));
    InMux I__11981 (
            .O(N__49722),
            .I(N__49662));
    LocalMux I__11980 (
            .O(N__49719),
            .I(N__49659));
    InMux I__11979 (
            .O(N__49716),
            .I(N__49656));
    LocalMux I__11978 (
            .O(N__49713),
            .I(N__49649));
    Span4Mux_h I__11977 (
            .O(N__49704),
            .I(N__49649));
    LocalMux I__11976 (
            .O(N__49701),
            .I(N__49649));
    InMux I__11975 (
            .O(N__49698),
            .I(N__49646));
    InMux I__11974 (
            .O(N__49697),
            .I(N__49643));
    Span12Mux_v I__11973 (
            .O(N__49694),
            .I(N__49638));
    LocalMux I__11972 (
            .O(N__49691),
            .I(N__49638));
    LocalMux I__11971 (
            .O(N__49688),
            .I(N__49633));
    LocalMux I__11970 (
            .O(N__49685),
            .I(N__49633));
    LocalMux I__11969 (
            .O(N__49680),
            .I(N__49620));
    Span4Mux_h I__11968 (
            .O(N__49677),
            .I(N__49620));
    LocalMux I__11967 (
            .O(N__49674),
            .I(N__49620));
    Span4Mux_h I__11966 (
            .O(N__49665),
            .I(N__49620));
    LocalMux I__11965 (
            .O(N__49662),
            .I(N__49620));
    Span4Mux_v I__11964 (
            .O(N__49659),
            .I(N__49620));
    LocalMux I__11963 (
            .O(N__49656),
            .I(N__49615));
    Span4Mux_v I__11962 (
            .O(N__49649),
            .I(N__49615));
    LocalMux I__11961 (
            .O(N__49646),
            .I(state_1));
    LocalMux I__11960 (
            .O(N__49643),
            .I(state_1));
    Odrv12 I__11959 (
            .O(N__49638),
            .I(state_1));
    Odrv4 I__11958 (
            .O(N__49633),
            .I(state_1));
    Odrv4 I__11957 (
            .O(N__49620),
            .I(state_1));
    Odrv4 I__11956 (
            .O(N__49615),
            .I(state_1));
    CascadeMux I__11955 (
            .O(N__49602),
            .I(N__49597));
    CascadeMux I__11954 (
            .O(N__49601),
            .I(N__49594));
    CascadeMux I__11953 (
            .O(N__49600),
            .I(N__49590));
    InMux I__11952 (
            .O(N__49597),
            .I(N__49585));
    InMux I__11951 (
            .O(N__49594),
            .I(N__49582));
    InMux I__11950 (
            .O(N__49593),
            .I(N__49577));
    InMux I__11949 (
            .O(N__49590),
            .I(N__49574));
    InMux I__11948 (
            .O(N__49589),
            .I(N__49571));
    CascadeMux I__11947 (
            .O(N__49588),
            .I(N__49567));
    LocalMux I__11946 (
            .O(N__49585),
            .I(N__49564));
    LocalMux I__11945 (
            .O(N__49582),
            .I(N__49561));
    InMux I__11944 (
            .O(N__49581),
            .I(N__49558));
    InMux I__11943 (
            .O(N__49580),
            .I(N__49555));
    LocalMux I__11942 (
            .O(N__49577),
            .I(N__49548));
    LocalMux I__11941 (
            .O(N__49574),
            .I(N__49548));
    LocalMux I__11940 (
            .O(N__49571),
            .I(N__49545));
    InMux I__11939 (
            .O(N__49570),
            .I(N__49542));
    InMux I__11938 (
            .O(N__49567),
            .I(N__49539));
    Span4Mux_v I__11937 (
            .O(N__49564),
            .I(N__49536));
    Span4Mux_v I__11936 (
            .O(N__49561),
            .I(N__49533));
    LocalMux I__11935 (
            .O(N__49558),
            .I(N__49528));
    LocalMux I__11934 (
            .O(N__49555),
            .I(N__49528));
    InMux I__11933 (
            .O(N__49554),
            .I(N__49521));
    InMux I__11932 (
            .O(N__49553),
            .I(N__49518));
    Span4Mux_v I__11931 (
            .O(N__49548),
            .I(N__49511));
    Span4Mux_v I__11930 (
            .O(N__49545),
            .I(N__49511));
    LocalMux I__11929 (
            .O(N__49542),
            .I(N__49503));
    LocalMux I__11928 (
            .O(N__49539),
            .I(N__49503));
    Sp12to4 I__11927 (
            .O(N__49536),
            .I(N__49498));
    Sp12to4 I__11926 (
            .O(N__49533),
            .I(N__49498));
    Span4Mux_v I__11925 (
            .O(N__49528),
            .I(N__49495));
    InMux I__11924 (
            .O(N__49527),
            .I(N__49490));
    InMux I__11923 (
            .O(N__49526),
            .I(N__49490));
    InMux I__11922 (
            .O(N__49525),
            .I(N__49484));
    InMux I__11921 (
            .O(N__49524),
            .I(N__49484));
    LocalMux I__11920 (
            .O(N__49521),
            .I(N__49481));
    LocalMux I__11919 (
            .O(N__49518),
            .I(N__49478));
    InMux I__11918 (
            .O(N__49517),
            .I(N__49475));
    InMux I__11917 (
            .O(N__49516),
            .I(N__49472));
    Sp12to4 I__11916 (
            .O(N__49511),
            .I(N__49469));
    InMux I__11915 (
            .O(N__49510),
            .I(N__49466));
    InMux I__11914 (
            .O(N__49509),
            .I(N__49463));
    InMux I__11913 (
            .O(N__49508),
            .I(N__49460));
    Span12Mux_h I__11912 (
            .O(N__49503),
            .I(N__49455));
    Span12Mux_h I__11911 (
            .O(N__49498),
            .I(N__49455));
    Span4Mux_h I__11910 (
            .O(N__49495),
            .I(N__49450));
    LocalMux I__11909 (
            .O(N__49490),
            .I(N__49450));
    InMux I__11908 (
            .O(N__49489),
            .I(N__49447));
    LocalMux I__11907 (
            .O(N__49484),
            .I(N__49444));
    Span4Mux_v I__11906 (
            .O(N__49481),
            .I(N__49435));
    Span4Mux_h I__11905 (
            .O(N__49478),
            .I(N__49435));
    LocalMux I__11904 (
            .O(N__49475),
            .I(N__49435));
    LocalMux I__11903 (
            .O(N__49472),
            .I(N__49435));
    Span12Mux_s11_h I__11902 (
            .O(N__49469),
            .I(N__49426));
    LocalMux I__11901 (
            .O(N__49466),
            .I(N__49426));
    LocalMux I__11900 (
            .O(N__49463),
            .I(N__49426));
    LocalMux I__11899 (
            .O(N__49460),
            .I(N__49426));
    Odrv12 I__11898 (
            .O(N__49455),
            .I(state_2));
    Odrv4 I__11897 (
            .O(N__49450),
            .I(state_2));
    LocalMux I__11896 (
            .O(N__49447),
            .I(state_2));
    Odrv4 I__11895 (
            .O(N__49444),
            .I(state_2));
    Odrv4 I__11894 (
            .O(N__49435),
            .I(state_2));
    Odrv12 I__11893 (
            .O(N__49426),
            .I(state_2));
    CascadeMux I__11892 (
            .O(N__49413),
            .I(N__49407));
    InMux I__11891 (
            .O(N__49412),
            .I(N__49403));
    InMux I__11890 (
            .O(N__49411),
            .I(N__49396));
    InMux I__11889 (
            .O(N__49410),
            .I(N__49396));
    InMux I__11888 (
            .O(N__49407),
            .I(N__49396));
    InMux I__11887 (
            .O(N__49406),
            .I(N__49393));
    LocalMux I__11886 (
            .O(N__49403),
            .I(N__49390));
    LocalMux I__11885 (
            .O(N__49396),
            .I(N__49387));
    LocalMux I__11884 (
            .O(N__49393),
            .I(N__49384));
    Span4Mux_h I__11883 (
            .O(N__49390),
            .I(N__49381));
    Span4Mux_h I__11882 (
            .O(N__49387),
            .I(N__49378));
    Span4Mux_h I__11881 (
            .O(N__49384),
            .I(N__49375));
    Odrv4 I__11880 (
            .O(N__49381),
            .I(n15_adj_721));
    Odrv4 I__11879 (
            .O(N__49378),
            .I(n15_adj_721));
    Odrv4 I__11878 (
            .O(N__49375),
            .I(n15_adj_721));
    InMux I__11877 (
            .O(N__49368),
            .I(N__49365));
    LocalMux I__11876 (
            .O(N__49365),
            .I(N__49362));
    Odrv4 I__11875 (
            .O(N__49362),
            .I(n2421));
    InMux I__11874 (
            .O(N__49359),
            .I(N__49356));
    LocalMux I__11873 (
            .O(N__49356),
            .I(N__49353));
    Odrv12 I__11872 (
            .O(N__49353),
            .I(n2373));
    CascadeMux I__11871 (
            .O(N__49350),
            .I(N__49346));
    CascadeMux I__11870 (
            .O(N__49349),
            .I(N__49343));
    InMux I__11869 (
            .O(N__49346),
            .I(N__49340));
    InMux I__11868 (
            .O(N__49343),
            .I(N__49337));
    LocalMux I__11867 (
            .O(N__49340),
            .I(N__49334));
    LocalMux I__11866 (
            .O(N__49337),
            .I(N__49331));
    Span4Mux_v I__11865 (
            .O(N__49334),
            .I(N__49326));
    Span4Mux_h I__11864 (
            .O(N__49331),
            .I(N__49326));
    Odrv4 I__11863 (
            .O(N__49326),
            .I(n11_adj_739));
    InMux I__11862 (
            .O(N__49323),
            .I(N__49320));
    LocalMux I__11861 (
            .O(N__49320),
            .I(N__49317));
    Span4Mux_h I__11860 (
            .O(N__49317),
            .I(N__49314));
    Odrv4 I__11859 (
            .O(N__49314),
            .I(n39));
    InMux I__11858 (
            .O(N__49311),
            .I(N__49308));
    LocalMux I__11857 (
            .O(N__49308),
            .I(n42));
    CascadeMux I__11856 (
            .O(N__49305),
            .I(n40_cascade_));
    InMux I__11855 (
            .O(N__49302),
            .I(N__49299));
    LocalMux I__11854 (
            .O(N__49299),
            .I(N__49296));
    Span4Mux_v I__11853 (
            .O(N__49296),
            .I(N__49293));
    Odrv4 I__11852 (
            .O(N__49293),
            .I(n41));
    InMux I__11851 (
            .O(N__49290),
            .I(N__49287));
    LocalMux I__11850 (
            .O(N__49287),
            .I(N__49284));
    Span4Mux_v I__11849 (
            .O(N__49284),
            .I(N__49280));
    InMux I__11848 (
            .O(N__49283),
            .I(N__49277));
    Sp12to4 I__11847 (
            .O(N__49280),
            .I(N__49272));
    LocalMux I__11846 (
            .O(N__49277),
            .I(N__49272));
    Span12Mux_h I__11845 (
            .O(N__49272),
            .I(N__49269));
    Span12Mux_v I__11844 (
            .O(N__49269),
            .I(N__49266));
    Odrv12 I__11843 (
            .O(N__49266),
            .I(pin_in_19));
    InMux I__11842 (
            .O(N__49263),
            .I(N__49260));
    LocalMux I__11841 (
            .O(N__49260),
            .I(N__49256));
    CascadeMux I__11840 (
            .O(N__49259),
            .I(N__49253));
    Span4Mux_v I__11839 (
            .O(N__49256),
            .I(N__49250));
    InMux I__11838 (
            .O(N__49253),
            .I(N__49247));
    Sp12to4 I__11837 (
            .O(N__49250),
            .I(N__49242));
    LocalMux I__11836 (
            .O(N__49247),
            .I(N__49242));
    Span12Mux_h I__11835 (
            .O(N__49242),
            .I(N__49239));
    Span12Mux_v I__11834 (
            .O(N__49239),
            .I(N__49236));
    Odrv12 I__11833 (
            .O(N__49236),
            .I(pin_in_18));
    CascadeMux I__11832 (
            .O(N__49233),
            .I(N__49230));
    InMux I__11831 (
            .O(N__49230),
            .I(N__49227));
    LocalMux I__11830 (
            .O(N__49227),
            .I(N__49223));
    InMux I__11829 (
            .O(N__49226),
            .I(N__49220));
    Span4Mux_h I__11828 (
            .O(N__49223),
            .I(N__49217));
    LocalMux I__11827 (
            .O(N__49220),
            .I(N__49214));
    Sp12to4 I__11826 (
            .O(N__49217),
            .I(N__49211));
    Span4Mux_v I__11825 (
            .O(N__49214),
            .I(N__49208));
    Span12Mux_v I__11824 (
            .O(N__49211),
            .I(N__49203));
    Sp12to4 I__11823 (
            .O(N__49208),
            .I(N__49203));
    Span12Mux_v I__11822 (
            .O(N__49203),
            .I(N__49200));
    Span12Mux_h I__11821 (
            .O(N__49200),
            .I(N__49197));
    Odrv12 I__11820 (
            .O(N__49197),
            .I(pin_in_16));
    CascadeMux I__11819 (
            .O(N__49194),
            .I(n13444_cascade_));
    InMux I__11818 (
            .O(N__49191),
            .I(N__49188));
    LocalMux I__11817 (
            .O(N__49188),
            .I(N__49184));
    InMux I__11816 (
            .O(N__49187),
            .I(N__49181));
    Span4Mux_v I__11815 (
            .O(N__49184),
            .I(N__49178));
    LocalMux I__11814 (
            .O(N__49181),
            .I(N__49175));
    Span4Mux_h I__11813 (
            .O(N__49178),
            .I(N__49172));
    Sp12to4 I__11812 (
            .O(N__49175),
            .I(N__49169));
    Sp12to4 I__11811 (
            .O(N__49172),
            .I(N__49166));
    Span12Mux_v I__11810 (
            .O(N__49169),
            .I(N__49163));
    Span12Mux_h I__11809 (
            .O(N__49166),
            .I(N__49160));
    Span12Mux_h I__11808 (
            .O(N__49163),
            .I(N__49157));
    Odrv12 I__11807 (
            .O(N__49160),
            .I(pin_in_17));
    Odrv12 I__11806 (
            .O(N__49157),
            .I(pin_in_17));
    InMux I__11805 (
            .O(N__49152),
            .I(N__49149));
    LocalMux I__11804 (
            .O(N__49149),
            .I(n13447));
    InMux I__11803 (
            .O(N__49146),
            .I(N__49138));
    InMux I__11802 (
            .O(N__49145),
            .I(N__49133));
    InMux I__11801 (
            .O(N__49144),
            .I(N__49133));
    InMux I__11800 (
            .O(N__49143),
            .I(N__49130));
    InMux I__11799 (
            .O(N__49142),
            .I(N__49127));
    InMux I__11798 (
            .O(N__49141),
            .I(N__49124));
    LocalMux I__11797 (
            .O(N__49138),
            .I(N__49120));
    LocalMux I__11796 (
            .O(N__49133),
            .I(N__49113));
    LocalMux I__11795 (
            .O(N__49130),
            .I(N__49113));
    LocalMux I__11794 (
            .O(N__49127),
            .I(N__49113));
    LocalMux I__11793 (
            .O(N__49124),
            .I(N__49110));
    InMux I__11792 (
            .O(N__49123),
            .I(N__49107));
    Span4Mux_v I__11791 (
            .O(N__49120),
            .I(N__49102));
    Span4Mux_v I__11790 (
            .O(N__49113),
            .I(N__49102));
    Odrv4 I__11789 (
            .O(N__49110),
            .I(n14_adj_752));
    LocalMux I__11788 (
            .O(N__49107),
            .I(n14_adj_752));
    Odrv4 I__11787 (
            .O(N__49102),
            .I(n14_adj_752));
    InMux I__11786 (
            .O(N__49095),
            .I(N__49092));
    LocalMux I__11785 (
            .O(N__49092),
            .I(N__49088));
    InMux I__11784 (
            .O(N__49091),
            .I(N__49085));
    Sp12to4 I__11783 (
            .O(N__49088),
            .I(N__49082));
    LocalMux I__11782 (
            .O(N__49085),
            .I(N__49079));
    Span12Mux_v I__11781 (
            .O(N__49082),
            .I(N__49076));
    Sp12to4 I__11780 (
            .O(N__49079),
            .I(N__49073));
    Span12Mux_h I__11779 (
            .O(N__49076),
            .I(N__49068));
    Span12Mux_v I__11778 (
            .O(N__49073),
            .I(N__49068));
    Odrv12 I__11777 (
            .O(N__49068),
            .I(pin_in_5));
    CascadeMux I__11776 (
            .O(N__49065),
            .I(n15_adj_749_cascade_));
    InMux I__11775 (
            .O(N__49062),
            .I(N__49059));
    LocalMux I__11774 (
            .O(N__49059),
            .I(n15_adj_750));
    InMux I__11773 (
            .O(N__49056),
            .I(N__49053));
    LocalMux I__11772 (
            .O(N__49053),
            .I(n37));
    CascadeMux I__11771 (
            .O(N__49050),
            .I(N__49045));
    CascadeMux I__11770 (
            .O(N__49049),
            .I(N__49037));
    CascadeMux I__11769 (
            .O(N__49048),
            .I(N__49034));
    InMux I__11768 (
            .O(N__49045),
            .I(N__49021));
    InMux I__11767 (
            .O(N__49044),
            .I(N__49021));
    InMux I__11766 (
            .O(N__49043),
            .I(N__49021));
    InMux I__11765 (
            .O(N__49042),
            .I(N__49021));
    InMux I__11764 (
            .O(N__49041),
            .I(N__49018));
    CascadeMux I__11763 (
            .O(N__49040),
            .I(N__49011));
    InMux I__11762 (
            .O(N__49037),
            .I(N__49008));
    InMux I__11761 (
            .O(N__49034),
            .I(N__49005));
    InMux I__11760 (
            .O(N__49033),
            .I(N__48989));
    InMux I__11759 (
            .O(N__49032),
            .I(N__48986));
    InMux I__11758 (
            .O(N__49031),
            .I(N__48979));
    InMux I__11757 (
            .O(N__49030),
            .I(N__48979));
    LocalMux I__11756 (
            .O(N__49021),
            .I(N__48976));
    LocalMux I__11755 (
            .O(N__49018),
            .I(N__48973));
    InMux I__11754 (
            .O(N__49017),
            .I(N__48970));
    InMux I__11753 (
            .O(N__49016),
            .I(N__48964));
    InMux I__11752 (
            .O(N__49015),
            .I(N__48961));
    InMux I__11751 (
            .O(N__49014),
            .I(N__48956));
    InMux I__11750 (
            .O(N__49011),
            .I(N__48956));
    LocalMux I__11749 (
            .O(N__49008),
            .I(N__48950));
    LocalMux I__11748 (
            .O(N__49005),
            .I(N__48950));
    InMux I__11747 (
            .O(N__49004),
            .I(N__48947));
    InMux I__11746 (
            .O(N__49003),
            .I(N__48940));
    InMux I__11745 (
            .O(N__49002),
            .I(N__48940));
    InMux I__11744 (
            .O(N__49001),
            .I(N__48940));
    InMux I__11743 (
            .O(N__49000),
            .I(N__48937));
    InMux I__11742 (
            .O(N__48999),
            .I(N__48928));
    InMux I__11741 (
            .O(N__48998),
            .I(N__48928));
    InMux I__11740 (
            .O(N__48997),
            .I(N__48928));
    InMux I__11739 (
            .O(N__48996),
            .I(N__48928));
    InMux I__11738 (
            .O(N__48995),
            .I(N__48925));
    CascadeMux I__11737 (
            .O(N__48994),
            .I(N__48922));
    InMux I__11736 (
            .O(N__48993),
            .I(N__48914));
    InMux I__11735 (
            .O(N__48992),
            .I(N__48914));
    LocalMux I__11734 (
            .O(N__48989),
            .I(N__48910));
    LocalMux I__11733 (
            .O(N__48986),
            .I(N__48907));
    InMux I__11732 (
            .O(N__48985),
            .I(N__48902));
    InMux I__11731 (
            .O(N__48984),
            .I(N__48902));
    LocalMux I__11730 (
            .O(N__48979),
            .I(N__48895));
    Span4Mux_v I__11729 (
            .O(N__48976),
            .I(N__48895));
    Span4Mux_h I__11728 (
            .O(N__48973),
            .I(N__48895));
    LocalMux I__11727 (
            .O(N__48970),
            .I(N__48891));
    InMux I__11726 (
            .O(N__48969),
            .I(N__48884));
    InMux I__11725 (
            .O(N__48968),
            .I(N__48884));
    InMux I__11724 (
            .O(N__48967),
            .I(N__48884));
    LocalMux I__11723 (
            .O(N__48964),
            .I(N__48877));
    LocalMux I__11722 (
            .O(N__48961),
            .I(N__48877));
    LocalMux I__11721 (
            .O(N__48956),
            .I(N__48877));
    InMux I__11720 (
            .O(N__48955),
            .I(N__48874));
    Span4Mux_v I__11719 (
            .O(N__48950),
            .I(N__48869));
    LocalMux I__11718 (
            .O(N__48947),
            .I(N__48869));
    LocalMux I__11717 (
            .O(N__48940),
            .I(N__48862));
    LocalMux I__11716 (
            .O(N__48937),
            .I(N__48862));
    LocalMux I__11715 (
            .O(N__48928),
            .I(N__48862));
    LocalMux I__11714 (
            .O(N__48925),
            .I(N__48859));
    InMux I__11713 (
            .O(N__48922),
            .I(N__48854));
    InMux I__11712 (
            .O(N__48921),
            .I(N__48854));
    InMux I__11711 (
            .O(N__48920),
            .I(N__48849));
    InMux I__11710 (
            .O(N__48919),
            .I(N__48849));
    LocalMux I__11709 (
            .O(N__48914),
            .I(N__48846));
    InMux I__11708 (
            .O(N__48913),
            .I(N__48839));
    Span4Mux_h I__11707 (
            .O(N__48910),
            .I(N__48836));
    Span4Mux_v I__11706 (
            .O(N__48907),
            .I(N__48829));
    LocalMux I__11705 (
            .O(N__48902),
            .I(N__48829));
    Span4Mux_h I__11704 (
            .O(N__48895),
            .I(N__48829));
    InMux I__11703 (
            .O(N__48894),
            .I(N__48826));
    Span4Mux_h I__11702 (
            .O(N__48891),
            .I(N__48819));
    LocalMux I__11701 (
            .O(N__48884),
            .I(N__48819));
    Span4Mux_h I__11700 (
            .O(N__48877),
            .I(N__48819));
    LocalMux I__11699 (
            .O(N__48874),
            .I(N__48810));
    Span4Mux_h I__11698 (
            .O(N__48869),
            .I(N__48810));
    Span4Mux_v I__11697 (
            .O(N__48862),
            .I(N__48810));
    Span4Mux_v I__11696 (
            .O(N__48859),
            .I(N__48810));
    LocalMux I__11695 (
            .O(N__48854),
            .I(N__48803));
    LocalMux I__11694 (
            .O(N__48849),
            .I(N__48803));
    Span12Mux_h I__11693 (
            .O(N__48846),
            .I(N__48803));
    InMux I__11692 (
            .O(N__48845),
            .I(N__48794));
    InMux I__11691 (
            .O(N__48844),
            .I(N__48794));
    InMux I__11690 (
            .O(N__48843),
            .I(N__48794));
    InMux I__11689 (
            .O(N__48842),
            .I(N__48794));
    LocalMux I__11688 (
            .O(N__48839),
            .I(N__48787));
    Span4Mux_h I__11687 (
            .O(N__48836),
            .I(N__48787));
    Span4Mux_h I__11686 (
            .O(N__48829),
            .I(N__48787));
    LocalMux I__11685 (
            .O(N__48826),
            .I(current_pin_0));
    Odrv4 I__11684 (
            .O(N__48819),
            .I(current_pin_0));
    Odrv4 I__11683 (
            .O(N__48810),
            .I(current_pin_0));
    Odrv12 I__11682 (
            .O(N__48803),
            .I(current_pin_0));
    LocalMux I__11681 (
            .O(N__48794),
            .I(current_pin_0));
    Odrv4 I__11680 (
            .O(N__48787),
            .I(current_pin_0));
    InMux I__11679 (
            .O(N__48774),
            .I(N__48770));
    InMux I__11678 (
            .O(N__48773),
            .I(N__48767));
    LocalMux I__11677 (
            .O(N__48770),
            .I(N__48764));
    LocalMux I__11676 (
            .O(N__48767),
            .I(N__48761));
    Span4Mux_h I__11675 (
            .O(N__48764),
            .I(N__48756));
    Span4Mux_h I__11674 (
            .O(N__48761),
            .I(N__48756));
    Span4Mux_h I__11673 (
            .O(N__48756),
            .I(N__48753));
    Sp12to4 I__11672 (
            .O(N__48753),
            .I(N__48750));
    Odrv12 I__11671 (
            .O(N__48750),
            .I(pin_in_21));
    InMux I__11670 (
            .O(N__48747),
            .I(N__48743));
    InMux I__11669 (
            .O(N__48746),
            .I(N__48740));
    LocalMux I__11668 (
            .O(N__48743),
            .I(N__48737));
    LocalMux I__11667 (
            .O(N__48740),
            .I(N__48734));
    Span4Mux_v I__11666 (
            .O(N__48737),
            .I(N__48731));
    Span4Mux_v I__11665 (
            .O(N__48734),
            .I(N__48728));
    Sp12to4 I__11664 (
            .O(N__48731),
            .I(N__48723));
    Sp12to4 I__11663 (
            .O(N__48728),
            .I(N__48723));
    Span12Mux_h I__11662 (
            .O(N__48723),
            .I(N__48720));
    Odrv12 I__11661 (
            .O(N__48720),
            .I(pin_in_20));
    InMux I__11660 (
            .O(N__48717),
            .I(N__48714));
    LocalMux I__11659 (
            .O(N__48714),
            .I(n19_adj_715));
    InMux I__11658 (
            .O(N__48711),
            .I(n10384));
    InMux I__11657 (
            .O(N__48708),
            .I(n10385));
    InMux I__11656 (
            .O(N__48705),
            .I(n10386));
    CascadeMux I__11655 (
            .O(N__48702),
            .I(N__48692));
    InMux I__11654 (
            .O(N__48701),
            .I(N__48686));
    InMux I__11653 (
            .O(N__48700),
            .I(N__48686));
    InMux I__11652 (
            .O(N__48699),
            .I(N__48683));
    InMux I__11651 (
            .O(N__48698),
            .I(N__48677));
    InMux I__11650 (
            .O(N__48697),
            .I(N__48672));
    InMux I__11649 (
            .O(N__48696),
            .I(N__48672));
    CascadeMux I__11648 (
            .O(N__48695),
            .I(N__48667));
    InMux I__11647 (
            .O(N__48692),
            .I(N__48663));
    InMux I__11646 (
            .O(N__48691),
            .I(N__48660));
    LocalMux I__11645 (
            .O(N__48686),
            .I(N__48657));
    LocalMux I__11644 (
            .O(N__48683),
            .I(N__48654));
    InMux I__11643 (
            .O(N__48682),
            .I(N__48651));
    InMux I__11642 (
            .O(N__48681),
            .I(N__48648));
    InMux I__11641 (
            .O(N__48680),
            .I(N__48642));
    LocalMux I__11640 (
            .O(N__48677),
            .I(N__48637));
    LocalMux I__11639 (
            .O(N__48672),
            .I(N__48637));
    InMux I__11638 (
            .O(N__48671),
            .I(N__48628));
    InMux I__11637 (
            .O(N__48670),
            .I(N__48628));
    InMux I__11636 (
            .O(N__48667),
            .I(N__48628));
    InMux I__11635 (
            .O(N__48666),
            .I(N__48628));
    LocalMux I__11634 (
            .O(N__48663),
            .I(N__48625));
    LocalMux I__11633 (
            .O(N__48660),
            .I(N__48620));
    Span4Mux_h I__11632 (
            .O(N__48657),
            .I(N__48620));
    Span4Mux_v I__11631 (
            .O(N__48654),
            .I(N__48613));
    LocalMux I__11630 (
            .O(N__48651),
            .I(N__48613));
    LocalMux I__11629 (
            .O(N__48648),
            .I(N__48613));
    InMux I__11628 (
            .O(N__48647),
            .I(N__48610));
    InMux I__11627 (
            .O(N__48646),
            .I(N__48607));
    InMux I__11626 (
            .O(N__48645),
            .I(N__48604));
    LocalMux I__11625 (
            .O(N__48642),
            .I(N__48597));
    Span4Mux_h I__11624 (
            .O(N__48637),
            .I(N__48597));
    LocalMux I__11623 (
            .O(N__48628),
            .I(N__48597));
    Span4Mux_h I__11622 (
            .O(N__48625),
            .I(N__48594));
    Span4Mux_h I__11621 (
            .O(N__48620),
            .I(N__48589));
    Span4Mux_h I__11620 (
            .O(N__48613),
            .I(N__48589));
    LocalMux I__11619 (
            .O(N__48610),
            .I(current_pin_4));
    LocalMux I__11618 (
            .O(N__48607),
            .I(current_pin_4));
    LocalMux I__11617 (
            .O(N__48604),
            .I(current_pin_4));
    Odrv4 I__11616 (
            .O(N__48597),
            .I(current_pin_4));
    Odrv4 I__11615 (
            .O(N__48594),
            .I(current_pin_4));
    Odrv4 I__11614 (
            .O(N__48589),
            .I(current_pin_4));
    InMux I__11613 (
            .O(N__48576),
            .I(n10387));
    InMux I__11612 (
            .O(N__48573),
            .I(N__48569));
    InMux I__11611 (
            .O(N__48572),
            .I(N__48566));
    LocalMux I__11610 (
            .O(N__48569),
            .I(N__48563));
    LocalMux I__11609 (
            .O(N__48566),
            .I(N__48560));
    Span4Mux_v I__11608 (
            .O(N__48563),
            .I(N__48554));
    Span4Mux_h I__11607 (
            .O(N__48560),
            .I(N__48554));
    InMux I__11606 (
            .O(N__48559),
            .I(N__48550));
    Span4Mux_h I__11605 (
            .O(N__48554),
            .I(N__48547));
    InMux I__11604 (
            .O(N__48553),
            .I(N__48544));
    LocalMux I__11603 (
            .O(N__48550),
            .I(current_pin_5));
    Odrv4 I__11602 (
            .O(N__48547),
            .I(current_pin_5));
    LocalMux I__11601 (
            .O(N__48544),
            .I(current_pin_5));
    InMux I__11600 (
            .O(N__48537),
            .I(n10388));
    InMux I__11599 (
            .O(N__48534),
            .I(N__48531));
    LocalMux I__11598 (
            .O(N__48531),
            .I(N__48528));
    Span4Mux_h I__11597 (
            .O(N__48528),
            .I(N__48523));
    InMux I__11596 (
            .O(N__48527),
            .I(N__48520));
    InMux I__11595 (
            .O(N__48526),
            .I(N__48516));
    Span4Mux_h I__11594 (
            .O(N__48523),
            .I(N__48513));
    LocalMux I__11593 (
            .O(N__48520),
            .I(N__48510));
    InMux I__11592 (
            .O(N__48519),
            .I(N__48507));
    LocalMux I__11591 (
            .O(N__48516),
            .I(current_pin_6));
    Odrv4 I__11590 (
            .O(N__48513),
            .I(current_pin_6));
    Odrv12 I__11589 (
            .O(N__48510),
            .I(current_pin_6));
    LocalMux I__11588 (
            .O(N__48507),
            .I(current_pin_6));
    InMux I__11587 (
            .O(N__48498),
            .I(n10389));
    InMux I__11586 (
            .O(N__48495),
            .I(n10390));
    CascadeMux I__11585 (
            .O(N__48492),
            .I(N__48489));
    InMux I__11584 (
            .O(N__48489),
            .I(N__48486));
    LocalMux I__11583 (
            .O(N__48486),
            .I(N__48483));
    Span4Mux_h I__11582 (
            .O(N__48483),
            .I(N__48478));
    InMux I__11581 (
            .O(N__48482),
            .I(N__48475));
    InMux I__11580 (
            .O(N__48481),
            .I(N__48471));
    Span4Mux_h I__11579 (
            .O(N__48478),
            .I(N__48468));
    LocalMux I__11578 (
            .O(N__48475),
            .I(N__48465));
    InMux I__11577 (
            .O(N__48474),
            .I(N__48462));
    LocalMux I__11576 (
            .O(N__48471),
            .I(current_pin_7));
    Odrv4 I__11575 (
            .O(N__48468),
            .I(current_pin_7));
    Odrv12 I__11574 (
            .O(N__48465),
            .I(current_pin_7));
    LocalMux I__11573 (
            .O(N__48462),
            .I(current_pin_7));
    ClkMux I__11572 (
            .O(N__48453),
            .I(N__48240));
    ClkMux I__11571 (
            .O(N__48452),
            .I(N__48240));
    ClkMux I__11570 (
            .O(N__48451),
            .I(N__48240));
    ClkMux I__11569 (
            .O(N__48450),
            .I(N__48240));
    ClkMux I__11568 (
            .O(N__48449),
            .I(N__48240));
    ClkMux I__11567 (
            .O(N__48448),
            .I(N__48240));
    ClkMux I__11566 (
            .O(N__48447),
            .I(N__48240));
    ClkMux I__11565 (
            .O(N__48446),
            .I(N__48240));
    ClkMux I__11564 (
            .O(N__48445),
            .I(N__48240));
    ClkMux I__11563 (
            .O(N__48444),
            .I(N__48240));
    ClkMux I__11562 (
            .O(N__48443),
            .I(N__48240));
    ClkMux I__11561 (
            .O(N__48442),
            .I(N__48240));
    ClkMux I__11560 (
            .O(N__48441),
            .I(N__48240));
    ClkMux I__11559 (
            .O(N__48440),
            .I(N__48240));
    ClkMux I__11558 (
            .O(N__48439),
            .I(N__48240));
    ClkMux I__11557 (
            .O(N__48438),
            .I(N__48240));
    ClkMux I__11556 (
            .O(N__48437),
            .I(N__48240));
    ClkMux I__11555 (
            .O(N__48436),
            .I(N__48240));
    ClkMux I__11554 (
            .O(N__48435),
            .I(N__48240));
    ClkMux I__11553 (
            .O(N__48434),
            .I(N__48240));
    ClkMux I__11552 (
            .O(N__48433),
            .I(N__48240));
    ClkMux I__11551 (
            .O(N__48432),
            .I(N__48240));
    ClkMux I__11550 (
            .O(N__48431),
            .I(N__48240));
    ClkMux I__11549 (
            .O(N__48430),
            .I(N__48240));
    ClkMux I__11548 (
            .O(N__48429),
            .I(N__48240));
    ClkMux I__11547 (
            .O(N__48428),
            .I(N__48240));
    ClkMux I__11546 (
            .O(N__48427),
            .I(N__48240));
    ClkMux I__11545 (
            .O(N__48426),
            .I(N__48240));
    ClkMux I__11544 (
            .O(N__48425),
            .I(N__48240));
    ClkMux I__11543 (
            .O(N__48424),
            .I(N__48240));
    ClkMux I__11542 (
            .O(N__48423),
            .I(N__48240));
    ClkMux I__11541 (
            .O(N__48422),
            .I(N__48240));
    ClkMux I__11540 (
            .O(N__48421),
            .I(N__48240));
    ClkMux I__11539 (
            .O(N__48420),
            .I(N__48240));
    ClkMux I__11538 (
            .O(N__48419),
            .I(N__48240));
    ClkMux I__11537 (
            .O(N__48418),
            .I(N__48240));
    ClkMux I__11536 (
            .O(N__48417),
            .I(N__48240));
    ClkMux I__11535 (
            .O(N__48416),
            .I(N__48240));
    ClkMux I__11534 (
            .O(N__48415),
            .I(N__48240));
    ClkMux I__11533 (
            .O(N__48414),
            .I(N__48240));
    ClkMux I__11532 (
            .O(N__48413),
            .I(N__48240));
    ClkMux I__11531 (
            .O(N__48412),
            .I(N__48240));
    ClkMux I__11530 (
            .O(N__48411),
            .I(N__48240));
    ClkMux I__11529 (
            .O(N__48410),
            .I(N__48240));
    ClkMux I__11528 (
            .O(N__48409),
            .I(N__48240));
    ClkMux I__11527 (
            .O(N__48408),
            .I(N__48240));
    ClkMux I__11526 (
            .O(N__48407),
            .I(N__48240));
    ClkMux I__11525 (
            .O(N__48406),
            .I(N__48240));
    ClkMux I__11524 (
            .O(N__48405),
            .I(N__48240));
    ClkMux I__11523 (
            .O(N__48404),
            .I(N__48240));
    ClkMux I__11522 (
            .O(N__48403),
            .I(N__48240));
    ClkMux I__11521 (
            .O(N__48402),
            .I(N__48240));
    ClkMux I__11520 (
            .O(N__48401),
            .I(N__48240));
    ClkMux I__11519 (
            .O(N__48400),
            .I(N__48240));
    ClkMux I__11518 (
            .O(N__48399),
            .I(N__48240));
    ClkMux I__11517 (
            .O(N__48398),
            .I(N__48240));
    ClkMux I__11516 (
            .O(N__48397),
            .I(N__48240));
    ClkMux I__11515 (
            .O(N__48396),
            .I(N__48240));
    ClkMux I__11514 (
            .O(N__48395),
            .I(N__48240));
    ClkMux I__11513 (
            .O(N__48394),
            .I(N__48240));
    ClkMux I__11512 (
            .O(N__48393),
            .I(N__48240));
    ClkMux I__11511 (
            .O(N__48392),
            .I(N__48240));
    ClkMux I__11510 (
            .O(N__48391),
            .I(N__48240));
    ClkMux I__11509 (
            .O(N__48390),
            .I(N__48240));
    ClkMux I__11508 (
            .O(N__48389),
            .I(N__48240));
    ClkMux I__11507 (
            .O(N__48388),
            .I(N__48240));
    ClkMux I__11506 (
            .O(N__48387),
            .I(N__48240));
    ClkMux I__11505 (
            .O(N__48386),
            .I(N__48240));
    ClkMux I__11504 (
            .O(N__48385),
            .I(N__48240));
    ClkMux I__11503 (
            .O(N__48384),
            .I(N__48240));
    ClkMux I__11502 (
            .O(N__48383),
            .I(N__48240));
    GlobalMux I__11501 (
            .O(N__48240),
            .I(N__48237));
    gio2CtrlBuf I__11500 (
            .O(N__48237),
            .I(CLK_c));
    CEMux I__11499 (
            .O(N__48234),
            .I(N__48230));
    InMux I__11498 (
            .O(N__48233),
            .I(N__48227));
    LocalMux I__11497 (
            .O(N__48230),
            .I(n7223));
    LocalMux I__11496 (
            .O(N__48227),
            .I(n7223));
    SRMux I__11495 (
            .O(N__48222),
            .I(N__48219));
    LocalMux I__11494 (
            .O(N__48219),
            .I(N__48216));
    Odrv4 I__11493 (
            .O(N__48216),
            .I(n7401));
    SRMux I__11492 (
            .O(N__48213),
            .I(N__48210));
    LocalMux I__11491 (
            .O(N__48210),
            .I(N__48207));
    Sp12to4 I__11490 (
            .O(N__48207),
            .I(N__48204));
    Odrv12 I__11489 (
            .O(N__48204),
            .I(n7409));
    CascadeMux I__11488 (
            .O(N__48201),
            .I(N__48198));
    InMux I__11487 (
            .O(N__48198),
            .I(N__48194));
    CascadeMux I__11486 (
            .O(N__48197),
            .I(N__48191));
    LocalMux I__11485 (
            .O(N__48194),
            .I(N__48188));
    InMux I__11484 (
            .O(N__48191),
            .I(N__48185));
    Span4Mux_h I__11483 (
            .O(N__48188),
            .I(N__48182));
    LocalMux I__11482 (
            .O(N__48185),
            .I(n11_adj_743));
    Odrv4 I__11481 (
            .O(N__48182),
            .I(n11_adj_743));
    InMux I__11480 (
            .O(N__48177),
            .I(N__48173));
    InMux I__11479 (
            .O(N__48176),
            .I(N__48170));
    LocalMux I__11478 (
            .O(N__48173),
            .I(counter_1));
    LocalMux I__11477 (
            .O(N__48170),
            .I(counter_1));
    CascadeMux I__11476 (
            .O(N__48165),
            .I(n10_adj_762_cascade_));
    InMux I__11475 (
            .O(N__48162),
            .I(N__48158));
    InMux I__11474 (
            .O(N__48161),
            .I(N__48155));
    LocalMux I__11473 (
            .O(N__48158),
            .I(counter_5));
    LocalMux I__11472 (
            .O(N__48155),
            .I(counter_5));
    InMux I__11471 (
            .O(N__48150),
            .I(N__48144));
    InMux I__11470 (
            .O(N__48149),
            .I(N__48141));
    InMux I__11469 (
            .O(N__48148),
            .I(N__48138));
    CascadeMux I__11468 (
            .O(N__48147),
            .I(N__48134));
    LocalMux I__11467 (
            .O(N__48144),
            .I(N__48129));
    LocalMux I__11466 (
            .O(N__48141),
            .I(N__48124));
    LocalMux I__11465 (
            .O(N__48138),
            .I(N__48124));
    InMux I__11464 (
            .O(N__48137),
            .I(N__48121));
    InMux I__11463 (
            .O(N__48134),
            .I(N__48116));
    InMux I__11462 (
            .O(N__48133),
            .I(N__48116));
    InMux I__11461 (
            .O(N__48132),
            .I(N__48113));
    Span4Mux_v I__11460 (
            .O(N__48129),
            .I(N__48108));
    Span4Mux_h I__11459 (
            .O(N__48124),
            .I(N__48108));
    LocalMux I__11458 (
            .O(N__48121),
            .I(N__48103));
    LocalMux I__11457 (
            .O(N__48116),
            .I(N__48103));
    LocalMux I__11456 (
            .O(N__48113),
            .I(n18_adj_742));
    Odrv4 I__11455 (
            .O(N__48108),
            .I(n18_adj_742));
    Odrv12 I__11454 (
            .O(N__48103),
            .I(n18_adj_742));
    InMux I__11453 (
            .O(N__48096),
            .I(N__48093));
    LocalMux I__11452 (
            .O(N__48093),
            .I(N__48090));
    Span4Mux_v I__11451 (
            .O(N__48090),
            .I(N__48087));
    Odrv4 I__11450 (
            .O(N__48087),
            .I(n4));
    IoInMux I__11449 (
            .O(N__48084),
            .I(N__48081));
    LocalMux I__11448 (
            .O(N__48081),
            .I(N__48078));
    IoSpan4Mux I__11447 (
            .O(N__48078),
            .I(N__48074));
    InMux I__11446 (
            .O(N__48077),
            .I(N__48070));
    Sp12to4 I__11445 (
            .O(N__48074),
            .I(N__48067));
    CascadeMux I__11444 (
            .O(N__48073),
            .I(N__48064));
    LocalMux I__11443 (
            .O(N__48070),
            .I(N__48061));
    Span12Mux_s9_h I__11442 (
            .O(N__48067),
            .I(N__48058));
    InMux I__11441 (
            .O(N__48064),
            .I(N__48055));
    Span4Mux_h I__11440 (
            .O(N__48061),
            .I(N__48052));
    Odrv12 I__11439 (
            .O(N__48058),
            .I(pin_out_13));
    LocalMux I__11438 (
            .O(N__48055),
            .I(pin_out_13));
    Odrv4 I__11437 (
            .O(N__48052),
            .I(pin_out_13));
    IoInMux I__11436 (
            .O(N__48045),
            .I(N__48042));
    LocalMux I__11435 (
            .O(N__48042),
            .I(N__48039));
    Span12Mux_s5_h I__11434 (
            .O(N__48039),
            .I(N__48035));
    InMux I__11433 (
            .O(N__48038),
            .I(N__48032));
    Span12Mux_h I__11432 (
            .O(N__48035),
            .I(N__48029));
    LocalMux I__11431 (
            .O(N__48032),
            .I(N__48025));
    Span12Mux_v I__11430 (
            .O(N__48029),
            .I(N__48022));
    InMux I__11429 (
            .O(N__48028),
            .I(N__48019));
    Span4Mux_h I__11428 (
            .O(N__48025),
            .I(N__48016));
    Odrv12 I__11427 (
            .O(N__48022),
            .I(pin_out_12));
    LocalMux I__11426 (
            .O(N__48019),
            .I(pin_out_12));
    Odrv4 I__11425 (
            .O(N__48016),
            .I(pin_out_12));
    CascadeMux I__11424 (
            .O(N__48009),
            .I(n13164_cascade_));
    InMux I__11423 (
            .O(N__48006),
            .I(N__48003));
    LocalMux I__11422 (
            .O(N__48003),
            .I(N__48000));
    Odrv4 I__11421 (
            .O(N__48000),
            .I(n13468));
    CascadeMux I__11420 (
            .O(N__47997),
            .I(N__47988));
    InMux I__11419 (
            .O(N__47996),
            .I(N__47985));
    InMux I__11418 (
            .O(N__47995),
            .I(N__47982));
    InMux I__11417 (
            .O(N__47994),
            .I(N__47978));
    InMux I__11416 (
            .O(N__47993),
            .I(N__47975));
    InMux I__11415 (
            .O(N__47992),
            .I(N__47970));
    InMux I__11414 (
            .O(N__47991),
            .I(N__47970));
    InMux I__11413 (
            .O(N__47988),
            .I(N__47967));
    LocalMux I__11412 (
            .O(N__47985),
            .I(N__47964));
    LocalMux I__11411 (
            .O(N__47982),
            .I(N__47961));
    InMux I__11410 (
            .O(N__47981),
            .I(N__47958));
    LocalMux I__11409 (
            .O(N__47978),
            .I(N__47955));
    LocalMux I__11408 (
            .O(N__47975),
            .I(N__47950));
    LocalMux I__11407 (
            .O(N__47970),
            .I(N__47950));
    LocalMux I__11406 (
            .O(N__47967),
            .I(N__47945));
    Span4Mux_v I__11405 (
            .O(N__47964),
            .I(N__47945));
    Span12Mux_v I__11404 (
            .O(N__47961),
            .I(N__47940));
    LocalMux I__11403 (
            .O(N__47958),
            .I(N__47940));
    Span4Mux_h I__11402 (
            .O(N__47955),
            .I(N__47935));
    Span4Mux_h I__11401 (
            .O(N__47950),
            .I(N__47935));
    Odrv4 I__11400 (
            .O(N__47945),
            .I(n6_adj_748));
    Odrv12 I__11399 (
            .O(N__47940),
            .I(n6_adj_748));
    Odrv4 I__11398 (
            .O(N__47935),
            .I(n6_adj_748));
    InMux I__11397 (
            .O(N__47928),
            .I(N__47924));
    CascadeMux I__11396 (
            .O(N__47927),
            .I(N__47921));
    LocalMux I__11395 (
            .O(N__47924),
            .I(N__47918));
    InMux I__11394 (
            .O(N__47921),
            .I(N__47915));
    Span4Mux_v I__11393 (
            .O(N__47918),
            .I(N__47912));
    LocalMux I__11392 (
            .O(N__47915),
            .I(N__47909));
    Sp12to4 I__11391 (
            .O(N__47912),
            .I(N__47906));
    Span4Mux_h I__11390 (
            .O(N__47909),
            .I(N__47903));
    Span12Mux_h I__11389 (
            .O(N__47906),
            .I(N__47900));
    Span4Mux_h I__11388 (
            .O(N__47903),
            .I(N__47897));
    Span12Mux_v I__11387 (
            .O(N__47900),
            .I(N__47894));
    Sp12to4 I__11386 (
            .O(N__47897),
            .I(N__47891));
    Odrv12 I__11385 (
            .O(N__47894),
            .I(pin_in_22));
    Odrv12 I__11384 (
            .O(N__47891),
            .I(pin_in_22));
    CascadeMux I__11383 (
            .O(N__47886),
            .I(n6_adj_748_cascade_));
    InMux I__11382 (
            .O(N__47883),
            .I(N__47879));
    IoInMux I__11381 (
            .O(N__47882),
            .I(N__47876));
    LocalMux I__11380 (
            .O(N__47879),
            .I(N__47873));
    LocalMux I__11379 (
            .O(N__47876),
            .I(N__47870));
    Span4Mux_h I__11378 (
            .O(N__47873),
            .I(N__47866));
    Span12Mux_s6_h I__11377 (
            .O(N__47870),
            .I(N__47863));
    InMux I__11376 (
            .O(N__47869),
            .I(N__47860));
    Span4Mux_v I__11375 (
            .O(N__47866),
            .I(N__47857));
    Odrv12 I__11374 (
            .O(N__47863),
            .I(pin_out_15));
    LocalMux I__11373 (
            .O(N__47860),
            .I(pin_out_15));
    Odrv4 I__11372 (
            .O(N__47857),
            .I(pin_out_15));
    IoInMux I__11371 (
            .O(N__47850),
            .I(N__47847));
    LocalMux I__11370 (
            .O(N__47847),
            .I(N__47844));
    Span12Mux_s5_h I__11369 (
            .O(N__47844),
            .I(N__47840));
    InMux I__11368 (
            .O(N__47843),
            .I(N__47836));
    Span12Mux_h I__11367 (
            .O(N__47840),
            .I(N__47833));
    InMux I__11366 (
            .O(N__47839),
            .I(N__47830));
    LocalMux I__11365 (
            .O(N__47836),
            .I(N__47827));
    Odrv12 I__11364 (
            .O(N__47833),
            .I(pin_out_14));
    LocalMux I__11363 (
            .O(N__47830),
            .I(pin_out_14));
    Odrv4 I__11362 (
            .O(N__47827),
            .I(pin_out_14));
    InMux I__11361 (
            .O(N__47820),
            .I(N__47817));
    LocalMux I__11360 (
            .O(N__47817),
            .I(n13165));
    InMux I__11359 (
            .O(N__47814),
            .I(bfn_17_17_0_));
    CascadeMux I__11358 (
            .O(N__47811),
            .I(n13144_cascade_));
    InMux I__11357 (
            .O(N__47808),
            .I(N__47805));
    LocalMux I__11356 (
            .O(N__47805),
            .I(N__47802));
    Odrv4 I__11355 (
            .O(N__47802),
            .I(n13279));
    InMux I__11354 (
            .O(N__47799),
            .I(N__47792));
    InMux I__11353 (
            .O(N__47798),
            .I(N__47789));
    InMux I__11352 (
            .O(N__47797),
            .I(N__47784));
    InMux I__11351 (
            .O(N__47796),
            .I(N__47784));
    InMux I__11350 (
            .O(N__47795),
            .I(N__47781));
    LocalMux I__11349 (
            .O(N__47792),
            .I(N__47775));
    LocalMux I__11348 (
            .O(N__47789),
            .I(N__47770));
    LocalMux I__11347 (
            .O(N__47784),
            .I(N__47770));
    LocalMux I__11346 (
            .O(N__47781),
            .I(N__47767));
    InMux I__11345 (
            .O(N__47780),
            .I(N__47760));
    InMux I__11344 (
            .O(N__47779),
            .I(N__47760));
    InMux I__11343 (
            .O(N__47778),
            .I(N__47760));
    Span4Mux_h I__11342 (
            .O(N__47775),
            .I(N__47757));
    Span4Mux_h I__11341 (
            .O(N__47770),
            .I(N__47754));
    Span4Mux_h I__11340 (
            .O(N__47767),
            .I(N__47749));
    LocalMux I__11339 (
            .O(N__47760),
            .I(N__47749));
    Odrv4 I__11338 (
            .O(N__47757),
            .I(n14_adj_717));
    Odrv4 I__11337 (
            .O(N__47754),
            .I(n14_adj_717));
    Odrv4 I__11336 (
            .O(N__47749),
            .I(n14_adj_717));
    InMux I__11335 (
            .O(N__47742),
            .I(N__47738));
    InMux I__11334 (
            .O(N__47741),
            .I(N__47735));
    LocalMux I__11333 (
            .O(N__47738),
            .I(N__47732));
    LocalMux I__11332 (
            .O(N__47735),
            .I(n11));
    Odrv4 I__11331 (
            .O(N__47732),
            .I(n11));
    InMux I__11330 (
            .O(N__47727),
            .I(N__47724));
    LocalMux I__11329 (
            .O(N__47724),
            .I(N__47721));
    Odrv12 I__11328 (
            .O(N__47721),
            .I(n30));
    InMux I__11327 (
            .O(N__47718),
            .I(N__47715));
    LocalMux I__11326 (
            .O(N__47715),
            .I(N__47712));
    Span4Mux_v I__11325 (
            .O(N__47712),
            .I(N__47708));
    InMux I__11324 (
            .O(N__47711),
            .I(N__47704));
    Span4Mux_v I__11323 (
            .O(N__47708),
            .I(N__47701));
    InMux I__11322 (
            .O(N__47707),
            .I(N__47698));
    LocalMux I__11321 (
            .O(N__47704),
            .I(N__47695));
    Span4Mux_h I__11320 (
            .O(N__47701),
            .I(N__47692));
    LocalMux I__11319 (
            .O(N__47698),
            .I(delay_counter_31));
    Odrv12 I__11318 (
            .O(N__47695),
            .I(delay_counter_31));
    Odrv4 I__11317 (
            .O(N__47692),
            .I(delay_counter_31));
    InMux I__11316 (
            .O(N__47685),
            .I(N__47682));
    LocalMux I__11315 (
            .O(N__47682),
            .I(N__47679));
    Span4Mux_v I__11314 (
            .O(N__47679),
            .I(N__47675));
    InMux I__11313 (
            .O(N__47678),
            .I(N__47672));
    Span4Mux_h I__11312 (
            .O(N__47675),
            .I(N__47669));
    LocalMux I__11311 (
            .O(N__47672),
            .I(n11612));
    Odrv4 I__11310 (
            .O(N__47669),
            .I(n11612));
    CascadeMux I__11309 (
            .O(N__47664),
            .I(N__47661));
    InMux I__11308 (
            .O(N__47661),
            .I(N__47658));
    LocalMux I__11307 (
            .O(N__47658),
            .I(N__47655));
    Span12Mux_h I__11306 (
            .O(N__47655),
            .I(N__47651));
    InMux I__11305 (
            .O(N__47654),
            .I(N__47648));
    Odrv12 I__11304 (
            .O(N__47651),
            .I(n11481));
    LocalMux I__11303 (
            .O(N__47648),
            .I(n11481));
    InMux I__11302 (
            .O(N__47643),
            .I(N__47640));
    LocalMux I__11301 (
            .O(N__47640),
            .I(N__47637));
    Span4Mux_v I__11300 (
            .O(N__47637),
            .I(N__47634));
    Odrv4 I__11299 (
            .O(N__47634),
            .I(n13273));
    InMux I__11298 (
            .O(N__47631),
            .I(N__47627));
    CascadeMux I__11297 (
            .O(N__47630),
            .I(N__47624));
    LocalMux I__11296 (
            .O(N__47627),
            .I(N__47621));
    InMux I__11295 (
            .O(N__47624),
            .I(N__47618));
    Span4Mux_v I__11294 (
            .O(N__47621),
            .I(N__47612));
    LocalMux I__11293 (
            .O(N__47618),
            .I(N__47612));
    InMux I__11292 (
            .O(N__47617),
            .I(N__47609));
    Span4Mux_v I__11291 (
            .O(N__47612),
            .I(N__47604));
    LocalMux I__11290 (
            .O(N__47609),
            .I(N__47604));
    Span4Mux_h I__11289 (
            .O(N__47604),
            .I(N__47601));
    Odrv4 I__11288 (
            .O(N__47601),
            .I(state_7_N_167_0));
    InMux I__11287 (
            .O(N__47598),
            .I(N__47594));
    InMux I__11286 (
            .O(N__47597),
            .I(N__47591));
    LocalMux I__11285 (
            .O(N__47594),
            .I(counter_3));
    LocalMux I__11284 (
            .O(N__47591),
            .I(counter_3));
    CascadeMux I__11283 (
            .O(N__47586),
            .I(N__47583));
    InMux I__11282 (
            .O(N__47583),
            .I(N__47579));
    InMux I__11281 (
            .O(N__47582),
            .I(N__47576));
    LocalMux I__11280 (
            .O(N__47579),
            .I(counter_4));
    LocalMux I__11279 (
            .O(N__47576),
            .I(counter_4));
    CascadeMux I__11278 (
            .O(N__47571),
            .I(N__47567));
    InMux I__11277 (
            .O(N__47570),
            .I(N__47564));
    InMux I__11276 (
            .O(N__47567),
            .I(N__47561));
    LocalMux I__11275 (
            .O(N__47564),
            .I(counter_0));
    LocalMux I__11274 (
            .O(N__47561),
            .I(counter_0));
    CascadeMux I__11273 (
            .O(N__47556),
            .I(N__47553));
    InMux I__11272 (
            .O(N__47553),
            .I(N__47550));
    LocalMux I__11271 (
            .O(N__47550),
            .I(N__47546));
    InMux I__11270 (
            .O(N__47549),
            .I(N__47543));
    Odrv4 I__11269 (
            .O(N__47546),
            .I(counter_2));
    LocalMux I__11268 (
            .O(N__47543),
            .I(counter_2));
    CEMux I__11267 (
            .O(N__47538),
            .I(N__47535));
    LocalMux I__11266 (
            .O(N__47535),
            .I(N__47531));
    CascadeMux I__11265 (
            .O(N__47534),
            .I(N__47520));
    Span4Mux_v I__11264 (
            .O(N__47531),
            .I(N__47515));
    CEMux I__11263 (
            .O(N__47530),
            .I(N__47512));
    InMux I__11262 (
            .O(N__47529),
            .I(N__47507));
    InMux I__11261 (
            .O(N__47528),
            .I(N__47507));
    CascadeMux I__11260 (
            .O(N__47527),
            .I(N__47498));
    InMux I__11259 (
            .O(N__47526),
            .I(N__47490));
    InMux I__11258 (
            .O(N__47525),
            .I(N__47487));
    InMux I__11257 (
            .O(N__47524),
            .I(N__47484));
    InMux I__11256 (
            .O(N__47523),
            .I(N__47477));
    InMux I__11255 (
            .O(N__47520),
            .I(N__47477));
    InMux I__11254 (
            .O(N__47519),
            .I(N__47477));
    InMux I__11253 (
            .O(N__47518),
            .I(N__47473));
    Span4Mux_v I__11252 (
            .O(N__47515),
            .I(N__47468));
    LocalMux I__11251 (
            .O(N__47512),
            .I(N__47468));
    LocalMux I__11250 (
            .O(N__47507),
            .I(N__47465));
    InMux I__11249 (
            .O(N__47506),
            .I(N__47462));
    InMux I__11248 (
            .O(N__47505),
            .I(N__47459));
    InMux I__11247 (
            .O(N__47504),
            .I(N__47455));
    InMux I__11246 (
            .O(N__47503),
            .I(N__47448));
    InMux I__11245 (
            .O(N__47502),
            .I(N__47448));
    InMux I__11244 (
            .O(N__47501),
            .I(N__47448));
    InMux I__11243 (
            .O(N__47498),
            .I(N__47445));
    InMux I__11242 (
            .O(N__47497),
            .I(N__47442));
    InMux I__11241 (
            .O(N__47496),
            .I(N__47437));
    InMux I__11240 (
            .O(N__47495),
            .I(N__47437));
    InMux I__11239 (
            .O(N__47494),
            .I(N__47432));
    InMux I__11238 (
            .O(N__47493),
            .I(N__47432));
    LocalMux I__11237 (
            .O(N__47490),
            .I(N__47423));
    LocalMux I__11236 (
            .O(N__47487),
            .I(N__47423));
    LocalMux I__11235 (
            .O(N__47484),
            .I(N__47423));
    LocalMux I__11234 (
            .O(N__47477),
            .I(N__47423));
    InMux I__11233 (
            .O(N__47476),
            .I(N__47419));
    LocalMux I__11232 (
            .O(N__47473),
            .I(N__47416));
    Span4Mux_v I__11231 (
            .O(N__47468),
            .I(N__47409));
    Span4Mux_h I__11230 (
            .O(N__47465),
            .I(N__47409));
    LocalMux I__11229 (
            .O(N__47462),
            .I(N__47409));
    LocalMux I__11228 (
            .O(N__47459),
            .I(N__47406));
    InMux I__11227 (
            .O(N__47458),
            .I(N__47403));
    LocalMux I__11226 (
            .O(N__47455),
            .I(N__47398));
    LocalMux I__11225 (
            .O(N__47448),
            .I(N__47398));
    LocalMux I__11224 (
            .O(N__47445),
            .I(N__47395));
    LocalMux I__11223 (
            .O(N__47442),
            .I(N__47390));
    LocalMux I__11222 (
            .O(N__47437),
            .I(N__47390));
    LocalMux I__11221 (
            .O(N__47432),
            .I(N__47385));
    Span4Mux_v I__11220 (
            .O(N__47423),
            .I(N__47385));
    InMux I__11219 (
            .O(N__47422),
            .I(N__47382));
    LocalMux I__11218 (
            .O(N__47419),
            .I(N__47379));
    Span4Mux_h I__11217 (
            .O(N__47416),
            .I(N__47374));
    Span4Mux_h I__11216 (
            .O(N__47409),
            .I(N__47374));
    Span4Mux_v I__11215 (
            .O(N__47406),
            .I(N__47369));
    LocalMux I__11214 (
            .O(N__47403),
            .I(N__47369));
    Span4Mux_v I__11213 (
            .O(N__47398),
            .I(N__47366));
    Span4Mux_v I__11212 (
            .O(N__47395),
            .I(N__47359));
    Span4Mux_v I__11211 (
            .O(N__47390),
            .I(N__47359));
    Span4Mux_h I__11210 (
            .O(N__47385),
            .I(N__47359));
    LocalMux I__11209 (
            .O(N__47382),
            .I(n7231));
    Odrv4 I__11208 (
            .O(N__47379),
            .I(n7231));
    Odrv4 I__11207 (
            .O(N__47374),
            .I(n7231));
    Odrv4 I__11206 (
            .O(N__47369),
            .I(n7231));
    Odrv4 I__11205 (
            .O(N__47366),
            .I(n7231));
    Odrv4 I__11204 (
            .O(N__47359),
            .I(n7231));
    InMux I__11203 (
            .O(N__47346),
            .I(N__47343));
    LocalMux I__11202 (
            .O(N__47343),
            .I(n12208));
    CascadeMux I__11201 (
            .O(N__47340),
            .I(n7500_cascade_));
    IoInMux I__11200 (
            .O(N__47337),
            .I(N__47334));
    LocalMux I__11199 (
            .O(N__47334),
            .I(N__47331));
    Span4Mux_s3_v I__11198 (
            .O(N__47331),
            .I(N__47328));
    Sp12to4 I__11197 (
            .O(N__47328),
            .I(N__47325));
    Span12Mux_h I__11196 (
            .O(N__47325),
            .I(N__47320));
    CascadeMux I__11195 (
            .O(N__47324),
            .I(N__47317));
    InMux I__11194 (
            .O(N__47323),
            .I(N__47314));
    Span12Mux_v I__11193 (
            .O(N__47320),
            .I(N__47311));
    InMux I__11192 (
            .O(N__47317),
            .I(N__47308));
    LocalMux I__11191 (
            .O(N__47314),
            .I(N__47305));
    Odrv12 I__11190 (
            .O(N__47311),
            .I(pin_out_22));
    LocalMux I__11189 (
            .O(N__47308),
            .I(pin_out_22));
    Odrv4 I__11188 (
            .O(N__47305),
            .I(pin_out_22));
    InMux I__11187 (
            .O(N__47298),
            .I(N__47295));
    LocalMux I__11186 (
            .O(N__47295),
            .I(N__47291));
    InMux I__11185 (
            .O(N__47294),
            .I(N__47287));
    Span4Mux_v I__11184 (
            .O(N__47291),
            .I(N__47284));
    InMux I__11183 (
            .O(N__47290),
            .I(N__47281));
    LocalMux I__11182 (
            .O(N__47287),
            .I(N__47278));
    Odrv4 I__11181 (
            .O(N__47284),
            .I(n8_adj_723));
    LocalMux I__11180 (
            .O(N__47281),
            .I(n8_adj_723));
    Odrv4 I__11179 (
            .O(N__47278),
            .I(n8_adj_723));
    InMux I__11178 (
            .O(N__47271),
            .I(N__47268));
    LocalMux I__11177 (
            .O(N__47268),
            .I(n4_adj_778));
    InMux I__11176 (
            .O(N__47265),
            .I(N__47260));
    InMux I__11175 (
            .O(N__47264),
            .I(N__47255));
    InMux I__11174 (
            .O(N__47263),
            .I(N__47255));
    LocalMux I__11173 (
            .O(N__47260),
            .I(N__47252));
    LocalMux I__11172 (
            .O(N__47255),
            .I(N__47249));
    Span4Mux_h I__11171 (
            .O(N__47252),
            .I(N__47246));
    Odrv4 I__11170 (
            .O(N__47249),
            .I(n7142));
    Odrv4 I__11169 (
            .O(N__47246),
            .I(n7142));
    CascadeMux I__11168 (
            .O(N__47241),
            .I(n7142_cascade_));
    InMux I__11167 (
            .O(N__47238),
            .I(N__47232));
    InMux I__11166 (
            .O(N__47237),
            .I(N__47226));
    InMux I__11165 (
            .O(N__47236),
            .I(N__47220));
    InMux I__11164 (
            .O(N__47235),
            .I(N__47220));
    LocalMux I__11163 (
            .O(N__47232),
            .I(N__47217));
    InMux I__11162 (
            .O(N__47231),
            .I(N__47212));
    InMux I__11161 (
            .O(N__47230),
            .I(N__47212));
    InMux I__11160 (
            .O(N__47229),
            .I(N__47209));
    LocalMux I__11159 (
            .O(N__47226),
            .I(N__47206));
    InMux I__11158 (
            .O(N__47225),
            .I(N__47203));
    LocalMux I__11157 (
            .O(N__47220),
            .I(N__47200));
    Span4Mux_h I__11156 (
            .O(N__47217),
            .I(N__47197));
    LocalMux I__11155 (
            .O(N__47212),
            .I(N__47194));
    LocalMux I__11154 (
            .O(N__47209),
            .I(counter_7));
    Odrv4 I__11153 (
            .O(N__47206),
            .I(counter_7));
    LocalMux I__11152 (
            .O(N__47203),
            .I(counter_7));
    Odrv4 I__11151 (
            .O(N__47200),
            .I(counter_7));
    Odrv4 I__11150 (
            .O(N__47197),
            .I(counter_7));
    Odrv12 I__11149 (
            .O(N__47194),
            .I(counter_7));
    CascadeMux I__11148 (
            .O(N__47181),
            .I(N__47177));
    CascadeMux I__11147 (
            .O(N__47180),
            .I(N__47173));
    InMux I__11146 (
            .O(N__47177),
            .I(N__47169));
    CascadeMux I__11145 (
            .O(N__47176),
            .I(N__47165));
    InMux I__11144 (
            .O(N__47173),
            .I(N__47160));
    CascadeMux I__11143 (
            .O(N__47172),
            .I(N__47157));
    LocalMux I__11142 (
            .O(N__47169),
            .I(N__47153));
    InMux I__11141 (
            .O(N__47168),
            .I(N__47148));
    InMux I__11140 (
            .O(N__47165),
            .I(N__47148));
    InMux I__11139 (
            .O(N__47164),
            .I(N__47143));
    InMux I__11138 (
            .O(N__47163),
            .I(N__47143));
    LocalMux I__11137 (
            .O(N__47160),
            .I(N__47140));
    InMux I__11136 (
            .O(N__47157),
            .I(N__47137));
    InMux I__11135 (
            .O(N__47156),
            .I(N__47134));
    Span4Mux_v I__11134 (
            .O(N__47153),
            .I(N__47129));
    LocalMux I__11133 (
            .O(N__47148),
            .I(N__47129));
    LocalMux I__11132 (
            .O(N__47143),
            .I(N__47126));
    Odrv4 I__11131 (
            .O(N__47140),
            .I(counter_6));
    LocalMux I__11130 (
            .O(N__47137),
            .I(counter_6));
    LocalMux I__11129 (
            .O(N__47134),
            .I(counter_6));
    Odrv4 I__11128 (
            .O(N__47129),
            .I(counter_6));
    Odrv12 I__11127 (
            .O(N__47126),
            .I(counter_6));
    SRMux I__11126 (
            .O(N__47115),
            .I(N__47112));
    LocalMux I__11125 (
            .O(N__47112),
            .I(N__47109));
    Span4Mux_v I__11124 (
            .O(N__47109),
            .I(N__47106));
    Sp12to4 I__11123 (
            .O(N__47106),
            .I(N__47102));
    InMux I__11122 (
            .O(N__47105),
            .I(N__47099));
    Span12Mux_s6_h I__11121 (
            .O(N__47102),
            .I(N__47096));
    LocalMux I__11120 (
            .O(N__47099),
            .I(N__47093));
    Odrv12 I__11119 (
            .O(N__47096),
            .I(n73));
    Odrv12 I__11118 (
            .O(N__47093),
            .I(n73));
    InMux I__11117 (
            .O(N__47088),
            .I(N__47085));
    LocalMux I__11116 (
            .O(N__47085),
            .I(N__47081));
    InMux I__11115 (
            .O(N__47084),
            .I(N__47078));
    Span4Mux_v I__11114 (
            .O(N__47081),
            .I(N__47075));
    LocalMux I__11113 (
            .O(N__47078),
            .I(N__47072));
    Span4Mux_v I__11112 (
            .O(N__47075),
            .I(N__47069));
    Span4Mux_v I__11111 (
            .O(N__47072),
            .I(N__47066));
    Span4Mux_v I__11110 (
            .O(N__47069),
            .I(N__47063));
    Span4Mux_v I__11109 (
            .O(N__47066),
            .I(N__47060));
    Sp12to4 I__11108 (
            .O(N__47063),
            .I(N__47057));
    Span4Mux_v I__11107 (
            .O(N__47060),
            .I(N__47054));
    Span12Mux_h I__11106 (
            .O(N__47057),
            .I(N__47051));
    Span4Mux_h I__11105 (
            .O(N__47054),
            .I(N__47048));
    Odrv12 I__11104 (
            .O(N__47051),
            .I(pin_in_7));
    Odrv4 I__11103 (
            .O(N__47048),
            .I(pin_in_7));
    InMux I__11102 (
            .O(N__47043),
            .I(N__47040));
    LocalMux I__11101 (
            .O(N__47040),
            .I(n2385));
    CascadeMux I__11100 (
            .O(N__47037),
            .I(n12123_cascade_));
    InMux I__11099 (
            .O(N__47034),
            .I(N__47031));
    LocalMux I__11098 (
            .O(N__47031),
            .I(N__47028));
    Span4Mux_v I__11097 (
            .O(N__47028),
            .I(N__47025));
    Odrv4 I__11096 (
            .O(N__47025),
            .I(n48_adj_771));
    InMux I__11095 (
            .O(N__47022),
            .I(N__47019));
    LocalMux I__11094 (
            .O(N__47019),
            .I(N__47016));
    Span4Mux_v I__11093 (
            .O(N__47016),
            .I(N__47012));
    InMux I__11092 (
            .O(N__47015),
            .I(N__47009));
    Sp12to4 I__11091 (
            .O(N__47012),
            .I(N__47006));
    LocalMux I__11090 (
            .O(N__47009),
            .I(N__47003));
    Span12Mux_h I__11089 (
            .O(N__47006),
            .I(N__46998));
    Span12Mux_s7_h I__11088 (
            .O(N__47003),
            .I(N__46998));
    Span12Mux_v I__11087 (
            .O(N__46998),
            .I(N__46995));
    Odrv12 I__11086 (
            .O(N__46995),
            .I(pin_in_4));
    InMux I__11085 (
            .O(N__46992),
            .I(N__46989));
    LocalMux I__11084 (
            .O(N__46989),
            .I(n2313));
    InMux I__11083 (
            .O(N__46986),
            .I(n10516));
    CascadeMux I__11082 (
            .O(N__46983),
            .I(n8_adj_763_cascade_));
    InMux I__11081 (
            .O(N__46980),
            .I(N__46974));
    CascadeMux I__11080 (
            .O(N__46979),
            .I(N__46971));
    CascadeMux I__11079 (
            .O(N__46978),
            .I(N__46966));
    InMux I__11078 (
            .O(N__46977),
            .I(N__46960));
    LocalMux I__11077 (
            .O(N__46974),
            .I(N__46955));
    InMux I__11076 (
            .O(N__46971),
            .I(N__46950));
    InMux I__11075 (
            .O(N__46970),
            .I(N__46950));
    InMux I__11074 (
            .O(N__46969),
            .I(N__46945));
    InMux I__11073 (
            .O(N__46966),
            .I(N__46945));
    InMux I__11072 (
            .O(N__46965),
            .I(N__46937));
    InMux I__11071 (
            .O(N__46964),
            .I(N__46932));
    InMux I__11070 (
            .O(N__46963),
            .I(N__46932));
    LocalMux I__11069 (
            .O(N__46960),
            .I(N__46924));
    CascadeMux I__11068 (
            .O(N__46959),
            .I(N__46920));
    CascadeMux I__11067 (
            .O(N__46958),
            .I(N__46917));
    Span4Mux_v I__11066 (
            .O(N__46955),
            .I(N__46908));
    LocalMux I__11065 (
            .O(N__46950),
            .I(N__46908));
    LocalMux I__11064 (
            .O(N__46945),
            .I(N__46908));
    InMux I__11063 (
            .O(N__46944),
            .I(N__46905));
    InMux I__11062 (
            .O(N__46943),
            .I(N__46898));
    InMux I__11061 (
            .O(N__46942),
            .I(N__46898));
    InMux I__11060 (
            .O(N__46941),
            .I(N__46898));
    InMux I__11059 (
            .O(N__46940),
            .I(N__46895));
    LocalMux I__11058 (
            .O(N__46937),
            .I(N__46890));
    LocalMux I__11057 (
            .O(N__46932),
            .I(N__46890));
    CascadeMux I__11056 (
            .O(N__46931),
            .I(N__46887));
    CascadeMux I__11055 (
            .O(N__46930),
            .I(N__46883));
    CascadeMux I__11054 (
            .O(N__46929),
            .I(N__46879));
    CascadeMux I__11053 (
            .O(N__46928),
            .I(N__46875));
    CascadeMux I__11052 (
            .O(N__46927),
            .I(N__46872));
    Sp12to4 I__11051 (
            .O(N__46924),
            .I(N__46868));
    InMux I__11050 (
            .O(N__46923),
            .I(N__46865));
    InMux I__11049 (
            .O(N__46920),
            .I(N__46862));
    InMux I__11048 (
            .O(N__46917),
            .I(N__46859));
    InMux I__11047 (
            .O(N__46916),
            .I(N__46856));
    InMux I__11046 (
            .O(N__46915),
            .I(N__46853));
    Span4Mux_v I__11045 (
            .O(N__46908),
            .I(N__46850));
    LocalMux I__11044 (
            .O(N__46905),
            .I(N__46841));
    LocalMux I__11043 (
            .O(N__46898),
            .I(N__46841));
    LocalMux I__11042 (
            .O(N__46895),
            .I(N__46841));
    Span4Mux_h I__11041 (
            .O(N__46890),
            .I(N__46841));
    InMux I__11040 (
            .O(N__46887),
            .I(N__46826));
    InMux I__11039 (
            .O(N__46886),
            .I(N__46826));
    InMux I__11038 (
            .O(N__46883),
            .I(N__46826));
    InMux I__11037 (
            .O(N__46882),
            .I(N__46826));
    InMux I__11036 (
            .O(N__46879),
            .I(N__46826));
    InMux I__11035 (
            .O(N__46878),
            .I(N__46826));
    InMux I__11034 (
            .O(N__46875),
            .I(N__46826));
    InMux I__11033 (
            .O(N__46872),
            .I(N__46821));
    InMux I__11032 (
            .O(N__46871),
            .I(N__46821));
    Span12Mux_v I__11031 (
            .O(N__46868),
            .I(N__46818));
    LocalMux I__11030 (
            .O(N__46865),
            .I(N__46807));
    LocalMux I__11029 (
            .O(N__46862),
            .I(N__46807));
    LocalMux I__11028 (
            .O(N__46859),
            .I(N__46807));
    LocalMux I__11027 (
            .O(N__46856),
            .I(N__46807));
    LocalMux I__11026 (
            .O(N__46853),
            .I(N__46807));
    Span4Mux_h I__11025 (
            .O(N__46850),
            .I(N__46804));
    Span4Mux_h I__11024 (
            .O(N__46841),
            .I(N__46801));
    LocalMux I__11023 (
            .O(N__46826),
            .I(current_pin_7__N_155));
    LocalMux I__11022 (
            .O(N__46821),
            .I(current_pin_7__N_155));
    Odrv12 I__11021 (
            .O(N__46818),
            .I(current_pin_7__N_155));
    Odrv12 I__11020 (
            .O(N__46807),
            .I(current_pin_7__N_155));
    Odrv4 I__11019 (
            .O(N__46804),
            .I(current_pin_7__N_155));
    Odrv4 I__11018 (
            .O(N__46801),
            .I(current_pin_7__N_155));
    InMux I__11017 (
            .O(N__46788),
            .I(N__46783));
    InMux I__11016 (
            .O(N__46787),
            .I(N__46778));
    InMux I__11015 (
            .O(N__46786),
            .I(N__46778));
    LocalMux I__11014 (
            .O(N__46783),
            .I(N__46769));
    LocalMux I__11013 (
            .O(N__46778),
            .I(N__46769));
    InMux I__11012 (
            .O(N__46777),
            .I(N__46766));
    InMux I__11011 (
            .O(N__46776),
            .I(N__46763));
    InMux I__11010 (
            .O(N__46775),
            .I(N__46758));
    InMux I__11009 (
            .O(N__46774),
            .I(N__46758));
    Span4Mux_h I__11008 (
            .O(N__46769),
            .I(N__46755));
    LocalMux I__11007 (
            .O(N__46766),
            .I(n7_adj_719));
    LocalMux I__11006 (
            .O(N__46763),
            .I(n7_adj_719));
    LocalMux I__11005 (
            .O(N__46758),
            .I(n7_adj_719));
    Odrv4 I__11004 (
            .O(N__46755),
            .I(n7_adj_719));
    CascadeMux I__11003 (
            .O(N__46746),
            .I(N__46740));
    CascadeMux I__11002 (
            .O(N__46745),
            .I(N__46737));
    InMux I__11001 (
            .O(N__46744),
            .I(N__46734));
    InMux I__11000 (
            .O(N__46743),
            .I(N__46729));
    InMux I__10999 (
            .O(N__46740),
            .I(N__46729));
    InMux I__10998 (
            .O(N__46737),
            .I(N__46726));
    LocalMux I__10997 (
            .O(N__46734),
            .I(N__46723));
    LocalMux I__10996 (
            .O(N__46729),
            .I(N__46719));
    LocalMux I__10995 (
            .O(N__46726),
            .I(N__46716));
    Span4Mux_h I__10994 (
            .O(N__46723),
            .I(N__46713));
    InMux I__10993 (
            .O(N__46722),
            .I(N__46710));
    Span4Mux_h I__10992 (
            .O(N__46719),
            .I(N__46705));
    Span4Mux_v I__10991 (
            .O(N__46716),
            .I(N__46705));
    Span4Mux_h I__10990 (
            .O(N__46713),
            .I(N__46702));
    LocalMux I__10989 (
            .O(N__46710),
            .I(n21));
    Odrv4 I__10988 (
            .O(N__46705),
            .I(n21));
    Odrv4 I__10987 (
            .O(N__46702),
            .I(n21));
    CascadeMux I__10986 (
            .O(N__46695),
            .I(current_pin_7__N_155_cascade_));
    CascadeMux I__10985 (
            .O(N__46692),
            .I(N__46689));
    InMux I__10984 (
            .O(N__46689),
            .I(N__46684));
    CascadeMux I__10983 (
            .O(N__46688),
            .I(N__46680));
    InMux I__10982 (
            .O(N__46687),
            .I(N__46674));
    LocalMux I__10981 (
            .O(N__46684),
            .I(N__46671));
    InMux I__10980 (
            .O(N__46683),
            .I(N__46666));
    InMux I__10979 (
            .O(N__46680),
            .I(N__46663));
    InMux I__10978 (
            .O(N__46679),
            .I(N__46658));
    InMux I__10977 (
            .O(N__46678),
            .I(N__46658));
    InMux I__10976 (
            .O(N__46677),
            .I(N__46654));
    LocalMux I__10975 (
            .O(N__46674),
            .I(N__46651));
    Span4Mux_v I__10974 (
            .O(N__46671),
            .I(N__46648));
    InMux I__10973 (
            .O(N__46670),
            .I(N__46643));
    InMux I__10972 (
            .O(N__46669),
            .I(N__46643));
    LocalMux I__10971 (
            .O(N__46666),
            .I(N__46639));
    LocalMux I__10970 (
            .O(N__46663),
            .I(N__46634));
    LocalMux I__10969 (
            .O(N__46658),
            .I(N__46634));
    InMux I__10968 (
            .O(N__46657),
            .I(N__46631));
    LocalMux I__10967 (
            .O(N__46654),
            .I(N__46626));
    Span4Mux_v I__10966 (
            .O(N__46651),
            .I(N__46626));
    Span4Mux_h I__10965 (
            .O(N__46648),
            .I(N__46621));
    LocalMux I__10964 (
            .O(N__46643),
            .I(N__46621));
    InMux I__10963 (
            .O(N__46642),
            .I(N__46618));
    Span4Mux_h I__10962 (
            .O(N__46639),
            .I(N__46613));
    Span4Mux_h I__10961 (
            .O(N__46634),
            .I(N__46613));
    LocalMux I__10960 (
            .O(N__46631),
            .I(n7166));
    Odrv4 I__10959 (
            .O(N__46626),
            .I(n7166));
    Odrv4 I__10958 (
            .O(N__46621),
            .I(n7166));
    LocalMux I__10957 (
            .O(N__46618),
            .I(n7166));
    Odrv4 I__10956 (
            .O(N__46613),
            .I(n7166));
    CascadeMux I__10955 (
            .O(N__46602),
            .I(N__46599));
    InMux I__10954 (
            .O(N__46599),
            .I(N__46596));
    LocalMux I__10953 (
            .O(N__46596),
            .I(N__46593));
    Span4Mux_h I__10952 (
            .O(N__46593),
            .I(N__46589));
    InMux I__10951 (
            .O(N__46592),
            .I(N__46586));
    Odrv4 I__10950 (
            .O(N__46589),
            .I(n6180));
    LocalMux I__10949 (
            .O(N__46586),
            .I(n6180));
    InMux I__10948 (
            .O(N__46581),
            .I(N__46571));
    InMux I__10947 (
            .O(N__46580),
            .I(N__46571));
    InMux I__10946 (
            .O(N__46579),
            .I(N__46571));
    InMux I__10945 (
            .O(N__46578),
            .I(N__46564));
    LocalMux I__10944 (
            .O(N__46571),
            .I(N__46561));
    InMux I__10943 (
            .O(N__46570),
            .I(N__46552));
    InMux I__10942 (
            .O(N__46569),
            .I(N__46552));
    InMux I__10941 (
            .O(N__46568),
            .I(N__46552));
    InMux I__10940 (
            .O(N__46567),
            .I(N__46552));
    LocalMux I__10939 (
            .O(N__46564),
            .I(N__46549));
    Odrv4 I__10938 (
            .O(N__46561),
            .I(n6971));
    LocalMux I__10937 (
            .O(N__46552),
            .I(n6971));
    Odrv4 I__10936 (
            .O(N__46549),
            .I(n6971));
    InMux I__10935 (
            .O(N__46542),
            .I(N__46539));
    LocalMux I__10934 (
            .O(N__46539),
            .I(n12135));
    InMux I__10933 (
            .O(N__46536),
            .I(N__46531));
    InMux I__10932 (
            .O(N__46535),
            .I(N__46525));
    InMux I__10931 (
            .O(N__46534),
            .I(N__46520));
    LocalMux I__10930 (
            .O(N__46531),
            .I(N__46512));
    InMux I__10929 (
            .O(N__46530),
            .I(N__46509));
    InMux I__10928 (
            .O(N__46529),
            .I(N__46506));
    InMux I__10927 (
            .O(N__46528),
            .I(N__46503));
    LocalMux I__10926 (
            .O(N__46525),
            .I(N__46500));
    InMux I__10925 (
            .O(N__46524),
            .I(N__46495));
    InMux I__10924 (
            .O(N__46523),
            .I(N__46495));
    LocalMux I__10923 (
            .O(N__46520),
            .I(N__46492));
    InMux I__10922 (
            .O(N__46519),
            .I(N__46489));
    InMux I__10921 (
            .O(N__46518),
            .I(N__46484));
    InMux I__10920 (
            .O(N__46517),
            .I(N__46476));
    InMux I__10919 (
            .O(N__46516),
            .I(N__46476));
    InMux I__10918 (
            .O(N__46515),
            .I(N__46472));
    Span4Mux_v I__10917 (
            .O(N__46512),
            .I(N__46467));
    LocalMux I__10916 (
            .O(N__46509),
            .I(N__46467));
    LocalMux I__10915 (
            .O(N__46506),
            .I(N__46464));
    LocalMux I__10914 (
            .O(N__46503),
            .I(N__46457));
    Span4Mux_h I__10913 (
            .O(N__46500),
            .I(N__46457));
    LocalMux I__10912 (
            .O(N__46495),
            .I(N__46457));
    Span4Mux_h I__10911 (
            .O(N__46492),
            .I(N__46452));
    LocalMux I__10910 (
            .O(N__46489),
            .I(N__46452));
    InMux I__10909 (
            .O(N__46488),
            .I(N__46445));
    InMux I__10908 (
            .O(N__46487),
            .I(N__46442));
    LocalMux I__10907 (
            .O(N__46484),
            .I(N__46439));
    InMux I__10906 (
            .O(N__46483),
            .I(N__46436));
    InMux I__10905 (
            .O(N__46482),
            .I(N__46431));
    InMux I__10904 (
            .O(N__46481),
            .I(N__46431));
    LocalMux I__10903 (
            .O(N__46476),
            .I(N__46428));
    InMux I__10902 (
            .O(N__46475),
            .I(N__46425));
    LocalMux I__10901 (
            .O(N__46472),
            .I(N__46422));
    Span4Mux_h I__10900 (
            .O(N__46467),
            .I(N__46417));
    Span4Mux_v I__10899 (
            .O(N__46464),
            .I(N__46417));
    Span4Mux_v I__10898 (
            .O(N__46457),
            .I(N__46414));
    Span4Mux_v I__10897 (
            .O(N__46452),
            .I(N__46411));
    InMux I__10896 (
            .O(N__46451),
            .I(N__46408));
    InMux I__10895 (
            .O(N__46450),
            .I(N__46401));
    InMux I__10894 (
            .O(N__46449),
            .I(N__46401));
    InMux I__10893 (
            .O(N__46448),
            .I(N__46401));
    LocalMux I__10892 (
            .O(N__46445),
            .I(N__46396));
    LocalMux I__10891 (
            .O(N__46442),
            .I(N__46396));
    Span4Mux_v I__10890 (
            .O(N__46439),
            .I(N__46393));
    LocalMux I__10889 (
            .O(N__46436),
            .I(N__46384));
    LocalMux I__10888 (
            .O(N__46431),
            .I(N__46384));
    Span4Mux_h I__10887 (
            .O(N__46428),
            .I(N__46384));
    LocalMux I__10886 (
            .O(N__46425),
            .I(N__46384));
    Span12Mux_v I__10885 (
            .O(N__46422),
            .I(N__46381));
    Span4Mux_h I__10884 (
            .O(N__46417),
            .I(N__46376));
    Span4Mux_h I__10883 (
            .O(N__46414),
            .I(N__46376));
    Span4Mux_h I__10882 (
            .O(N__46411),
            .I(N__46371));
    LocalMux I__10881 (
            .O(N__46408),
            .I(N__46371));
    LocalMux I__10880 (
            .O(N__46401),
            .I(n149));
    Odrv12 I__10879 (
            .O(N__46396),
            .I(n149));
    Odrv4 I__10878 (
            .O(N__46393),
            .I(n149));
    Odrv4 I__10877 (
            .O(N__46384),
            .I(n149));
    Odrv12 I__10876 (
            .O(N__46381),
            .I(n149));
    Odrv4 I__10875 (
            .O(N__46376),
            .I(n149));
    Odrv4 I__10874 (
            .O(N__46371),
            .I(n149));
    InMux I__10873 (
            .O(N__46356),
            .I(n10572));
    InMux I__10872 (
            .O(N__46353),
            .I(N__46349));
    InMux I__10871 (
            .O(N__46352),
            .I(N__46346));
    LocalMux I__10870 (
            .O(N__46349),
            .I(blink_counter_25));
    LocalMux I__10869 (
            .O(N__46346),
            .I(blink_counter_25));
    InMux I__10868 (
            .O(N__46341),
            .I(N__46338));
    LocalMux I__10867 (
            .O(N__46338),
            .I(n45));
    InMux I__10866 (
            .O(N__46335),
            .I(bfn_16_15_0_));
    InMux I__10865 (
            .O(N__46332),
            .I(n10510));
    InMux I__10864 (
            .O(N__46329),
            .I(n10511));
    InMux I__10863 (
            .O(N__46326),
            .I(n10512));
    InMux I__10862 (
            .O(N__46323),
            .I(n10513));
    InMux I__10861 (
            .O(N__46320),
            .I(n10514));
    InMux I__10860 (
            .O(N__46317),
            .I(n10515));
    InMux I__10859 (
            .O(N__46314),
            .I(N__46311));
    LocalMux I__10858 (
            .O(N__46311),
            .I(n9));
    InMux I__10857 (
            .O(N__46308),
            .I(n10564));
    InMux I__10856 (
            .O(N__46305),
            .I(N__46302));
    LocalMux I__10855 (
            .O(N__46302),
            .I(n8_adj_755));
    InMux I__10854 (
            .O(N__46299),
            .I(n10565));
    InMux I__10853 (
            .O(N__46296),
            .I(N__46293));
    LocalMux I__10852 (
            .O(N__46293),
            .I(n7));
    InMux I__10851 (
            .O(N__46290),
            .I(n10566));
    InMux I__10850 (
            .O(N__46287),
            .I(N__46284));
    LocalMux I__10849 (
            .O(N__46284),
            .I(n6_adj_756));
    InMux I__10848 (
            .O(N__46281),
            .I(n10567));
    CascadeMux I__10847 (
            .O(N__46278),
            .I(N__46275));
    InMux I__10846 (
            .O(N__46275),
            .I(N__46268));
    InMux I__10845 (
            .O(N__46274),
            .I(N__46268));
    InMux I__10844 (
            .O(N__46273),
            .I(N__46265));
    LocalMux I__10843 (
            .O(N__46268),
            .I(blink_counter_21));
    LocalMux I__10842 (
            .O(N__46265),
            .I(blink_counter_21));
    InMux I__10841 (
            .O(N__46260),
            .I(n10568));
    InMux I__10840 (
            .O(N__46257),
            .I(N__46250));
    InMux I__10839 (
            .O(N__46256),
            .I(N__46250));
    InMux I__10838 (
            .O(N__46255),
            .I(N__46247));
    LocalMux I__10837 (
            .O(N__46250),
            .I(blink_counter_22));
    LocalMux I__10836 (
            .O(N__46247),
            .I(blink_counter_22));
    InMux I__10835 (
            .O(N__46242),
            .I(n10569));
    CascadeMux I__10834 (
            .O(N__46239),
            .I(N__46235));
    InMux I__10833 (
            .O(N__46238),
            .I(N__46229));
    InMux I__10832 (
            .O(N__46235),
            .I(N__46229));
    InMux I__10831 (
            .O(N__46234),
            .I(N__46226));
    LocalMux I__10830 (
            .O(N__46229),
            .I(blink_counter_23));
    LocalMux I__10829 (
            .O(N__46226),
            .I(blink_counter_23));
    InMux I__10828 (
            .O(N__46221),
            .I(n10570));
    InMux I__10827 (
            .O(N__46218),
            .I(N__46211));
    InMux I__10826 (
            .O(N__46217),
            .I(N__46211));
    InMux I__10825 (
            .O(N__46216),
            .I(N__46208));
    LocalMux I__10824 (
            .O(N__46211),
            .I(blink_counter_24));
    LocalMux I__10823 (
            .O(N__46208),
            .I(blink_counter_24));
    InMux I__10822 (
            .O(N__46203),
            .I(bfn_15_29_0_));
    InMux I__10821 (
            .O(N__46200),
            .I(N__46197));
    LocalMux I__10820 (
            .O(N__46197),
            .I(n18));
    InMux I__10819 (
            .O(N__46194),
            .I(bfn_15_27_0_));
    InMux I__10818 (
            .O(N__46191),
            .I(N__46188));
    LocalMux I__10817 (
            .O(N__46188),
            .I(n17));
    InMux I__10816 (
            .O(N__46185),
            .I(n10556));
    InMux I__10815 (
            .O(N__46182),
            .I(N__46179));
    LocalMux I__10814 (
            .O(N__46179),
            .I(n16));
    InMux I__10813 (
            .O(N__46176),
            .I(n10557));
    InMux I__10812 (
            .O(N__46173),
            .I(N__46170));
    LocalMux I__10811 (
            .O(N__46170),
            .I(n15_adj_759));
    InMux I__10810 (
            .O(N__46167),
            .I(n10558));
    InMux I__10809 (
            .O(N__46164),
            .I(N__46161));
    LocalMux I__10808 (
            .O(N__46161),
            .I(n14_adj_745));
    InMux I__10807 (
            .O(N__46158),
            .I(n10559));
    InMux I__10806 (
            .O(N__46155),
            .I(N__46152));
    LocalMux I__10805 (
            .O(N__46152),
            .I(n13));
    InMux I__10804 (
            .O(N__46149),
            .I(n10560));
    InMux I__10803 (
            .O(N__46146),
            .I(N__46143));
    LocalMux I__10802 (
            .O(N__46143),
            .I(n12));
    InMux I__10801 (
            .O(N__46140),
            .I(n10561));
    InMux I__10800 (
            .O(N__46137),
            .I(N__46134));
    LocalMux I__10799 (
            .O(N__46134),
            .I(n11_adj_758));
    InMux I__10798 (
            .O(N__46131),
            .I(n10562));
    InMux I__10797 (
            .O(N__46128),
            .I(N__46125));
    LocalMux I__10796 (
            .O(N__46125),
            .I(n10_adj_757));
    InMux I__10795 (
            .O(N__46122),
            .I(bfn_15_28_0_));
    InMux I__10794 (
            .O(N__46119),
            .I(N__46116));
    LocalMux I__10793 (
            .O(N__46116),
            .I(n26));
    InMux I__10792 (
            .O(N__46113),
            .I(bfn_15_26_0_));
    InMux I__10791 (
            .O(N__46110),
            .I(N__46107));
    LocalMux I__10790 (
            .O(N__46107),
            .I(n25));
    InMux I__10789 (
            .O(N__46104),
            .I(n10548));
    InMux I__10788 (
            .O(N__46101),
            .I(N__46098));
    LocalMux I__10787 (
            .O(N__46098),
            .I(n24));
    InMux I__10786 (
            .O(N__46095),
            .I(n10549));
    InMux I__10785 (
            .O(N__46092),
            .I(N__46089));
    LocalMux I__10784 (
            .O(N__46089),
            .I(n23));
    InMux I__10783 (
            .O(N__46086),
            .I(n10550));
    InMux I__10782 (
            .O(N__46083),
            .I(N__46080));
    LocalMux I__10781 (
            .O(N__46080),
            .I(n22));
    InMux I__10780 (
            .O(N__46077),
            .I(n10551));
    InMux I__10779 (
            .O(N__46074),
            .I(N__46071));
    LocalMux I__10778 (
            .O(N__46071),
            .I(n21_adj_737));
    InMux I__10777 (
            .O(N__46068),
            .I(n10552));
    InMux I__10776 (
            .O(N__46065),
            .I(N__46062));
    LocalMux I__10775 (
            .O(N__46062),
            .I(n20));
    InMux I__10774 (
            .O(N__46059),
            .I(n10553));
    InMux I__10773 (
            .O(N__46056),
            .I(N__46053));
    LocalMux I__10772 (
            .O(N__46053),
            .I(n19_adj_718));
    InMux I__10771 (
            .O(N__46050),
            .I(n10554));
    InMux I__10770 (
            .O(N__46047),
            .I(N__46043));
    CascadeMux I__10769 (
            .O(N__46046),
            .I(N__46040));
    LocalMux I__10768 (
            .O(N__46043),
            .I(N__46036));
    InMux I__10767 (
            .O(N__46040),
            .I(N__46033));
    InMux I__10766 (
            .O(N__46039),
            .I(N__46030));
    Odrv4 I__10765 (
            .O(N__46036),
            .I(\nx.n2298 ));
    LocalMux I__10764 (
            .O(N__46033),
            .I(\nx.n2298 ));
    LocalMux I__10763 (
            .O(N__46030),
            .I(\nx.n2298 ));
    CascadeMux I__10762 (
            .O(N__46023),
            .I(N__46020));
    InMux I__10761 (
            .O(N__46020),
            .I(N__46017));
    LocalMux I__10760 (
            .O(N__46017),
            .I(N__46014));
    Odrv4 I__10759 (
            .O(N__46014),
            .I(\nx.n2365 ));
    InMux I__10758 (
            .O(N__46011),
            .I(\nx.n10719 ));
    CascadeMux I__10757 (
            .O(N__46008),
            .I(N__46004));
    CascadeMux I__10756 (
            .O(N__46007),
            .I(N__46001));
    InMux I__10755 (
            .O(N__46004),
            .I(N__45998));
    InMux I__10754 (
            .O(N__46001),
            .I(N__45995));
    LocalMux I__10753 (
            .O(N__45998),
            .I(\nx.n2297 ));
    LocalMux I__10752 (
            .O(N__45995),
            .I(\nx.n2297 ));
    InMux I__10751 (
            .O(N__45990),
            .I(N__45987));
    LocalMux I__10750 (
            .O(N__45987),
            .I(\nx.n2364 ));
    InMux I__10749 (
            .O(N__45984),
            .I(\nx.n10720 ));
    CascadeMux I__10748 (
            .O(N__45981),
            .I(N__45978));
    InMux I__10747 (
            .O(N__45978),
            .I(N__45975));
    LocalMux I__10746 (
            .O(N__45975),
            .I(N__45972));
    Span4Mux_v I__10745 (
            .O(N__45972),
            .I(N__45968));
    InMux I__10744 (
            .O(N__45971),
            .I(N__45965));
    Odrv4 I__10743 (
            .O(N__45968),
            .I(\nx.n2296 ));
    LocalMux I__10742 (
            .O(N__45965),
            .I(\nx.n2296 ));
    InMux I__10741 (
            .O(N__45960),
            .I(N__45957));
    LocalMux I__10740 (
            .O(N__45957),
            .I(N__45954));
    Span4Mux_h I__10739 (
            .O(N__45954),
            .I(N__45951));
    Odrv4 I__10738 (
            .O(N__45951),
            .I(\nx.n2363 ));
    InMux I__10737 (
            .O(N__45948),
            .I(\nx.n10721 ));
    CascadeMux I__10736 (
            .O(N__45945),
            .I(N__45942));
    InMux I__10735 (
            .O(N__45942),
            .I(N__45939));
    LocalMux I__10734 (
            .O(N__45939),
            .I(N__45935));
    InMux I__10733 (
            .O(N__45938),
            .I(N__45931));
    Span4Mux_h I__10732 (
            .O(N__45935),
            .I(N__45928));
    InMux I__10731 (
            .O(N__45934),
            .I(N__45925));
    LocalMux I__10730 (
            .O(N__45931),
            .I(\nx.n2295 ));
    Odrv4 I__10729 (
            .O(N__45928),
            .I(\nx.n2295 ));
    LocalMux I__10728 (
            .O(N__45925),
            .I(\nx.n2295 ));
    CascadeMux I__10727 (
            .O(N__45918),
            .I(N__45915));
    InMux I__10726 (
            .O(N__45915),
            .I(N__45912));
    LocalMux I__10725 (
            .O(N__45912),
            .I(N__45909));
    Span4Mux_h I__10724 (
            .O(N__45909),
            .I(N__45906));
    Span4Mux_h I__10723 (
            .O(N__45906),
            .I(N__45903));
    Odrv4 I__10722 (
            .O(N__45903),
            .I(\nx.n2362 ));
    InMux I__10721 (
            .O(N__45900),
            .I(\nx.n10722 ));
    CascadeMux I__10720 (
            .O(N__45897),
            .I(N__45894));
    InMux I__10719 (
            .O(N__45894),
            .I(N__45891));
    LocalMux I__10718 (
            .O(N__45891),
            .I(N__45887));
    InMux I__10717 (
            .O(N__45890),
            .I(N__45883));
    Span4Mux_h I__10716 (
            .O(N__45887),
            .I(N__45880));
    InMux I__10715 (
            .O(N__45886),
            .I(N__45877));
    LocalMux I__10714 (
            .O(N__45883),
            .I(\nx.n2294 ));
    Odrv4 I__10713 (
            .O(N__45880),
            .I(\nx.n2294 ));
    LocalMux I__10712 (
            .O(N__45877),
            .I(\nx.n2294 ));
    InMux I__10711 (
            .O(N__45870),
            .I(N__45867));
    LocalMux I__10710 (
            .O(N__45867),
            .I(N__45864));
    Span4Mux_h I__10709 (
            .O(N__45864),
            .I(N__45861));
    Span4Mux_h I__10708 (
            .O(N__45861),
            .I(N__45858));
    Odrv4 I__10707 (
            .O(N__45858),
            .I(\nx.n2361 ));
    InMux I__10706 (
            .O(N__45855),
            .I(bfn_15_25_0_));
    CascadeMux I__10705 (
            .O(N__45852),
            .I(N__45849));
    InMux I__10704 (
            .O(N__45849),
            .I(N__45845));
    CascadeMux I__10703 (
            .O(N__45848),
            .I(N__45842));
    LocalMux I__10702 (
            .O(N__45845),
            .I(N__45839));
    InMux I__10701 (
            .O(N__45842),
            .I(N__45836));
    Span4Mux_h I__10700 (
            .O(N__45839),
            .I(N__45833));
    LocalMux I__10699 (
            .O(N__45836),
            .I(\nx.n2293 ));
    Odrv4 I__10698 (
            .O(N__45833),
            .I(\nx.n2293 ));
    InMux I__10697 (
            .O(N__45828),
            .I(N__45825));
    LocalMux I__10696 (
            .O(N__45825),
            .I(N__45822));
    Span4Mux_h I__10695 (
            .O(N__45822),
            .I(N__45819));
    Span4Mux_h I__10694 (
            .O(N__45819),
            .I(N__45816));
    Odrv4 I__10693 (
            .O(N__45816),
            .I(\nx.n2360 ));
    InMux I__10692 (
            .O(N__45813),
            .I(\nx.n10724 ));
    CascadeMux I__10691 (
            .O(N__45810),
            .I(N__45807));
    InMux I__10690 (
            .O(N__45807),
            .I(N__45802));
    CascadeMux I__10689 (
            .O(N__45806),
            .I(N__45799));
    CascadeMux I__10688 (
            .O(N__45805),
            .I(N__45796));
    LocalMux I__10687 (
            .O(N__45802),
            .I(N__45793));
    InMux I__10686 (
            .O(N__45799),
            .I(N__45790));
    InMux I__10685 (
            .O(N__45796),
            .I(N__45787));
    Span4Mux_h I__10684 (
            .O(N__45793),
            .I(N__45784));
    LocalMux I__10683 (
            .O(N__45790),
            .I(\nx.n2292 ));
    LocalMux I__10682 (
            .O(N__45787),
            .I(\nx.n2292 ));
    Odrv4 I__10681 (
            .O(N__45784),
            .I(\nx.n2292 ));
    InMux I__10680 (
            .O(N__45777),
            .I(N__45774));
    LocalMux I__10679 (
            .O(N__45774),
            .I(N__45771));
    Odrv4 I__10678 (
            .O(N__45771),
            .I(\nx.n2359 ));
    InMux I__10677 (
            .O(N__45768),
            .I(\nx.n10725 ));
    CascadeMux I__10676 (
            .O(N__45765),
            .I(N__45734));
    CascadeMux I__10675 (
            .O(N__45764),
            .I(N__45724));
    CascadeMux I__10674 (
            .O(N__45763),
            .I(N__45721));
    CascadeMux I__10673 (
            .O(N__45762),
            .I(N__45717));
    CascadeMux I__10672 (
            .O(N__45761),
            .I(N__45714));
    CascadeMux I__10671 (
            .O(N__45760),
            .I(N__45711));
    CascadeMux I__10670 (
            .O(N__45759),
            .I(N__45708));
    CascadeMux I__10669 (
            .O(N__45758),
            .I(N__45705));
    InMux I__10668 (
            .O(N__45757),
            .I(N__45701));
    CascadeMux I__10667 (
            .O(N__45756),
            .I(N__45681));
    CascadeMux I__10666 (
            .O(N__45755),
            .I(N__45673));
    CascadeMux I__10665 (
            .O(N__45754),
            .I(N__45667));
    CascadeMux I__10664 (
            .O(N__45753),
            .I(N__45662));
    CascadeMux I__10663 (
            .O(N__45752),
            .I(N__45651));
    CascadeMux I__10662 (
            .O(N__45751),
            .I(N__45639));
    CascadeMux I__10661 (
            .O(N__45750),
            .I(N__45636));
    InMux I__10660 (
            .O(N__45749),
            .I(N__45616));
    InMux I__10659 (
            .O(N__45748),
            .I(N__45616));
    InMux I__10658 (
            .O(N__45747),
            .I(N__45616));
    InMux I__10657 (
            .O(N__45746),
            .I(N__45616));
    InMux I__10656 (
            .O(N__45745),
            .I(N__45607));
    InMux I__10655 (
            .O(N__45744),
            .I(N__45607));
    InMux I__10654 (
            .O(N__45743),
            .I(N__45607));
    InMux I__10653 (
            .O(N__45742),
            .I(N__45607));
    InMux I__10652 (
            .O(N__45741),
            .I(N__45600));
    InMux I__10651 (
            .O(N__45740),
            .I(N__45600));
    InMux I__10650 (
            .O(N__45739),
            .I(N__45600));
    InMux I__10649 (
            .O(N__45738),
            .I(N__45591));
    InMux I__10648 (
            .O(N__45737),
            .I(N__45591));
    InMux I__10647 (
            .O(N__45734),
            .I(N__45591));
    InMux I__10646 (
            .O(N__45733),
            .I(N__45591));
    CascadeMux I__10645 (
            .O(N__45732),
            .I(N__45581));
    CascadeMux I__10644 (
            .O(N__45731),
            .I(N__45573));
    CascadeMux I__10643 (
            .O(N__45730),
            .I(N__45559));
    CascadeMux I__10642 (
            .O(N__45729),
            .I(N__45544));
    CascadeMux I__10641 (
            .O(N__45728),
            .I(N__45536));
    CascadeMux I__10640 (
            .O(N__45727),
            .I(N__45527));
    InMux I__10639 (
            .O(N__45724),
            .I(N__45514));
    InMux I__10638 (
            .O(N__45721),
            .I(N__45514));
    InMux I__10637 (
            .O(N__45720),
            .I(N__45514));
    InMux I__10636 (
            .O(N__45717),
            .I(N__45514));
    InMux I__10635 (
            .O(N__45714),
            .I(N__45514));
    InMux I__10634 (
            .O(N__45711),
            .I(N__45507));
    InMux I__10633 (
            .O(N__45708),
            .I(N__45507));
    InMux I__10632 (
            .O(N__45705),
            .I(N__45507));
    CascadeMux I__10631 (
            .O(N__45704),
            .I(N__45498));
    LocalMux I__10630 (
            .O(N__45701),
            .I(N__45493));
    InMux I__10629 (
            .O(N__45700),
            .I(N__45486));
    InMux I__10628 (
            .O(N__45699),
            .I(N__45486));
    InMux I__10627 (
            .O(N__45698),
            .I(N__45486));
    InMux I__10626 (
            .O(N__45697),
            .I(N__45479));
    InMux I__10625 (
            .O(N__45696),
            .I(N__45479));
    InMux I__10624 (
            .O(N__45695),
            .I(N__45479));
    InMux I__10623 (
            .O(N__45694),
            .I(N__45470));
    InMux I__10622 (
            .O(N__45693),
            .I(N__45470));
    InMux I__10621 (
            .O(N__45692),
            .I(N__45470));
    InMux I__10620 (
            .O(N__45691),
            .I(N__45470));
    InMux I__10619 (
            .O(N__45690),
            .I(N__45463));
    InMux I__10618 (
            .O(N__45689),
            .I(N__45463));
    InMux I__10617 (
            .O(N__45688),
            .I(N__45463));
    InMux I__10616 (
            .O(N__45687),
            .I(N__45456));
    InMux I__10615 (
            .O(N__45686),
            .I(N__45456));
    InMux I__10614 (
            .O(N__45685),
            .I(N__45456));
    InMux I__10613 (
            .O(N__45684),
            .I(N__45423));
    InMux I__10612 (
            .O(N__45681),
            .I(N__45423));
    InMux I__10611 (
            .O(N__45680),
            .I(N__45423));
    InMux I__10610 (
            .O(N__45679),
            .I(N__45423));
    InMux I__10609 (
            .O(N__45678),
            .I(N__45418));
    InMux I__10608 (
            .O(N__45677),
            .I(N__45418));
    InMux I__10607 (
            .O(N__45676),
            .I(N__45402));
    InMux I__10606 (
            .O(N__45673),
            .I(N__45402));
    InMux I__10605 (
            .O(N__45672),
            .I(N__45402));
    InMux I__10604 (
            .O(N__45671),
            .I(N__45402));
    CascadeMux I__10603 (
            .O(N__45670),
            .I(N__45396));
    InMux I__10602 (
            .O(N__45667),
            .I(N__45386));
    InMux I__10601 (
            .O(N__45666),
            .I(N__45386));
    InMux I__10600 (
            .O(N__45665),
            .I(N__45375));
    InMux I__10599 (
            .O(N__45662),
            .I(N__45375));
    InMux I__10598 (
            .O(N__45661),
            .I(N__45375));
    InMux I__10597 (
            .O(N__45660),
            .I(N__45375));
    InMux I__10596 (
            .O(N__45659),
            .I(N__45375));
    InMux I__10595 (
            .O(N__45658),
            .I(N__45368));
    InMux I__10594 (
            .O(N__45657),
            .I(N__45368));
    InMux I__10593 (
            .O(N__45656),
            .I(N__45368));
    InMux I__10592 (
            .O(N__45655),
            .I(N__45357));
    InMux I__10591 (
            .O(N__45654),
            .I(N__45357));
    InMux I__10590 (
            .O(N__45651),
            .I(N__45357));
    InMux I__10589 (
            .O(N__45650),
            .I(N__45357));
    InMux I__10588 (
            .O(N__45649),
            .I(N__45357));
    InMux I__10587 (
            .O(N__45648),
            .I(N__45348));
    InMux I__10586 (
            .O(N__45647),
            .I(N__45348));
    InMux I__10585 (
            .O(N__45646),
            .I(N__45348));
    InMux I__10584 (
            .O(N__45645),
            .I(N__45348));
    InMux I__10583 (
            .O(N__45644),
            .I(N__45339));
    InMux I__10582 (
            .O(N__45643),
            .I(N__45339));
    InMux I__10581 (
            .O(N__45642),
            .I(N__45339));
    InMux I__10580 (
            .O(N__45639),
            .I(N__45339));
    InMux I__10579 (
            .O(N__45636),
            .I(N__45333));
    InMux I__10578 (
            .O(N__45635),
            .I(N__45333));
    InMux I__10577 (
            .O(N__45634),
            .I(N__45326));
    InMux I__10576 (
            .O(N__45633),
            .I(N__45326));
    InMux I__10575 (
            .O(N__45632),
            .I(N__45326));
    CascadeMux I__10574 (
            .O(N__45631),
            .I(N__45319));
    CascadeMux I__10573 (
            .O(N__45630),
            .I(N__45314));
    CascadeMux I__10572 (
            .O(N__45629),
            .I(N__45304));
    CascadeMux I__10571 (
            .O(N__45628),
            .I(N__45299));
    CascadeMux I__10570 (
            .O(N__45627),
            .I(N__45293));
    CascadeMux I__10569 (
            .O(N__45626),
            .I(N__45289));
    CascadeMux I__10568 (
            .O(N__45625),
            .I(N__45286));
    LocalMux I__10567 (
            .O(N__45616),
            .I(N__45276));
    LocalMux I__10566 (
            .O(N__45607),
            .I(N__45269));
    LocalMux I__10565 (
            .O(N__45600),
            .I(N__45269));
    LocalMux I__10564 (
            .O(N__45591),
            .I(N__45269));
    InMux I__10563 (
            .O(N__45590),
            .I(N__45262));
    InMux I__10562 (
            .O(N__45589),
            .I(N__45262));
    InMux I__10561 (
            .O(N__45588),
            .I(N__45262));
    InMux I__10560 (
            .O(N__45587),
            .I(N__45251));
    InMux I__10559 (
            .O(N__45586),
            .I(N__45251));
    InMux I__10558 (
            .O(N__45585),
            .I(N__45251));
    InMux I__10557 (
            .O(N__45584),
            .I(N__45251));
    InMux I__10556 (
            .O(N__45581),
            .I(N__45251));
    InMux I__10555 (
            .O(N__45580),
            .I(N__45244));
    InMux I__10554 (
            .O(N__45579),
            .I(N__45244));
    InMux I__10553 (
            .O(N__45578),
            .I(N__45244));
    InMux I__10552 (
            .O(N__45577),
            .I(N__45239));
    InMux I__10551 (
            .O(N__45576),
            .I(N__45239));
    InMux I__10550 (
            .O(N__45573),
            .I(N__45232));
    InMux I__10549 (
            .O(N__45572),
            .I(N__45232));
    InMux I__10548 (
            .O(N__45571),
            .I(N__45232));
    CascadeMux I__10547 (
            .O(N__45570),
            .I(N__45228));
    CascadeMux I__10546 (
            .O(N__45569),
            .I(N__45224));
    CascadeMux I__10545 (
            .O(N__45568),
            .I(N__45220));
    InMux I__10544 (
            .O(N__45567),
            .I(N__45211));
    InMux I__10543 (
            .O(N__45566),
            .I(N__45211));
    InMux I__10542 (
            .O(N__45565),
            .I(N__45211));
    InMux I__10541 (
            .O(N__45564),
            .I(N__45206));
    InMux I__10540 (
            .O(N__45563),
            .I(N__45206));
    InMux I__10539 (
            .O(N__45562),
            .I(N__45197));
    InMux I__10538 (
            .O(N__45559),
            .I(N__45197));
    InMux I__10537 (
            .O(N__45558),
            .I(N__45197));
    InMux I__10536 (
            .O(N__45557),
            .I(N__45197));
    InMux I__10535 (
            .O(N__45556),
            .I(N__45190));
    InMux I__10534 (
            .O(N__45555),
            .I(N__45190));
    InMux I__10533 (
            .O(N__45554),
            .I(N__45190));
    InMux I__10532 (
            .O(N__45553),
            .I(N__45183));
    InMux I__10531 (
            .O(N__45552),
            .I(N__45183));
    InMux I__10530 (
            .O(N__45551),
            .I(N__45183));
    InMux I__10529 (
            .O(N__45550),
            .I(N__45174));
    InMux I__10528 (
            .O(N__45549),
            .I(N__45174));
    InMux I__10527 (
            .O(N__45548),
            .I(N__45174));
    InMux I__10526 (
            .O(N__45547),
            .I(N__45174));
    InMux I__10525 (
            .O(N__45544),
            .I(N__45163));
    InMux I__10524 (
            .O(N__45543),
            .I(N__45163));
    InMux I__10523 (
            .O(N__45542),
            .I(N__45163));
    InMux I__10522 (
            .O(N__45541),
            .I(N__45163));
    InMux I__10521 (
            .O(N__45540),
            .I(N__45163));
    InMux I__10520 (
            .O(N__45539),
            .I(N__45152));
    InMux I__10519 (
            .O(N__45536),
            .I(N__45152));
    InMux I__10518 (
            .O(N__45535),
            .I(N__45152));
    InMux I__10517 (
            .O(N__45534),
            .I(N__45152));
    InMux I__10516 (
            .O(N__45533),
            .I(N__45152));
    InMux I__10515 (
            .O(N__45532),
            .I(N__45145));
    InMux I__10514 (
            .O(N__45531),
            .I(N__45145));
    InMux I__10513 (
            .O(N__45530),
            .I(N__45145));
    InMux I__10512 (
            .O(N__45527),
            .I(N__45142));
    InMux I__10511 (
            .O(N__45526),
            .I(N__45131));
    InMux I__10510 (
            .O(N__45525),
            .I(N__45128));
    LocalMux I__10509 (
            .O(N__45514),
            .I(N__45123));
    LocalMux I__10508 (
            .O(N__45507),
            .I(N__45123));
    InMux I__10507 (
            .O(N__45506),
            .I(N__45116));
    InMux I__10506 (
            .O(N__45505),
            .I(N__45116));
    InMux I__10505 (
            .O(N__45504),
            .I(N__45116));
    InMux I__10504 (
            .O(N__45503),
            .I(N__45105));
    InMux I__10503 (
            .O(N__45502),
            .I(N__45105));
    InMux I__10502 (
            .O(N__45501),
            .I(N__45105));
    InMux I__10501 (
            .O(N__45498),
            .I(N__45105));
    InMux I__10500 (
            .O(N__45497),
            .I(N__45105));
    CascadeMux I__10499 (
            .O(N__45496),
            .I(N__45101));
    Span4Mux_v I__10498 (
            .O(N__45493),
            .I(N__45087));
    LocalMux I__10497 (
            .O(N__45486),
            .I(N__45082));
    LocalMux I__10496 (
            .O(N__45479),
            .I(N__45082));
    LocalMux I__10495 (
            .O(N__45470),
            .I(N__45079));
    LocalMux I__10494 (
            .O(N__45463),
            .I(N__45074));
    LocalMux I__10493 (
            .O(N__45456),
            .I(N__45074));
    InMux I__10492 (
            .O(N__45455),
            .I(N__45067));
    InMux I__10491 (
            .O(N__45454),
            .I(N__45067));
    InMux I__10490 (
            .O(N__45453),
            .I(N__45067));
    InMux I__10489 (
            .O(N__45452),
            .I(N__45060));
    InMux I__10488 (
            .O(N__45451),
            .I(N__45060));
    InMux I__10487 (
            .O(N__45450),
            .I(N__45060));
    InMux I__10486 (
            .O(N__45449),
            .I(N__45053));
    InMux I__10485 (
            .O(N__45448),
            .I(N__45053));
    InMux I__10484 (
            .O(N__45447),
            .I(N__45053));
    InMux I__10483 (
            .O(N__45446),
            .I(N__45046));
    InMux I__10482 (
            .O(N__45445),
            .I(N__45046));
    InMux I__10481 (
            .O(N__45444),
            .I(N__45046));
    InMux I__10480 (
            .O(N__45443),
            .I(N__45037));
    InMux I__10479 (
            .O(N__45442),
            .I(N__45037));
    InMux I__10478 (
            .O(N__45441),
            .I(N__45037));
    InMux I__10477 (
            .O(N__45440),
            .I(N__45037));
    CascadeMux I__10476 (
            .O(N__45439),
            .I(N__45033));
    CascadeMux I__10475 (
            .O(N__45438),
            .I(N__45030));
    CascadeMux I__10474 (
            .O(N__45437),
            .I(N__45020));
    InMux I__10473 (
            .O(N__45436),
            .I(N__45007));
    InMux I__10472 (
            .O(N__45435),
            .I(N__45007));
    InMux I__10471 (
            .O(N__45434),
            .I(N__45007));
    InMux I__10470 (
            .O(N__45433),
            .I(N__45007));
    InMux I__10469 (
            .O(N__45432),
            .I(N__45004));
    LocalMux I__10468 (
            .O(N__45423),
            .I(N__44999));
    LocalMux I__10467 (
            .O(N__45418),
            .I(N__44999));
    InMux I__10466 (
            .O(N__45417),
            .I(N__44990));
    InMux I__10465 (
            .O(N__45416),
            .I(N__44990));
    InMux I__10464 (
            .O(N__45415),
            .I(N__44990));
    InMux I__10463 (
            .O(N__45414),
            .I(N__44990));
    InMux I__10462 (
            .O(N__45413),
            .I(N__44983));
    InMux I__10461 (
            .O(N__45412),
            .I(N__44983));
    InMux I__10460 (
            .O(N__45411),
            .I(N__44983));
    LocalMux I__10459 (
            .O(N__45402),
            .I(N__44980));
    InMux I__10458 (
            .O(N__45401),
            .I(N__44973));
    InMux I__10457 (
            .O(N__45400),
            .I(N__44973));
    InMux I__10456 (
            .O(N__45399),
            .I(N__44973));
    InMux I__10455 (
            .O(N__45396),
            .I(N__44962));
    InMux I__10454 (
            .O(N__45395),
            .I(N__44962));
    InMux I__10453 (
            .O(N__45394),
            .I(N__44962));
    InMux I__10452 (
            .O(N__45393),
            .I(N__44962));
    InMux I__10451 (
            .O(N__45392),
            .I(N__44962));
    CascadeMux I__10450 (
            .O(N__45391),
            .I(N__44959));
    LocalMux I__10449 (
            .O(N__45386),
            .I(N__44950));
    LocalMux I__10448 (
            .O(N__45375),
            .I(N__44950));
    LocalMux I__10447 (
            .O(N__45368),
            .I(N__44941));
    LocalMux I__10446 (
            .O(N__45357),
            .I(N__44941));
    LocalMux I__10445 (
            .O(N__45348),
            .I(N__44941));
    LocalMux I__10444 (
            .O(N__45339),
            .I(N__44941));
    InMux I__10443 (
            .O(N__45338),
            .I(N__44938));
    LocalMux I__10442 (
            .O(N__45333),
            .I(N__44918));
    LocalMux I__10441 (
            .O(N__45326),
            .I(N__44918));
    InMux I__10440 (
            .O(N__45325),
            .I(N__44907));
    InMux I__10439 (
            .O(N__45324),
            .I(N__44907));
    InMux I__10438 (
            .O(N__45323),
            .I(N__44907));
    InMux I__10437 (
            .O(N__45322),
            .I(N__44907));
    InMux I__10436 (
            .O(N__45319),
            .I(N__44907));
    InMux I__10435 (
            .O(N__45318),
            .I(N__44900));
    InMux I__10434 (
            .O(N__45317),
            .I(N__44900));
    InMux I__10433 (
            .O(N__45314),
            .I(N__44900));
    InMux I__10432 (
            .O(N__45313),
            .I(N__44893));
    InMux I__10431 (
            .O(N__45312),
            .I(N__44893));
    InMux I__10430 (
            .O(N__45311),
            .I(N__44893));
    InMux I__10429 (
            .O(N__45310),
            .I(N__44886));
    InMux I__10428 (
            .O(N__45309),
            .I(N__44886));
    InMux I__10427 (
            .O(N__45308),
            .I(N__44886));
    InMux I__10426 (
            .O(N__45307),
            .I(N__44879));
    InMux I__10425 (
            .O(N__45304),
            .I(N__44879));
    InMux I__10424 (
            .O(N__45303),
            .I(N__44879));
    InMux I__10423 (
            .O(N__45302),
            .I(N__44872));
    InMux I__10422 (
            .O(N__45299),
            .I(N__44872));
    InMux I__10421 (
            .O(N__45298),
            .I(N__44872));
    InMux I__10420 (
            .O(N__45297),
            .I(N__44864));
    InMux I__10419 (
            .O(N__45296),
            .I(N__44864));
    InMux I__10418 (
            .O(N__45293),
            .I(N__44856));
    InMux I__10417 (
            .O(N__45292),
            .I(N__44849));
    InMux I__10416 (
            .O(N__45289),
            .I(N__44849));
    InMux I__10415 (
            .O(N__45286),
            .I(N__44849));
    InMux I__10414 (
            .O(N__45285),
            .I(N__44844));
    InMux I__10413 (
            .O(N__45284),
            .I(N__44844));
    InMux I__10412 (
            .O(N__45283),
            .I(N__44835));
    InMux I__10411 (
            .O(N__45282),
            .I(N__44835));
    InMux I__10410 (
            .O(N__45281),
            .I(N__44835));
    InMux I__10409 (
            .O(N__45280),
            .I(N__44835));
    CascadeMux I__10408 (
            .O(N__45279),
            .I(N__44829));
    Span4Mux_v I__10407 (
            .O(N__45276),
            .I(N__44823));
    Span4Mux_v I__10406 (
            .O(N__45269),
            .I(N__44823));
    LocalMux I__10405 (
            .O(N__45262),
            .I(N__44812));
    LocalMux I__10404 (
            .O(N__45251),
            .I(N__44812));
    LocalMux I__10403 (
            .O(N__45244),
            .I(N__44812));
    LocalMux I__10402 (
            .O(N__45239),
            .I(N__44812));
    LocalMux I__10401 (
            .O(N__45232),
            .I(N__44812));
    InMux I__10400 (
            .O(N__45231),
            .I(N__44805));
    InMux I__10399 (
            .O(N__45228),
            .I(N__44805));
    InMux I__10398 (
            .O(N__45227),
            .I(N__44805));
    InMux I__10397 (
            .O(N__45224),
            .I(N__44794));
    InMux I__10396 (
            .O(N__45223),
            .I(N__44794));
    InMux I__10395 (
            .O(N__45220),
            .I(N__44794));
    InMux I__10394 (
            .O(N__45219),
            .I(N__44794));
    InMux I__10393 (
            .O(N__45218),
            .I(N__44794));
    LocalMux I__10392 (
            .O(N__45211),
            .I(N__44791));
    LocalMux I__10391 (
            .O(N__45206),
            .I(N__44774));
    LocalMux I__10390 (
            .O(N__45197),
            .I(N__44774));
    LocalMux I__10389 (
            .O(N__45190),
            .I(N__44774));
    LocalMux I__10388 (
            .O(N__45183),
            .I(N__44774));
    LocalMux I__10387 (
            .O(N__45174),
            .I(N__44774));
    LocalMux I__10386 (
            .O(N__45163),
            .I(N__44774));
    LocalMux I__10385 (
            .O(N__45152),
            .I(N__44774));
    LocalMux I__10384 (
            .O(N__45145),
            .I(N__44774));
    LocalMux I__10383 (
            .O(N__45142),
            .I(N__44771));
    InMux I__10382 (
            .O(N__45141),
            .I(N__44762));
    InMux I__10381 (
            .O(N__45140),
            .I(N__44762));
    InMux I__10380 (
            .O(N__45139),
            .I(N__44762));
    InMux I__10379 (
            .O(N__45138),
            .I(N__44762));
    InMux I__10378 (
            .O(N__45137),
            .I(N__44753));
    InMux I__10377 (
            .O(N__45136),
            .I(N__44753));
    InMux I__10376 (
            .O(N__45135),
            .I(N__44753));
    InMux I__10375 (
            .O(N__45134),
            .I(N__44753));
    LocalMux I__10374 (
            .O(N__45131),
            .I(N__44748));
    LocalMux I__10373 (
            .O(N__45128),
            .I(N__44748));
    Span4Mux_s1_h I__10372 (
            .O(N__45123),
            .I(N__44743));
    LocalMux I__10371 (
            .O(N__45116),
            .I(N__44743));
    LocalMux I__10370 (
            .O(N__45105),
            .I(N__44740));
    InMux I__10369 (
            .O(N__45104),
            .I(N__44737));
    InMux I__10368 (
            .O(N__45101),
            .I(N__44730));
    InMux I__10367 (
            .O(N__45100),
            .I(N__44730));
    InMux I__10366 (
            .O(N__45099),
            .I(N__44730));
    InMux I__10365 (
            .O(N__45098),
            .I(N__44723));
    InMux I__10364 (
            .O(N__45097),
            .I(N__44723));
    InMux I__10363 (
            .O(N__45096),
            .I(N__44723));
    CascadeMux I__10362 (
            .O(N__45095),
            .I(N__44719));
    CascadeMux I__10361 (
            .O(N__45094),
            .I(N__44711));
    CascadeMux I__10360 (
            .O(N__45093),
            .I(N__44707));
    InMux I__10359 (
            .O(N__45092),
            .I(N__44699));
    InMux I__10358 (
            .O(N__45091),
            .I(N__44699));
    InMux I__10357 (
            .O(N__45090),
            .I(N__44699));
    Span4Mux_h I__10356 (
            .O(N__45087),
            .I(N__44692));
    Span4Mux_v I__10355 (
            .O(N__45082),
            .I(N__44692));
    Span4Mux_h I__10354 (
            .O(N__45079),
            .I(N__44692));
    Span4Mux_h I__10353 (
            .O(N__45074),
            .I(N__44685));
    LocalMux I__10352 (
            .O(N__45067),
            .I(N__44685));
    LocalMux I__10351 (
            .O(N__45060),
            .I(N__44685));
    LocalMux I__10350 (
            .O(N__45053),
            .I(N__44678));
    LocalMux I__10349 (
            .O(N__45046),
            .I(N__44678));
    LocalMux I__10348 (
            .O(N__45037),
            .I(N__44678));
    InMux I__10347 (
            .O(N__45036),
            .I(N__44671));
    InMux I__10346 (
            .O(N__45033),
            .I(N__44671));
    InMux I__10345 (
            .O(N__45030),
            .I(N__44671));
    CascadeMux I__10344 (
            .O(N__45029),
            .I(N__44667));
    InMux I__10343 (
            .O(N__45028),
            .I(N__44656));
    InMux I__10342 (
            .O(N__45027),
            .I(N__44656));
    InMux I__10341 (
            .O(N__45026),
            .I(N__44656));
    InMux I__10340 (
            .O(N__45025),
            .I(N__44656));
    InMux I__10339 (
            .O(N__45024),
            .I(N__44649));
    InMux I__10338 (
            .O(N__45023),
            .I(N__44649));
    InMux I__10337 (
            .O(N__45020),
            .I(N__44649));
    CascadeMux I__10336 (
            .O(N__45019),
            .I(N__44646));
    InMux I__10335 (
            .O(N__45018),
            .I(N__44637));
    InMux I__10334 (
            .O(N__45017),
            .I(N__44637));
    InMux I__10333 (
            .O(N__45016),
            .I(N__44637));
    LocalMux I__10332 (
            .O(N__45007),
            .I(N__44625));
    LocalMux I__10331 (
            .O(N__45004),
            .I(N__44625));
    Span4Mux_h I__10330 (
            .O(N__44999),
            .I(N__44618));
    LocalMux I__10329 (
            .O(N__44990),
            .I(N__44618));
    LocalMux I__10328 (
            .O(N__44983),
            .I(N__44618));
    Span4Mux_s2_h I__10327 (
            .O(N__44980),
            .I(N__44611));
    LocalMux I__10326 (
            .O(N__44973),
            .I(N__44611));
    LocalMux I__10325 (
            .O(N__44962),
            .I(N__44611));
    InMux I__10324 (
            .O(N__44959),
            .I(N__44602));
    InMux I__10323 (
            .O(N__44958),
            .I(N__44602));
    InMux I__10322 (
            .O(N__44957),
            .I(N__44602));
    InMux I__10321 (
            .O(N__44956),
            .I(N__44602));
    CascadeMux I__10320 (
            .O(N__44955),
            .I(N__44597));
    Span4Mux_h I__10319 (
            .O(N__44950),
            .I(N__44589));
    Span4Mux_v I__10318 (
            .O(N__44941),
            .I(N__44589));
    LocalMux I__10317 (
            .O(N__44938),
            .I(N__44589));
    InMux I__10316 (
            .O(N__44937),
            .I(N__44582));
    InMux I__10315 (
            .O(N__44936),
            .I(N__44582));
    InMux I__10314 (
            .O(N__44935),
            .I(N__44582));
    InMux I__10313 (
            .O(N__44934),
            .I(N__44575));
    InMux I__10312 (
            .O(N__44933),
            .I(N__44575));
    InMux I__10311 (
            .O(N__44932),
            .I(N__44575));
    InMux I__10310 (
            .O(N__44931),
            .I(N__44568));
    InMux I__10309 (
            .O(N__44930),
            .I(N__44568));
    InMux I__10308 (
            .O(N__44929),
            .I(N__44568));
    InMux I__10307 (
            .O(N__44928),
            .I(N__44561));
    InMux I__10306 (
            .O(N__44927),
            .I(N__44561));
    InMux I__10305 (
            .O(N__44926),
            .I(N__44561));
    InMux I__10304 (
            .O(N__44925),
            .I(N__44554));
    InMux I__10303 (
            .O(N__44924),
            .I(N__44554));
    InMux I__10302 (
            .O(N__44923),
            .I(N__44554));
    Span4Mux_v I__10301 (
            .O(N__44918),
            .I(N__44547));
    LocalMux I__10300 (
            .O(N__44907),
            .I(N__44547));
    LocalMux I__10299 (
            .O(N__44900),
            .I(N__44547));
    LocalMux I__10298 (
            .O(N__44893),
            .I(N__44538));
    LocalMux I__10297 (
            .O(N__44886),
            .I(N__44538));
    LocalMux I__10296 (
            .O(N__44879),
            .I(N__44538));
    LocalMux I__10295 (
            .O(N__44872),
            .I(N__44538));
    InMux I__10294 (
            .O(N__44871),
            .I(N__44531));
    InMux I__10293 (
            .O(N__44870),
            .I(N__44531));
    InMux I__10292 (
            .O(N__44869),
            .I(N__44531));
    LocalMux I__10291 (
            .O(N__44864),
            .I(N__44528));
    InMux I__10290 (
            .O(N__44863),
            .I(N__44523));
    InMux I__10289 (
            .O(N__44862),
            .I(N__44523));
    InMux I__10288 (
            .O(N__44861),
            .I(N__44513));
    InMux I__10287 (
            .O(N__44860),
            .I(N__44513));
    InMux I__10286 (
            .O(N__44859),
            .I(N__44510));
    LocalMux I__10285 (
            .O(N__44856),
            .I(N__44507));
    LocalMux I__10284 (
            .O(N__44849),
            .I(N__44500));
    LocalMux I__10283 (
            .O(N__44844),
            .I(N__44500));
    LocalMux I__10282 (
            .O(N__44835),
            .I(N__44500));
    InMux I__10281 (
            .O(N__44834),
            .I(N__44495));
    InMux I__10280 (
            .O(N__44833),
            .I(N__44495));
    InMux I__10279 (
            .O(N__44832),
            .I(N__44492));
    InMux I__10278 (
            .O(N__44829),
            .I(N__44487));
    InMux I__10277 (
            .O(N__44828),
            .I(N__44487));
    Span4Mux_v I__10276 (
            .O(N__44823),
            .I(N__44474));
    Span4Mux_v I__10275 (
            .O(N__44812),
            .I(N__44474));
    LocalMux I__10274 (
            .O(N__44805),
            .I(N__44474));
    LocalMux I__10273 (
            .O(N__44794),
            .I(N__44474));
    Span4Mux_h I__10272 (
            .O(N__44791),
            .I(N__44463));
    Span4Mux_v I__10271 (
            .O(N__44774),
            .I(N__44463));
    Span4Mux_v I__10270 (
            .O(N__44771),
            .I(N__44463));
    LocalMux I__10269 (
            .O(N__44762),
            .I(N__44463));
    LocalMux I__10268 (
            .O(N__44753),
            .I(N__44463));
    Span4Mux_v I__10267 (
            .O(N__44748),
            .I(N__44450));
    Span4Mux_h I__10266 (
            .O(N__44743),
            .I(N__44450));
    Span4Mux_v I__10265 (
            .O(N__44740),
            .I(N__44450));
    LocalMux I__10264 (
            .O(N__44737),
            .I(N__44450));
    LocalMux I__10263 (
            .O(N__44730),
            .I(N__44450));
    LocalMux I__10262 (
            .O(N__44723),
            .I(N__44450));
    InMux I__10261 (
            .O(N__44722),
            .I(N__44441));
    InMux I__10260 (
            .O(N__44719),
            .I(N__44441));
    InMux I__10259 (
            .O(N__44718),
            .I(N__44441));
    InMux I__10258 (
            .O(N__44717),
            .I(N__44441));
    CascadeMux I__10257 (
            .O(N__44716),
            .I(N__44437));
    InMux I__10256 (
            .O(N__44715),
            .I(N__44426));
    InMux I__10255 (
            .O(N__44714),
            .I(N__44426));
    InMux I__10254 (
            .O(N__44711),
            .I(N__44426));
    InMux I__10253 (
            .O(N__44710),
            .I(N__44419));
    InMux I__10252 (
            .O(N__44707),
            .I(N__44419));
    InMux I__10251 (
            .O(N__44706),
            .I(N__44419));
    LocalMux I__10250 (
            .O(N__44699),
            .I(N__44416));
    Span4Mux_h I__10249 (
            .O(N__44692),
            .I(N__44407));
    Span4Mux_v I__10248 (
            .O(N__44685),
            .I(N__44407));
    Span4Mux_h I__10247 (
            .O(N__44678),
            .I(N__44407));
    LocalMux I__10246 (
            .O(N__44671),
            .I(N__44407));
    InMux I__10245 (
            .O(N__44670),
            .I(N__44398));
    InMux I__10244 (
            .O(N__44667),
            .I(N__44398));
    InMux I__10243 (
            .O(N__44666),
            .I(N__44398));
    InMux I__10242 (
            .O(N__44665),
            .I(N__44398));
    LocalMux I__10241 (
            .O(N__44656),
            .I(N__44393));
    LocalMux I__10240 (
            .O(N__44649),
            .I(N__44393));
    InMux I__10239 (
            .O(N__44646),
            .I(N__44386));
    InMux I__10238 (
            .O(N__44645),
            .I(N__44386));
    InMux I__10237 (
            .O(N__44644),
            .I(N__44386));
    LocalMux I__10236 (
            .O(N__44637),
            .I(N__44382));
    InMux I__10235 (
            .O(N__44636),
            .I(N__44375));
    InMux I__10234 (
            .O(N__44635),
            .I(N__44375));
    InMux I__10233 (
            .O(N__44634),
            .I(N__44375));
    InMux I__10232 (
            .O(N__44633),
            .I(N__44368));
    InMux I__10231 (
            .O(N__44632),
            .I(N__44368));
    InMux I__10230 (
            .O(N__44631),
            .I(N__44368));
    InMux I__10229 (
            .O(N__44630),
            .I(N__44365));
    Span4Mux_v I__10228 (
            .O(N__44625),
            .I(N__44360));
    Span4Mux_v I__10227 (
            .O(N__44618),
            .I(N__44360));
    Span4Mux_h I__10226 (
            .O(N__44611),
            .I(N__44355));
    LocalMux I__10225 (
            .O(N__44602),
            .I(N__44355));
    InMux I__10224 (
            .O(N__44601),
            .I(N__44346));
    InMux I__10223 (
            .O(N__44600),
            .I(N__44346));
    InMux I__10222 (
            .O(N__44597),
            .I(N__44346));
    InMux I__10221 (
            .O(N__44596),
            .I(N__44346));
    Span4Mux_v I__10220 (
            .O(N__44589),
            .I(N__44339));
    LocalMux I__10219 (
            .O(N__44582),
            .I(N__44339));
    LocalMux I__10218 (
            .O(N__44575),
            .I(N__44339));
    LocalMux I__10217 (
            .O(N__44568),
            .I(N__44332));
    LocalMux I__10216 (
            .O(N__44561),
            .I(N__44332));
    LocalMux I__10215 (
            .O(N__44554),
            .I(N__44332));
    Span4Mux_v I__10214 (
            .O(N__44547),
            .I(N__44325));
    Span4Mux_s2_h I__10213 (
            .O(N__44538),
            .I(N__44325));
    LocalMux I__10212 (
            .O(N__44531),
            .I(N__44325));
    Span4Mux_h I__10211 (
            .O(N__44528),
            .I(N__44320));
    LocalMux I__10210 (
            .O(N__44523),
            .I(N__44320));
    InMux I__10209 (
            .O(N__44522),
            .I(N__44313));
    InMux I__10208 (
            .O(N__44521),
            .I(N__44313));
    InMux I__10207 (
            .O(N__44520),
            .I(N__44313));
    InMux I__10206 (
            .O(N__44519),
            .I(N__44308));
    InMux I__10205 (
            .O(N__44518),
            .I(N__44308));
    LocalMux I__10204 (
            .O(N__44513),
            .I(N__44305));
    LocalMux I__10203 (
            .O(N__44510),
            .I(N__44302));
    Span4Mux_v I__10202 (
            .O(N__44507),
            .I(N__44291));
    Span4Mux_v I__10201 (
            .O(N__44500),
            .I(N__44291));
    LocalMux I__10200 (
            .O(N__44495),
            .I(N__44291));
    LocalMux I__10199 (
            .O(N__44492),
            .I(N__44291));
    LocalMux I__10198 (
            .O(N__44487),
            .I(N__44291));
    InMux I__10197 (
            .O(N__44486),
            .I(N__44288));
    InMux I__10196 (
            .O(N__44485),
            .I(N__44281));
    InMux I__10195 (
            .O(N__44484),
            .I(N__44281));
    InMux I__10194 (
            .O(N__44483),
            .I(N__44281));
    Span4Mux_h I__10193 (
            .O(N__44474),
            .I(N__44272));
    Span4Mux_h I__10192 (
            .O(N__44463),
            .I(N__44272));
    Span4Mux_h I__10191 (
            .O(N__44450),
            .I(N__44272));
    LocalMux I__10190 (
            .O(N__44441),
            .I(N__44272));
    InMux I__10189 (
            .O(N__44440),
            .I(N__44265));
    InMux I__10188 (
            .O(N__44437),
            .I(N__44265));
    InMux I__10187 (
            .O(N__44436),
            .I(N__44265));
    InMux I__10186 (
            .O(N__44435),
            .I(N__44258));
    InMux I__10185 (
            .O(N__44434),
            .I(N__44258));
    InMux I__10184 (
            .O(N__44433),
            .I(N__44258));
    LocalMux I__10183 (
            .O(N__44426),
            .I(N__44251));
    LocalMux I__10182 (
            .O(N__44419),
            .I(N__44251));
    Sp12to4 I__10181 (
            .O(N__44416),
            .I(N__44251));
    Span4Mux_v I__10180 (
            .O(N__44407),
            .I(N__44248));
    LocalMux I__10179 (
            .O(N__44398),
            .I(N__44245));
    Sp12to4 I__10178 (
            .O(N__44393),
            .I(N__44240));
    LocalMux I__10177 (
            .O(N__44386),
            .I(N__44240));
    InMux I__10176 (
            .O(N__44385),
            .I(N__44237));
    Span12Mux_s8_h I__10175 (
            .O(N__44382),
            .I(N__44228));
    LocalMux I__10174 (
            .O(N__44375),
            .I(N__44228));
    LocalMux I__10173 (
            .O(N__44368),
            .I(N__44228));
    LocalMux I__10172 (
            .O(N__44365),
            .I(N__44228));
    Span4Mux_h I__10171 (
            .O(N__44360),
            .I(N__44221));
    Span4Mux_h I__10170 (
            .O(N__44355),
            .I(N__44221));
    LocalMux I__10169 (
            .O(N__44346),
            .I(N__44221));
    Span4Mux_v I__10168 (
            .O(N__44339),
            .I(N__44208));
    Span4Mux_h I__10167 (
            .O(N__44332),
            .I(N__44208));
    Span4Mux_h I__10166 (
            .O(N__44325),
            .I(N__44208));
    Span4Mux_v I__10165 (
            .O(N__44320),
            .I(N__44208));
    LocalMux I__10164 (
            .O(N__44313),
            .I(N__44208));
    LocalMux I__10163 (
            .O(N__44308),
            .I(N__44208));
    Span4Mux_v I__10162 (
            .O(N__44305),
            .I(N__44203));
    Span4Mux_v I__10161 (
            .O(N__44302),
            .I(N__44203));
    Span4Mux_h I__10160 (
            .O(N__44291),
            .I(N__44196));
    LocalMux I__10159 (
            .O(N__44288),
            .I(N__44196));
    LocalMux I__10158 (
            .O(N__44281),
            .I(N__44196));
    Span4Mux_v I__10157 (
            .O(N__44272),
            .I(N__44189));
    LocalMux I__10156 (
            .O(N__44265),
            .I(N__44189));
    LocalMux I__10155 (
            .O(N__44258),
            .I(N__44189));
    Span12Mux_s10_h I__10154 (
            .O(N__44251),
            .I(N__44186));
    Span4Mux_v I__10153 (
            .O(N__44248),
            .I(N__44183));
    Span12Mux_v I__10152 (
            .O(N__44245),
            .I(N__44176));
    Span12Mux_v I__10151 (
            .O(N__44240),
            .I(N__44176));
    LocalMux I__10150 (
            .O(N__44237),
            .I(N__44176));
    Span12Mux_v I__10149 (
            .O(N__44228),
            .I(N__44173));
    Span4Mux_v I__10148 (
            .O(N__44221),
            .I(N__44168));
    Span4Mux_h I__10147 (
            .O(N__44208),
            .I(N__44168));
    Span4Mux_v I__10146 (
            .O(N__44203),
            .I(N__44161));
    Span4Mux_h I__10145 (
            .O(N__44196),
            .I(N__44161));
    Span4Mux_v I__10144 (
            .O(N__44189),
            .I(N__44161));
    Odrv12 I__10143 (
            .O(N__44186),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__10142 (
            .O(N__44183),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__10141 (
            .O(N__44176),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__10140 (
            .O(N__44173),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__10139 (
            .O(N__44168),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__10138 (
            .O(N__44161),
            .I(CONSTANT_ONE_NET));
    InMux I__10137 (
            .O(N__44148),
            .I(N__44144));
    InMux I__10136 (
            .O(N__44147),
            .I(N__44141));
    LocalMux I__10135 (
            .O(N__44144),
            .I(N__44138));
    LocalMux I__10134 (
            .O(N__44141),
            .I(N__44135));
    Odrv4 I__10133 (
            .O(N__44138),
            .I(\nx.n2291 ));
    Odrv4 I__10132 (
            .O(N__44135),
            .I(\nx.n2291 ));
    CascadeMux I__10131 (
            .O(N__44130),
            .I(N__44124));
    CascadeMux I__10130 (
            .O(N__44129),
            .I(N__44119));
    CascadeMux I__10129 (
            .O(N__44128),
            .I(N__44110));
    InMux I__10128 (
            .O(N__44127),
            .I(N__44106));
    InMux I__10127 (
            .O(N__44124),
            .I(N__44103));
    CascadeMux I__10126 (
            .O(N__44123),
            .I(N__44100));
    InMux I__10125 (
            .O(N__44122),
            .I(N__44091));
    InMux I__10124 (
            .O(N__44119),
            .I(N__44091));
    InMux I__10123 (
            .O(N__44118),
            .I(N__44091));
    CascadeMux I__10122 (
            .O(N__44117),
            .I(N__44087));
    CascadeMux I__10121 (
            .O(N__44116),
            .I(N__44083));
    InMux I__10120 (
            .O(N__44115),
            .I(N__44070));
    InMux I__10119 (
            .O(N__44114),
            .I(N__44070));
    InMux I__10118 (
            .O(N__44113),
            .I(N__44070));
    InMux I__10117 (
            .O(N__44110),
            .I(N__44070));
    InMux I__10116 (
            .O(N__44109),
            .I(N__44070));
    LocalMux I__10115 (
            .O(N__44106),
            .I(N__44067));
    LocalMux I__10114 (
            .O(N__44103),
            .I(N__44064));
    InMux I__10113 (
            .O(N__44100),
            .I(N__44061));
    InMux I__10112 (
            .O(N__44099),
            .I(N__44058));
    InMux I__10111 (
            .O(N__44098),
            .I(N__44055));
    LocalMux I__10110 (
            .O(N__44091),
            .I(N__44052));
    InMux I__10109 (
            .O(N__44090),
            .I(N__44045));
    InMux I__10108 (
            .O(N__44087),
            .I(N__44045));
    InMux I__10107 (
            .O(N__44086),
            .I(N__44045));
    InMux I__10106 (
            .O(N__44083),
            .I(N__44038));
    InMux I__10105 (
            .O(N__44082),
            .I(N__44038));
    InMux I__10104 (
            .O(N__44081),
            .I(N__44038));
    LocalMux I__10103 (
            .O(N__44070),
            .I(N__44035));
    Span4Mux_h I__10102 (
            .O(N__44067),
            .I(N__44026));
    Span4Mux_h I__10101 (
            .O(N__44064),
            .I(N__44026));
    LocalMux I__10100 (
            .O(N__44061),
            .I(N__44026));
    LocalMux I__10099 (
            .O(N__44058),
            .I(N__44026));
    LocalMux I__10098 (
            .O(N__44055),
            .I(\nx.n2324 ));
    Odrv4 I__10097 (
            .O(N__44052),
            .I(\nx.n2324 ));
    LocalMux I__10096 (
            .O(N__44045),
            .I(\nx.n2324 ));
    LocalMux I__10095 (
            .O(N__44038),
            .I(\nx.n2324 ));
    Odrv4 I__10094 (
            .O(N__44035),
            .I(\nx.n2324 ));
    Odrv4 I__10093 (
            .O(N__44026),
            .I(\nx.n2324 ));
    InMux I__10092 (
            .O(N__44013),
            .I(\nx.n10726 ));
    InMux I__10091 (
            .O(N__44010),
            .I(N__44007));
    LocalMux I__10090 (
            .O(N__44007),
            .I(N__44003));
    InMux I__10089 (
            .O(N__44006),
            .I(N__44000));
    Span4Mux_h I__10088 (
            .O(N__44003),
            .I(N__43997));
    LocalMux I__10087 (
            .O(N__44000),
            .I(N__43992));
    Span4Mux_h I__10086 (
            .O(N__43997),
            .I(N__43992));
    Odrv4 I__10085 (
            .O(N__43992),
            .I(\nx.n2390 ));
    InMux I__10084 (
            .O(N__43989),
            .I(\nx.n10711 ));
    CascadeMux I__10083 (
            .O(N__43986),
            .I(N__43982));
    CascadeMux I__10082 (
            .O(N__43985),
            .I(N__43979));
    InMux I__10081 (
            .O(N__43982),
            .I(N__43976));
    InMux I__10080 (
            .O(N__43979),
            .I(N__43972));
    LocalMux I__10079 (
            .O(N__43976),
            .I(N__43969));
    InMux I__10078 (
            .O(N__43975),
            .I(N__43966));
    LocalMux I__10077 (
            .O(N__43972),
            .I(N__43963));
    Odrv4 I__10076 (
            .O(N__43969),
            .I(\nx.n2305 ));
    LocalMux I__10075 (
            .O(N__43966),
            .I(\nx.n2305 ));
    Odrv4 I__10074 (
            .O(N__43963),
            .I(\nx.n2305 ));
    InMux I__10073 (
            .O(N__43956),
            .I(N__43953));
    LocalMux I__10072 (
            .O(N__43953),
            .I(N__43950));
    Span4Mux_h I__10071 (
            .O(N__43950),
            .I(N__43947));
    Odrv4 I__10070 (
            .O(N__43947),
            .I(\nx.n2372 ));
    InMux I__10069 (
            .O(N__43944),
            .I(\nx.n10712 ));
    InMux I__10068 (
            .O(N__43941),
            .I(N__43937));
    InMux I__10067 (
            .O(N__43940),
            .I(N__43933));
    LocalMux I__10066 (
            .O(N__43937),
            .I(N__43930));
    InMux I__10065 (
            .O(N__43936),
            .I(N__43927));
    LocalMux I__10064 (
            .O(N__43933),
            .I(N__43924));
    Odrv4 I__10063 (
            .O(N__43930),
            .I(\nx.n2304 ));
    LocalMux I__10062 (
            .O(N__43927),
            .I(\nx.n2304 ));
    Odrv12 I__10061 (
            .O(N__43924),
            .I(\nx.n2304 ));
    CascadeMux I__10060 (
            .O(N__43917),
            .I(N__43914));
    InMux I__10059 (
            .O(N__43914),
            .I(N__43911));
    LocalMux I__10058 (
            .O(N__43911),
            .I(N__43908));
    Span4Mux_h I__10057 (
            .O(N__43908),
            .I(N__43905));
    Odrv4 I__10056 (
            .O(N__43905),
            .I(\nx.n2371 ));
    InMux I__10055 (
            .O(N__43902),
            .I(\nx.n10713 ));
    InMux I__10054 (
            .O(N__43899),
            .I(N__43895));
    CascadeMux I__10053 (
            .O(N__43898),
            .I(N__43891));
    LocalMux I__10052 (
            .O(N__43895),
            .I(N__43888));
    InMux I__10051 (
            .O(N__43894),
            .I(N__43885));
    InMux I__10050 (
            .O(N__43891),
            .I(N__43882));
    Span4Mux_h I__10049 (
            .O(N__43888),
            .I(N__43879));
    LocalMux I__10048 (
            .O(N__43885),
            .I(\nx.n2303 ));
    LocalMux I__10047 (
            .O(N__43882),
            .I(\nx.n2303 ));
    Odrv4 I__10046 (
            .O(N__43879),
            .I(\nx.n2303 ));
    CascadeMux I__10045 (
            .O(N__43872),
            .I(N__43869));
    InMux I__10044 (
            .O(N__43869),
            .I(N__43866));
    LocalMux I__10043 (
            .O(N__43866),
            .I(\nx.n2370 ));
    InMux I__10042 (
            .O(N__43863),
            .I(\nx.n10714 ));
    CascadeMux I__10041 (
            .O(N__43860),
            .I(N__43857));
    InMux I__10040 (
            .O(N__43857),
            .I(N__43854));
    LocalMux I__10039 (
            .O(N__43854),
            .I(N__43849));
    InMux I__10038 (
            .O(N__43853),
            .I(N__43846));
    InMux I__10037 (
            .O(N__43852),
            .I(N__43843));
    Span4Mux_v I__10036 (
            .O(N__43849),
            .I(N__43840));
    LocalMux I__10035 (
            .O(N__43846),
            .I(\nx.n2302 ));
    LocalMux I__10034 (
            .O(N__43843),
            .I(\nx.n2302 ));
    Odrv4 I__10033 (
            .O(N__43840),
            .I(\nx.n2302 ));
    CascadeMux I__10032 (
            .O(N__43833),
            .I(N__43830));
    InMux I__10031 (
            .O(N__43830),
            .I(N__43827));
    LocalMux I__10030 (
            .O(N__43827),
            .I(N__43824));
    Span4Mux_h I__10029 (
            .O(N__43824),
            .I(N__43821));
    Odrv4 I__10028 (
            .O(N__43821),
            .I(\nx.n2369 ));
    InMux I__10027 (
            .O(N__43818),
            .I(bfn_15_24_0_));
    CascadeMux I__10026 (
            .O(N__43815),
            .I(N__43812));
    InMux I__10025 (
            .O(N__43812),
            .I(N__43807));
    CascadeMux I__10024 (
            .O(N__43811),
            .I(N__43804));
    InMux I__10023 (
            .O(N__43810),
            .I(N__43801));
    LocalMux I__10022 (
            .O(N__43807),
            .I(N__43798));
    InMux I__10021 (
            .O(N__43804),
            .I(N__43795));
    LocalMux I__10020 (
            .O(N__43801),
            .I(N__43792));
    Odrv4 I__10019 (
            .O(N__43798),
            .I(\nx.n2301 ));
    LocalMux I__10018 (
            .O(N__43795),
            .I(\nx.n2301 ));
    Odrv4 I__10017 (
            .O(N__43792),
            .I(\nx.n2301 ));
    InMux I__10016 (
            .O(N__43785),
            .I(N__43782));
    LocalMux I__10015 (
            .O(N__43782),
            .I(N__43779));
    Odrv4 I__10014 (
            .O(N__43779),
            .I(\nx.n2368 ));
    InMux I__10013 (
            .O(N__43776),
            .I(\nx.n10716 ));
    CascadeMux I__10012 (
            .O(N__43773),
            .I(N__43770));
    InMux I__10011 (
            .O(N__43770),
            .I(N__43767));
    LocalMux I__10010 (
            .O(N__43767),
            .I(N__43763));
    InMux I__10009 (
            .O(N__43766),
            .I(N__43760));
    Span4Mux_v I__10008 (
            .O(N__43763),
            .I(N__43757));
    LocalMux I__10007 (
            .O(N__43760),
            .I(\nx.n2300 ));
    Odrv4 I__10006 (
            .O(N__43757),
            .I(\nx.n2300 ));
    InMux I__10005 (
            .O(N__43752),
            .I(N__43749));
    LocalMux I__10004 (
            .O(N__43749),
            .I(N__43746));
    Span4Mux_h I__10003 (
            .O(N__43746),
            .I(N__43743));
    Odrv4 I__10002 (
            .O(N__43743),
            .I(\nx.n2367 ));
    InMux I__10001 (
            .O(N__43740),
            .I(\nx.n10717 ));
    CascadeMux I__10000 (
            .O(N__43737),
            .I(N__43734));
    InMux I__9999 (
            .O(N__43734),
            .I(N__43730));
    CascadeMux I__9998 (
            .O(N__43733),
            .I(N__43727));
    LocalMux I__9997 (
            .O(N__43730),
            .I(N__43723));
    InMux I__9996 (
            .O(N__43727),
            .I(N__43720));
    InMux I__9995 (
            .O(N__43726),
            .I(N__43717));
    Odrv4 I__9994 (
            .O(N__43723),
            .I(\nx.n2299 ));
    LocalMux I__9993 (
            .O(N__43720),
            .I(\nx.n2299 ));
    LocalMux I__9992 (
            .O(N__43717),
            .I(\nx.n2299 ));
    InMux I__9991 (
            .O(N__43710),
            .I(N__43707));
    LocalMux I__9990 (
            .O(N__43707),
            .I(N__43704));
    Odrv4 I__9989 (
            .O(N__43704),
            .I(\nx.n2366 ));
    InMux I__9988 (
            .O(N__43701),
            .I(\nx.n10718 ));
    CascadeMux I__9987 (
            .O(N__43698),
            .I(N__43695));
    InMux I__9986 (
            .O(N__43695),
            .I(N__43692));
    LocalMux I__9985 (
            .O(N__43692),
            .I(N__43689));
    Span4Mux_h I__9984 (
            .O(N__43689),
            .I(N__43685));
    CascadeMux I__9983 (
            .O(N__43688),
            .I(N__43682));
    Span4Mux_h I__9982 (
            .O(N__43685),
            .I(N__43679));
    InMux I__9981 (
            .O(N__43682),
            .I(N__43676));
    Odrv4 I__9980 (
            .O(N__43679),
            .I(\nx.n2400 ));
    LocalMux I__9979 (
            .O(N__43676),
            .I(\nx.n2400 ));
    CascadeMux I__9978 (
            .O(N__43671),
            .I(\nx.n2400_cascade_ ));
    InMux I__9977 (
            .O(N__43668),
            .I(N__43664));
    CascadeMux I__9976 (
            .O(N__43667),
            .I(N__43660));
    LocalMux I__9975 (
            .O(N__43664),
            .I(N__43657));
    InMux I__9974 (
            .O(N__43663),
            .I(N__43654));
    InMux I__9973 (
            .O(N__43660),
            .I(N__43651));
    Span4Mux_h I__9972 (
            .O(N__43657),
            .I(N__43648));
    LocalMux I__9971 (
            .O(N__43654),
            .I(\nx.n2403 ));
    LocalMux I__9970 (
            .O(N__43651),
            .I(\nx.n2403 ));
    Odrv4 I__9969 (
            .O(N__43648),
            .I(\nx.n2403 ));
    InMux I__9968 (
            .O(N__43641),
            .I(N__43638));
    LocalMux I__9967 (
            .O(N__43638),
            .I(N__43635));
    Span4Mux_h I__9966 (
            .O(N__43635),
            .I(N__43632));
    Span4Mux_h I__9965 (
            .O(N__43632),
            .I(N__43629));
    Odrv4 I__9964 (
            .O(N__43629),
            .I(\nx.n35_adj_658 ));
    CascadeMux I__9963 (
            .O(N__43626),
            .I(N__43623));
    InMux I__9962 (
            .O(N__43623),
            .I(N__43620));
    LocalMux I__9961 (
            .O(N__43620),
            .I(N__43617));
    Span4Mux_h I__9960 (
            .O(N__43617),
            .I(N__43612));
    InMux I__9959 (
            .O(N__43616),
            .I(N__43609));
    InMux I__9958 (
            .O(N__43615),
            .I(N__43606));
    Odrv4 I__9957 (
            .O(N__43612),
            .I(\nx.n2402 ));
    LocalMux I__9956 (
            .O(N__43609),
            .I(\nx.n2402 ));
    LocalMux I__9955 (
            .O(N__43606),
            .I(\nx.n2402 ));
    InMux I__9954 (
            .O(N__43599),
            .I(N__43596));
    LocalMux I__9953 (
            .O(N__43596),
            .I(N__43592));
    CascadeMux I__9952 (
            .O(N__43595),
            .I(N__43588));
    Span4Mux_h I__9951 (
            .O(N__43592),
            .I(N__43585));
    InMux I__9950 (
            .O(N__43591),
            .I(N__43582));
    InMux I__9949 (
            .O(N__43588),
            .I(N__43579));
    Odrv4 I__9948 (
            .O(N__43585),
            .I(\nx.n2406 ));
    LocalMux I__9947 (
            .O(N__43582),
            .I(\nx.n2406 ));
    LocalMux I__9946 (
            .O(N__43579),
            .I(\nx.n2406 ));
    InMux I__9945 (
            .O(N__43572),
            .I(N__43568));
    InMux I__9944 (
            .O(N__43571),
            .I(N__43564));
    LocalMux I__9943 (
            .O(N__43568),
            .I(N__43561));
    InMux I__9942 (
            .O(N__43567),
            .I(N__43558));
    LocalMux I__9941 (
            .O(N__43564),
            .I(N__43555));
    Span4Mux_v I__9940 (
            .O(N__43561),
            .I(N__43552));
    LocalMux I__9939 (
            .O(N__43558),
            .I(N__43549));
    Span4Mux_v I__9938 (
            .O(N__43555),
            .I(N__43545));
    Span4Mux_h I__9937 (
            .O(N__43552),
            .I(N__43540));
    Span4Mux_h I__9936 (
            .O(N__43549),
            .I(N__43540));
    InMux I__9935 (
            .O(N__43548),
            .I(N__43536));
    Span4Mux_h I__9934 (
            .O(N__43545),
            .I(N__43533));
    Span4Mux_h I__9933 (
            .O(N__43540),
            .I(N__43530));
    InMux I__9932 (
            .O(N__43539),
            .I(N__43527));
    LocalMux I__9931 (
            .O(N__43536),
            .I(N__43524));
    Span4Mux_h I__9930 (
            .O(N__43533),
            .I(N__43521));
    Span4Mux_h I__9929 (
            .O(N__43530),
            .I(N__43518));
    LocalMux I__9928 (
            .O(N__43527),
            .I(\nx.bit_ctr_12 ));
    Odrv4 I__9927 (
            .O(N__43524),
            .I(\nx.bit_ctr_12 ));
    Odrv4 I__9926 (
            .O(N__43521),
            .I(\nx.bit_ctr_12 ));
    Odrv4 I__9925 (
            .O(N__43518),
            .I(\nx.bit_ctr_12 ));
    InMux I__9924 (
            .O(N__43509),
            .I(N__43506));
    LocalMux I__9923 (
            .O(N__43506),
            .I(N__43503));
    Span4Mux_h I__9922 (
            .O(N__43503),
            .I(N__43500));
    Odrv4 I__9921 (
            .O(N__43500),
            .I(\nx.n2377 ));
    InMux I__9920 (
            .O(N__43497),
            .I(bfn_15_23_0_));
    CascadeMux I__9919 (
            .O(N__43494),
            .I(N__43491));
    InMux I__9918 (
            .O(N__43491),
            .I(N__43487));
    InMux I__9917 (
            .O(N__43490),
            .I(N__43483));
    LocalMux I__9916 (
            .O(N__43487),
            .I(N__43480));
    InMux I__9915 (
            .O(N__43486),
            .I(N__43477));
    LocalMux I__9914 (
            .O(N__43483),
            .I(\nx.n2309 ));
    Odrv4 I__9913 (
            .O(N__43480),
            .I(\nx.n2309 ));
    LocalMux I__9912 (
            .O(N__43477),
            .I(\nx.n2309 ));
    CascadeMux I__9911 (
            .O(N__43470),
            .I(N__43467));
    InMux I__9910 (
            .O(N__43467),
            .I(N__43464));
    LocalMux I__9909 (
            .O(N__43464),
            .I(N__43461));
    Span4Mux_v I__9908 (
            .O(N__43461),
            .I(N__43458));
    Odrv4 I__9907 (
            .O(N__43458),
            .I(\nx.n2376 ));
    InMux I__9906 (
            .O(N__43455),
            .I(\nx.n10708 ));
    CascadeMux I__9905 (
            .O(N__43452),
            .I(N__43448));
    CascadeMux I__9904 (
            .O(N__43451),
            .I(N__43444));
    InMux I__9903 (
            .O(N__43448),
            .I(N__43441));
    InMux I__9902 (
            .O(N__43447),
            .I(N__43438));
    InMux I__9901 (
            .O(N__43444),
            .I(N__43435));
    LocalMux I__9900 (
            .O(N__43441),
            .I(N__43432));
    LocalMux I__9899 (
            .O(N__43438),
            .I(\nx.n2308 ));
    LocalMux I__9898 (
            .O(N__43435),
            .I(\nx.n2308 ));
    Odrv4 I__9897 (
            .O(N__43432),
            .I(\nx.n2308 ));
    InMux I__9896 (
            .O(N__43425),
            .I(N__43422));
    LocalMux I__9895 (
            .O(N__43422),
            .I(N__43419));
    Span4Mux_h I__9894 (
            .O(N__43419),
            .I(N__43416));
    Odrv4 I__9893 (
            .O(N__43416),
            .I(\nx.n2375 ));
    InMux I__9892 (
            .O(N__43413),
            .I(\nx.n10709 ));
    InMux I__9891 (
            .O(N__43410),
            .I(N__43406));
    CascadeMux I__9890 (
            .O(N__43409),
            .I(N__43403));
    LocalMux I__9889 (
            .O(N__43406),
            .I(N__43400));
    InMux I__9888 (
            .O(N__43403),
            .I(N__43396));
    Span4Mux_h I__9887 (
            .O(N__43400),
            .I(N__43393));
    InMux I__9886 (
            .O(N__43399),
            .I(N__43390));
    LocalMux I__9885 (
            .O(N__43396),
            .I(N__43387));
    Odrv4 I__9884 (
            .O(N__43393),
            .I(\nx.n2307 ));
    LocalMux I__9883 (
            .O(N__43390),
            .I(\nx.n2307 ));
    Odrv12 I__9882 (
            .O(N__43387),
            .I(\nx.n2307 ));
    InMux I__9881 (
            .O(N__43380),
            .I(N__43377));
    LocalMux I__9880 (
            .O(N__43377),
            .I(\nx.n2374 ));
    InMux I__9879 (
            .O(N__43374),
            .I(\nx.n10710 ));
    CascadeMux I__9878 (
            .O(N__43371),
            .I(N__43366));
    InMux I__9877 (
            .O(N__43370),
            .I(N__43361));
    InMux I__9876 (
            .O(N__43369),
            .I(N__43361));
    InMux I__9875 (
            .O(N__43366),
            .I(N__43358));
    LocalMux I__9874 (
            .O(N__43361),
            .I(\nx.n2306 ));
    LocalMux I__9873 (
            .O(N__43358),
            .I(\nx.n2306 ));
    InMux I__9872 (
            .O(N__43353),
            .I(N__43350));
    LocalMux I__9871 (
            .O(N__43350),
            .I(N__43347));
    Span4Mux_h I__9870 (
            .O(N__43347),
            .I(N__43344));
    Odrv4 I__9869 (
            .O(N__43344),
            .I(\nx.n2373 ));
    CascadeMux I__9868 (
            .O(N__43341),
            .I(n19_adj_735_cascade_));
    InMux I__9867 (
            .O(N__43338),
            .I(N__43335));
    LocalMux I__9866 (
            .O(N__43335),
            .I(n13141));
    CascadeMux I__9865 (
            .O(N__43332),
            .I(N__43329));
    InMux I__9864 (
            .O(N__43329),
            .I(N__43326));
    LocalMux I__9863 (
            .O(N__43326),
            .I(n1));
    InMux I__9862 (
            .O(N__43323),
            .I(N__43320));
    LocalMux I__9861 (
            .O(N__43320),
            .I(N__43315));
    InMux I__9860 (
            .O(N__43319),
            .I(N__43312));
    InMux I__9859 (
            .O(N__43318),
            .I(N__43309));
    Span4Mux_v I__9858 (
            .O(N__43315),
            .I(N__43304));
    LocalMux I__9857 (
            .O(N__43312),
            .I(N__43304));
    LocalMux I__9856 (
            .O(N__43309),
            .I(n8_adj_747));
    Odrv4 I__9855 (
            .O(N__43304),
            .I(n8_adj_747));
    CascadeMux I__9854 (
            .O(N__43299),
            .I(N__43296));
    InMux I__9853 (
            .O(N__43296),
            .I(N__43290));
    InMux I__9852 (
            .O(N__43295),
            .I(N__43286));
    InMux I__9851 (
            .O(N__43294),
            .I(N__43283));
    InMux I__9850 (
            .O(N__43293),
            .I(N__43280));
    LocalMux I__9849 (
            .O(N__43290),
            .I(N__43277));
    InMux I__9848 (
            .O(N__43289),
            .I(N__43274));
    LocalMux I__9847 (
            .O(N__43286),
            .I(N__43269));
    LocalMux I__9846 (
            .O(N__43283),
            .I(N__43269));
    LocalMux I__9845 (
            .O(N__43280),
            .I(N__43266));
    Span4Mux_v I__9844 (
            .O(N__43277),
            .I(N__43259));
    LocalMux I__9843 (
            .O(N__43274),
            .I(N__43259));
    Span4Mux_v I__9842 (
            .O(N__43269),
            .I(N__43259));
    Span4Mux_v I__9841 (
            .O(N__43266),
            .I(N__43256));
    Odrv4 I__9840 (
            .O(N__43259),
            .I(n9426));
    Odrv4 I__9839 (
            .O(N__43256),
            .I(n9426));
    InMux I__9838 (
            .O(N__43251),
            .I(N__43245));
    InMux I__9837 (
            .O(N__43250),
            .I(N__43245));
    LocalMux I__9836 (
            .O(N__43245),
            .I(N__43242));
    Span4Mux_v I__9835 (
            .O(N__43242),
            .I(N__43239));
    Odrv4 I__9834 (
            .O(N__43239),
            .I(n6178));
    CascadeMux I__9833 (
            .O(N__43236),
            .I(n7310_cascade_));
    InMux I__9832 (
            .O(N__43233),
            .I(N__43229));
    InMux I__9831 (
            .O(N__43232),
            .I(N__43225));
    LocalMux I__9830 (
            .O(N__43229),
            .I(N__43222));
    CascadeMux I__9829 (
            .O(N__43228),
            .I(N__43219));
    LocalMux I__9828 (
            .O(N__43225),
            .I(N__43216));
    Span4Mux_h I__9827 (
            .O(N__43222),
            .I(N__43213));
    InMux I__9826 (
            .O(N__43219),
            .I(N__43210));
    Span4Mux_v I__9825 (
            .O(N__43216),
            .I(N__43207));
    Odrv4 I__9824 (
            .O(N__43213),
            .I(\nx.n2398 ));
    LocalMux I__9823 (
            .O(N__43210),
            .I(\nx.n2398 ));
    Odrv4 I__9822 (
            .O(N__43207),
            .I(\nx.n2398 ));
    InMux I__9821 (
            .O(N__43200),
            .I(N__43195));
    InMux I__9820 (
            .O(N__43199),
            .I(N__43192));
    CascadeMux I__9819 (
            .O(N__43198),
            .I(N__43189));
    LocalMux I__9818 (
            .O(N__43195),
            .I(N__43186));
    LocalMux I__9817 (
            .O(N__43192),
            .I(N__43183));
    InMux I__9816 (
            .O(N__43189),
            .I(N__43180));
    Span4Mux_v I__9815 (
            .O(N__43186),
            .I(N__43175));
    Span4Mux_h I__9814 (
            .O(N__43183),
            .I(N__43175));
    LocalMux I__9813 (
            .O(N__43180),
            .I(N__43170));
    Span4Mux_h I__9812 (
            .O(N__43175),
            .I(N__43170));
    Odrv4 I__9811 (
            .O(N__43170),
            .I(\nx.n2397 ));
    InMux I__9810 (
            .O(N__43167),
            .I(N__43164));
    LocalMux I__9809 (
            .O(N__43164),
            .I(N__43161));
    Span4Mux_v I__9808 (
            .O(N__43161),
            .I(N__43156));
    InMux I__9807 (
            .O(N__43160),
            .I(N__43153));
    InMux I__9806 (
            .O(N__43159),
            .I(N__43150));
    Span4Mux_h I__9805 (
            .O(N__43156),
            .I(N__43146));
    LocalMux I__9804 (
            .O(N__43153),
            .I(N__43143));
    LocalMux I__9803 (
            .O(N__43150),
            .I(N__43140));
    InMux I__9802 (
            .O(N__43149),
            .I(N__43137));
    Sp12to4 I__9801 (
            .O(N__43146),
            .I(N__43132));
    Span12Mux_v I__9800 (
            .O(N__43143),
            .I(N__43132));
    Odrv12 I__9799 (
            .O(N__43140),
            .I(neopxl_color_14));
    LocalMux I__9798 (
            .O(N__43137),
            .I(neopxl_color_14));
    Odrv12 I__9797 (
            .O(N__43132),
            .I(neopxl_color_14));
    CascadeMux I__9796 (
            .O(N__43125),
            .I(N__43122));
    InMux I__9795 (
            .O(N__43122),
            .I(N__43119));
    LocalMux I__9794 (
            .O(N__43119),
            .I(N__43116));
    Span4Mux_v I__9793 (
            .O(N__43116),
            .I(N__43113));
    Span4Mux_h I__9792 (
            .O(N__43113),
            .I(N__43110));
    Span4Mux_h I__9791 (
            .O(N__43110),
            .I(N__43107));
    Span4Mux_h I__9790 (
            .O(N__43107),
            .I(N__43104));
    Odrv4 I__9789 (
            .O(N__43104),
            .I(neopxl_color_prev_14));
    IoInMux I__9788 (
            .O(N__43101),
            .I(N__43098));
    LocalMux I__9787 (
            .O(N__43098),
            .I(N__43095));
    Span4Mux_s1_h I__9786 (
            .O(N__43095),
            .I(N__43092));
    Sp12to4 I__9785 (
            .O(N__43092),
            .I(N__43089));
    Span12Mux_v I__9784 (
            .O(N__43089),
            .I(N__43086));
    Span12Mux_h I__9783 (
            .O(N__43086),
            .I(N__43081));
    InMux I__9782 (
            .O(N__43085),
            .I(N__43078));
    InMux I__9781 (
            .O(N__43084),
            .I(N__43075));
    Odrv12 I__9780 (
            .O(N__43081),
            .I(pin_out_16));
    LocalMux I__9779 (
            .O(N__43078),
            .I(pin_out_16));
    LocalMux I__9778 (
            .O(N__43075),
            .I(pin_out_16));
    CascadeMux I__9777 (
            .O(N__43068),
            .I(n13438_cascade_));
    IoInMux I__9776 (
            .O(N__43065),
            .I(N__43062));
    LocalMux I__9775 (
            .O(N__43062),
            .I(N__43059));
    Span4Mux_s2_v I__9774 (
            .O(N__43059),
            .I(N__43056));
    Sp12to4 I__9773 (
            .O(N__43056),
            .I(N__43053));
    Span12Mux_s7_h I__9772 (
            .O(N__43053),
            .I(N__43049));
    InMux I__9771 (
            .O(N__43052),
            .I(N__43045));
    Span12Mux_v I__9770 (
            .O(N__43049),
            .I(N__43042));
    InMux I__9769 (
            .O(N__43048),
            .I(N__43039));
    LocalMux I__9768 (
            .O(N__43045),
            .I(N__43036));
    Odrv12 I__9767 (
            .O(N__43042),
            .I(pin_out_17));
    LocalMux I__9766 (
            .O(N__43039),
            .I(pin_out_17));
    Odrv4 I__9765 (
            .O(N__43036),
            .I(pin_out_17));
    CascadeMux I__9764 (
            .O(N__43029),
            .I(n13441_cascade_));
    CascadeMux I__9763 (
            .O(N__43026),
            .I(n13142_cascade_));
    InMux I__9762 (
            .O(N__43023),
            .I(N__43020));
    LocalMux I__9761 (
            .O(N__43020),
            .I(N__43017));
    Odrv4 I__9760 (
            .O(N__43017),
            .I(n13362));
    CascadeMux I__9759 (
            .O(N__43014),
            .I(n149_cascade_));
    IoInMux I__9758 (
            .O(N__43011),
            .I(N__43008));
    LocalMux I__9757 (
            .O(N__43008),
            .I(N__43005));
    IoSpan4Mux I__9756 (
            .O(N__43005),
            .I(N__43002));
    Span4Mux_s2_v I__9755 (
            .O(N__43002),
            .I(N__42999));
    Sp12to4 I__9754 (
            .O(N__42999),
            .I(N__42995));
    CascadeMux I__9753 (
            .O(N__42998),
            .I(N__42991));
    Span12Mux_v I__9752 (
            .O(N__42995),
            .I(N__42988));
    InMux I__9751 (
            .O(N__42994),
            .I(N__42983));
    InMux I__9750 (
            .O(N__42991),
            .I(N__42983));
    Odrv12 I__9749 (
            .O(N__42988),
            .I(pin_out_19));
    LocalMux I__9748 (
            .O(N__42983),
            .I(pin_out_19));
    InMux I__9747 (
            .O(N__42978),
            .I(N__42975));
    LocalMux I__9746 (
            .O(N__42975),
            .I(N__42969));
    InMux I__9745 (
            .O(N__42974),
            .I(N__42966));
    InMux I__9744 (
            .O(N__42973),
            .I(N__42963));
    InMux I__9743 (
            .O(N__42972),
            .I(N__42960));
    Span4Mux_v I__9742 (
            .O(N__42969),
            .I(N__42955));
    LocalMux I__9741 (
            .O(N__42966),
            .I(N__42955));
    LocalMux I__9740 (
            .O(N__42963),
            .I(n8_adj_746));
    LocalMux I__9739 (
            .O(N__42960),
            .I(n8_adj_746));
    Odrv4 I__9738 (
            .O(N__42955),
            .I(n8_adj_746));
    InMux I__9737 (
            .O(N__42948),
            .I(N__42942));
    InMux I__9736 (
            .O(N__42947),
            .I(N__42942));
    LocalMux I__9735 (
            .O(N__42942),
            .I(N__42939));
    Span4Mux_h I__9734 (
            .O(N__42939),
            .I(N__42936));
    Odrv4 I__9733 (
            .O(N__42936),
            .I(n6186));
    InMux I__9732 (
            .O(N__42933),
            .I(N__42930));
    LocalMux I__9731 (
            .O(N__42930),
            .I(n7326));
    InMux I__9730 (
            .O(N__42927),
            .I(N__42924));
    LocalMux I__9729 (
            .O(N__42924),
            .I(n11_adj_734));
    CascadeMux I__9728 (
            .O(N__42921),
            .I(n11_adj_734_cascade_));
    InMux I__9727 (
            .O(N__42918),
            .I(N__42915));
    LocalMux I__9726 (
            .O(N__42915),
            .I(N__42912));
    Odrv4 I__9725 (
            .O(N__42912),
            .I(n36_adj_773));
    IoInMux I__9724 (
            .O(N__42909),
            .I(N__42906));
    LocalMux I__9723 (
            .O(N__42906),
            .I(N__42903));
    Span4Mux_s2_v I__9722 (
            .O(N__42903),
            .I(N__42900));
    Span4Mux_v I__9721 (
            .O(N__42900),
            .I(N__42895));
    CascadeMux I__9720 (
            .O(N__42899),
            .I(N__42892));
    InMux I__9719 (
            .O(N__42898),
            .I(N__42889));
    Sp12to4 I__9718 (
            .O(N__42895),
            .I(N__42886));
    InMux I__9717 (
            .O(N__42892),
            .I(N__42883));
    LocalMux I__9716 (
            .O(N__42889),
            .I(N__42880));
    Span12Mux_h I__9715 (
            .O(N__42886),
            .I(N__42877));
    LocalMux I__9714 (
            .O(N__42883),
            .I(N__42872));
    Span4Mux_v I__9713 (
            .O(N__42880),
            .I(N__42872));
    Odrv12 I__9712 (
            .O(N__42877),
            .I(pin_out_21));
    Odrv4 I__9711 (
            .O(N__42872),
            .I(pin_out_21));
    IoInMux I__9710 (
            .O(N__42867),
            .I(N__42864));
    LocalMux I__9709 (
            .O(N__42864),
            .I(N__42860));
    CascadeMux I__9708 (
            .O(N__42863),
            .I(N__42857));
    Span12Mux_s6_v I__9707 (
            .O(N__42860),
            .I(N__42853));
    InMux I__9706 (
            .O(N__42857),
            .I(N__42850));
    InMux I__9705 (
            .O(N__42856),
            .I(N__42847));
    Span12Mux_h I__9704 (
            .O(N__42853),
            .I(N__42844));
    LocalMux I__9703 (
            .O(N__42850),
            .I(N__42841));
    LocalMux I__9702 (
            .O(N__42847),
            .I(N__42838));
    Odrv12 I__9701 (
            .O(N__42844),
            .I(pin_out_20));
    Odrv4 I__9700 (
            .O(N__42841),
            .I(pin_out_20));
    Odrv4 I__9699 (
            .O(N__42838),
            .I(pin_out_20));
    InMux I__9698 (
            .O(N__42831),
            .I(N__42827));
    InMux I__9697 (
            .O(N__42830),
            .I(N__42824));
    LocalMux I__9696 (
            .O(N__42827),
            .I(N__42821));
    LocalMux I__9695 (
            .O(N__42824),
            .I(N__42818));
    Span4Mux_v I__9694 (
            .O(N__42821),
            .I(N__42815));
    Span4Mux_v I__9693 (
            .O(N__42818),
            .I(N__42812));
    Odrv4 I__9692 (
            .O(N__42815),
            .I(n10_adj_736));
    Odrv4 I__9691 (
            .O(N__42812),
            .I(n10_adj_736));
    InMux I__9690 (
            .O(N__42807),
            .I(N__42804));
    LocalMux I__9689 (
            .O(N__42804),
            .I(N__42801));
    Span4Mux_v I__9688 (
            .O(N__42801),
            .I(N__42797));
    InMux I__9687 (
            .O(N__42800),
            .I(N__42794));
    Span4Mux_h I__9686 (
            .O(N__42797),
            .I(N__42791));
    LocalMux I__9685 (
            .O(N__42794),
            .I(N__42788));
    Sp12to4 I__9684 (
            .O(N__42791),
            .I(N__42785));
    Span12Mux_h I__9683 (
            .O(N__42788),
            .I(N__42782));
    Span12Mux_h I__9682 (
            .O(N__42785),
            .I(N__42779));
    Span12Mux_v I__9681 (
            .O(N__42782),
            .I(N__42776));
    Span12Mux_v I__9680 (
            .O(N__42779),
            .I(N__42771));
    Span12Mux_h I__9679 (
            .O(N__42776),
            .I(N__42771));
    Odrv12 I__9678 (
            .O(N__42771),
            .I(pin_in_14));
    CascadeMux I__9677 (
            .O(N__42768),
            .I(N__42762));
    InMux I__9676 (
            .O(N__42767),
            .I(N__42759));
    InMux I__9675 (
            .O(N__42766),
            .I(N__42756));
    InMux I__9674 (
            .O(N__42765),
            .I(N__42753));
    InMux I__9673 (
            .O(N__42762),
            .I(N__42750));
    LocalMux I__9672 (
            .O(N__42759),
            .I(N__42747));
    LocalMux I__9671 (
            .O(N__42756),
            .I(N__42742));
    LocalMux I__9670 (
            .O(N__42753),
            .I(N__42742));
    LocalMux I__9669 (
            .O(N__42750),
            .I(n7145));
    Odrv4 I__9668 (
            .O(N__42747),
            .I(n7145));
    Odrv4 I__9667 (
            .O(N__42742),
            .I(n7145));
    InMux I__9666 (
            .O(N__42735),
            .I(N__42732));
    LocalMux I__9665 (
            .O(N__42732),
            .I(N__42729));
    Odrv4 I__9664 (
            .O(N__42729),
            .I(n7314));
    InMux I__9663 (
            .O(N__42726),
            .I(N__42722));
    CascadeMux I__9662 (
            .O(N__42725),
            .I(N__42719));
    LocalMux I__9661 (
            .O(N__42722),
            .I(N__42716));
    InMux I__9660 (
            .O(N__42719),
            .I(N__42712));
    Span4Mux_h I__9659 (
            .O(N__42716),
            .I(N__42709));
    InMux I__9658 (
            .O(N__42715),
            .I(N__42706));
    LocalMux I__9657 (
            .O(N__42712),
            .I(N__42703));
    Span4Mux_h I__9656 (
            .O(N__42709),
            .I(N__42696));
    LocalMux I__9655 (
            .O(N__42706),
            .I(N__42696));
    Span4Mux_h I__9654 (
            .O(N__42703),
            .I(N__42693));
    CascadeMux I__9653 (
            .O(N__42702),
            .I(N__42690));
    CascadeMux I__9652 (
            .O(N__42701),
            .I(N__42687));
    Span4Mux_v I__9651 (
            .O(N__42696),
            .I(N__42684));
    Span4Mux_h I__9650 (
            .O(N__42693),
            .I(N__42681));
    InMux I__9649 (
            .O(N__42690),
            .I(N__42676));
    InMux I__9648 (
            .O(N__42687),
            .I(N__42676));
    Span4Mux_h I__9647 (
            .O(N__42684),
            .I(N__42673));
    Odrv4 I__9646 (
            .O(N__42681),
            .I(n6));
    LocalMux I__9645 (
            .O(N__42676),
            .I(n6));
    Odrv4 I__9644 (
            .O(N__42673),
            .I(n6));
    InMux I__9643 (
            .O(N__42666),
            .I(N__42660));
    InMux I__9642 (
            .O(N__42665),
            .I(N__42660));
    LocalMux I__9641 (
            .O(N__42660),
            .I(N__42657));
    Span4Mux_v I__9640 (
            .O(N__42657),
            .I(N__42654));
    Span4Mux_h I__9639 (
            .O(N__42654),
            .I(N__42651));
    Odrv4 I__9638 (
            .O(N__42651),
            .I(n6182));
    CascadeMux I__9637 (
            .O(N__42648),
            .I(n7318_cascade_));
    CascadeMux I__9636 (
            .O(N__42645),
            .I(N__42642));
    InMux I__9635 (
            .O(N__42642),
            .I(N__42637));
    CascadeMux I__9634 (
            .O(N__42641),
            .I(N__42634));
    InMux I__9633 (
            .O(N__42640),
            .I(N__42630));
    LocalMux I__9632 (
            .O(N__42637),
            .I(N__42627));
    InMux I__9631 (
            .O(N__42634),
            .I(N__42622));
    CascadeMux I__9630 (
            .O(N__42633),
            .I(N__42619));
    LocalMux I__9629 (
            .O(N__42630),
            .I(N__42614));
    Span4Mux_v I__9628 (
            .O(N__42627),
            .I(N__42614));
    CascadeMux I__9627 (
            .O(N__42626),
            .I(N__42611));
    InMux I__9626 (
            .O(N__42625),
            .I(N__42606));
    LocalMux I__9625 (
            .O(N__42622),
            .I(N__42603));
    InMux I__9624 (
            .O(N__42619),
            .I(N__42600));
    Span4Mux_h I__9623 (
            .O(N__42614),
            .I(N__42597));
    InMux I__9622 (
            .O(N__42611),
            .I(N__42594));
    InMux I__9621 (
            .O(N__42610),
            .I(N__42589));
    InMux I__9620 (
            .O(N__42609),
            .I(N__42589));
    LocalMux I__9619 (
            .O(N__42606),
            .I(n9_adj_733));
    Odrv4 I__9618 (
            .O(N__42603),
            .I(n9_adj_733));
    LocalMux I__9617 (
            .O(N__42600),
            .I(n9_adj_733));
    Odrv4 I__9616 (
            .O(N__42597),
            .I(n9_adj_733));
    LocalMux I__9615 (
            .O(N__42594),
            .I(n9_adj_733));
    LocalMux I__9614 (
            .O(N__42589),
            .I(n9_adj_733));
    CascadeMux I__9613 (
            .O(N__42576),
            .I(N__42572));
    InMux I__9612 (
            .O(N__42575),
            .I(N__42567));
    InMux I__9611 (
            .O(N__42572),
            .I(N__42567));
    LocalMux I__9610 (
            .O(N__42567),
            .I(N__42564));
    Odrv4 I__9609 (
            .O(N__42564),
            .I(n6188));
    InMux I__9608 (
            .O(N__42561),
            .I(N__42558));
    LocalMux I__9607 (
            .O(N__42558),
            .I(n7330));
    IoInMux I__9606 (
            .O(N__42555),
            .I(N__42552));
    LocalMux I__9605 (
            .O(N__42552),
            .I(N__42549));
    IoSpan4Mux I__9604 (
            .O(N__42549),
            .I(N__42546));
    Sp12to4 I__9603 (
            .O(N__42546),
            .I(N__42543));
    Span12Mux_v I__9602 (
            .O(N__42543),
            .I(N__42539));
    InMux I__9601 (
            .O(N__42542),
            .I(N__42535));
    Span12Mux_h I__9600 (
            .O(N__42539),
            .I(N__42532));
    InMux I__9599 (
            .O(N__42538),
            .I(N__42529));
    LocalMux I__9598 (
            .O(N__42535),
            .I(N__42526));
    Odrv12 I__9597 (
            .O(N__42532),
            .I(pin_out_18));
    LocalMux I__9596 (
            .O(N__42529),
            .I(pin_out_18));
    Odrv4 I__9595 (
            .O(N__42526),
            .I(pin_out_18));
    InMux I__9594 (
            .O(N__42519),
            .I(N__42513));
    InMux I__9593 (
            .O(N__42518),
            .I(N__42513));
    LocalMux I__9592 (
            .O(N__42513),
            .I(n6176));
    CascadeMux I__9591 (
            .O(N__42510),
            .I(n7306_cascade_));
    IoInMux I__9590 (
            .O(N__42507),
            .I(N__42504));
    LocalMux I__9589 (
            .O(N__42504),
            .I(N__42501));
    Span4Mux_s2_v I__9588 (
            .O(N__42501),
            .I(N__42498));
    Sp12to4 I__9587 (
            .O(N__42498),
            .I(N__42495));
    Span12Mux_s8_h I__9586 (
            .O(N__42495),
            .I(N__42491));
    CascadeMux I__9585 (
            .O(N__42494),
            .I(N__42488));
    Span12Mux_v I__9584 (
            .O(N__42491),
            .I(N__42484));
    InMux I__9583 (
            .O(N__42488),
            .I(N__42481));
    InMux I__9582 (
            .O(N__42487),
            .I(N__42478));
    Odrv12 I__9581 (
            .O(N__42484),
            .I(pin_out_9));
    LocalMux I__9580 (
            .O(N__42481),
            .I(pin_out_9));
    LocalMux I__9579 (
            .O(N__42478),
            .I(pin_out_9));
    InMux I__9578 (
            .O(N__42471),
            .I(N__42468));
    LocalMux I__9577 (
            .O(N__42468),
            .I(N__42465));
    Span4Mux_v I__9576 (
            .O(N__42465),
            .I(N__42462));
    Odrv4 I__9575 (
            .O(N__42462),
            .I(n13162));
    CascadeMux I__9574 (
            .O(N__42459),
            .I(n13161_cascade_));
    InMux I__9573 (
            .O(N__42456),
            .I(N__42451));
    InMux I__9572 (
            .O(N__42455),
            .I(N__42448));
    InMux I__9571 (
            .O(N__42454),
            .I(N__42445));
    LocalMux I__9570 (
            .O(N__42451),
            .I(N__42442));
    LocalMux I__9569 (
            .O(N__42448),
            .I(N__42439));
    LocalMux I__9568 (
            .O(N__42445),
            .I(N__42436));
    Span4Mux_h I__9567 (
            .O(N__42442),
            .I(N__42433));
    Odrv4 I__9566 (
            .O(N__42439),
            .I(n8_adj_751));
    Odrv4 I__9565 (
            .O(N__42436),
            .I(n8_adj_751));
    Odrv4 I__9564 (
            .O(N__42433),
            .I(n8_adj_751));
    InMux I__9563 (
            .O(N__42426),
            .I(N__42422));
    InMux I__9562 (
            .O(N__42425),
            .I(N__42419));
    LocalMux I__9561 (
            .O(N__42422),
            .I(n6164));
    LocalMux I__9560 (
            .O(N__42419),
            .I(n6164));
    CascadeMux I__9559 (
            .O(N__42414),
            .I(n7282_cascade_));
    IoInMux I__9558 (
            .O(N__42411),
            .I(N__42408));
    LocalMux I__9557 (
            .O(N__42408),
            .I(N__42405));
    Span12Mux_s4_v I__9556 (
            .O(N__42405),
            .I(N__42402));
    Span12Mux_v I__9555 (
            .O(N__42402),
            .I(N__42397));
    InMux I__9554 (
            .O(N__42401),
            .I(N__42392));
    InMux I__9553 (
            .O(N__42400),
            .I(N__42392));
    Odrv12 I__9552 (
            .O(N__42397),
            .I(pin_out_8));
    LocalMux I__9551 (
            .O(N__42392),
            .I(pin_out_8));
    CascadeMux I__9550 (
            .O(N__42387),
            .I(N__42383));
    InMux I__9549 (
            .O(N__42386),
            .I(N__42380));
    InMux I__9548 (
            .O(N__42383),
            .I(N__42377));
    LocalMux I__9547 (
            .O(N__42380),
            .I(n6184));
    LocalMux I__9546 (
            .O(N__42377),
            .I(n6184));
    CascadeMux I__9545 (
            .O(N__42372),
            .I(n7322_cascade_));
    InMux I__9544 (
            .O(N__42369),
            .I(N__42366));
    LocalMux I__9543 (
            .O(N__42366),
            .I(n13471));
    InMux I__9542 (
            .O(N__42363),
            .I(N__42360));
    LocalMux I__9541 (
            .O(N__42360),
            .I(N__42357));
    Odrv12 I__9540 (
            .O(N__42357),
            .I(n13465));
    CascadeMux I__9539 (
            .O(N__42354),
            .I(n13177_cascade_));
    IoInMux I__9538 (
            .O(N__42351),
            .I(N__42348));
    LocalMux I__9537 (
            .O(N__42348),
            .I(N__42345));
    Span4Mux_s0_v I__9536 (
            .O(N__42345),
            .I(N__42342));
    Sp12to4 I__9535 (
            .O(N__42342),
            .I(N__42339));
    Span12Mux_h I__9534 (
            .O(N__42339),
            .I(N__42336));
    Odrv12 I__9533 (
            .O(N__42336),
            .I(LED_c));
    InMux I__9532 (
            .O(N__42333),
            .I(N__42330));
    LocalMux I__9531 (
            .O(N__42330),
            .I(n13176));
    InMux I__9530 (
            .O(N__42327),
            .I(N__42321));
    InMux I__9529 (
            .O(N__42326),
            .I(N__42318));
    InMux I__9528 (
            .O(N__42325),
            .I(N__42315));
    InMux I__9527 (
            .O(N__42324),
            .I(N__42312));
    LocalMux I__9526 (
            .O(N__42321),
            .I(n21_adj_741));
    LocalMux I__9525 (
            .O(N__42318),
            .I(n21_adj_741));
    LocalMux I__9524 (
            .O(N__42315),
            .I(n21_adj_741));
    LocalMux I__9523 (
            .O(N__42312),
            .I(n21_adj_741));
    InMux I__9522 (
            .O(N__42303),
            .I(N__42300));
    LocalMux I__9521 (
            .O(N__42300),
            .I(n6172));
    InMux I__9520 (
            .O(N__42297),
            .I(N__42294));
    LocalMux I__9519 (
            .O(N__42294),
            .I(n7298));
    CascadeMux I__9518 (
            .O(N__42291),
            .I(n6172_cascade_));
    CascadeMux I__9517 (
            .O(N__42288),
            .I(N__42285));
    InMux I__9516 (
            .O(N__42285),
            .I(N__42281));
    InMux I__9515 (
            .O(N__42284),
            .I(N__42278));
    LocalMux I__9514 (
            .O(N__42281),
            .I(N__42275));
    LocalMux I__9513 (
            .O(N__42278),
            .I(n6174));
    Odrv12 I__9512 (
            .O(N__42275),
            .I(n6174));
    InMux I__9511 (
            .O(N__42270),
            .I(N__42267));
    LocalMux I__9510 (
            .O(N__42267),
            .I(n7302));
    CascadeMux I__9509 (
            .O(N__42264),
            .I(N__42257));
    CascadeMux I__9508 (
            .O(N__42263),
            .I(N__42253));
    InMux I__9507 (
            .O(N__42262),
            .I(N__42249));
    InMux I__9506 (
            .O(N__42261),
            .I(N__42246));
    InMux I__9505 (
            .O(N__42260),
            .I(N__42241));
    InMux I__9504 (
            .O(N__42257),
            .I(N__42241));
    InMux I__9503 (
            .O(N__42256),
            .I(N__42236));
    InMux I__9502 (
            .O(N__42253),
            .I(N__42236));
    InMux I__9501 (
            .O(N__42252),
            .I(N__42233));
    LocalMux I__9500 (
            .O(N__42249),
            .I(n7_adj_753));
    LocalMux I__9499 (
            .O(N__42246),
            .I(n7_adj_753));
    LocalMux I__9498 (
            .O(N__42241),
            .I(n7_adj_753));
    LocalMux I__9497 (
            .O(N__42236),
            .I(n7_adj_753));
    LocalMux I__9496 (
            .O(N__42233),
            .I(n7_adj_753));
    InMux I__9495 (
            .O(N__42222),
            .I(N__42219));
    LocalMux I__9494 (
            .O(N__42219),
            .I(N__42216));
    Odrv4 I__9493 (
            .O(N__42216),
            .I(\nx.n2271 ));
    CascadeMux I__9492 (
            .O(N__42213),
            .I(N__42210));
    InMux I__9491 (
            .O(N__42210),
            .I(N__42205));
    InMux I__9490 (
            .O(N__42209),
            .I(N__42202));
    InMux I__9489 (
            .O(N__42208),
            .I(N__42199));
    LocalMux I__9488 (
            .O(N__42205),
            .I(N__42194));
    LocalMux I__9487 (
            .O(N__42202),
            .I(N__42194));
    LocalMux I__9486 (
            .O(N__42199),
            .I(\nx.n2204 ));
    Odrv4 I__9485 (
            .O(N__42194),
            .I(\nx.n2204 ));
    InMux I__9484 (
            .O(N__42189),
            .I(N__42186));
    LocalMux I__9483 (
            .O(N__42186),
            .I(\nx.n2265 ));
    InMux I__9482 (
            .O(N__42183),
            .I(N__42179));
    CascadeMux I__9481 (
            .O(N__42182),
            .I(N__42176));
    LocalMux I__9480 (
            .O(N__42179),
            .I(N__42173));
    InMux I__9479 (
            .O(N__42176),
            .I(N__42170));
    Span4Mux_h I__9478 (
            .O(N__42173),
            .I(N__42164));
    LocalMux I__9477 (
            .O(N__42170),
            .I(N__42164));
    InMux I__9476 (
            .O(N__42169),
            .I(N__42161));
    Odrv4 I__9475 (
            .O(N__42164),
            .I(\nx.n2198 ));
    LocalMux I__9474 (
            .O(N__42161),
            .I(\nx.n2198 ));
    CascadeMux I__9473 (
            .O(N__42156),
            .I(\nx.n2297_cascade_ ));
    InMux I__9472 (
            .O(N__42153),
            .I(N__42150));
    LocalMux I__9471 (
            .O(N__42150),
            .I(N__42147));
    Odrv4 I__9470 (
            .O(N__42147),
            .I(\nx.n9650 ));
    InMux I__9469 (
            .O(N__42144),
            .I(N__42141));
    LocalMux I__9468 (
            .O(N__42141),
            .I(N__42138));
    Odrv4 I__9467 (
            .O(N__42138),
            .I(\nx.n31_adj_645 ));
    InMux I__9466 (
            .O(N__42135),
            .I(N__42132));
    LocalMux I__9465 (
            .O(N__42132),
            .I(\nx.n2269 ));
    CascadeMux I__9464 (
            .O(N__42129),
            .I(N__42125));
    InMux I__9463 (
            .O(N__42128),
            .I(N__42121));
    InMux I__9462 (
            .O(N__42125),
            .I(N__42118));
    CascadeMux I__9461 (
            .O(N__42124),
            .I(N__42115));
    LocalMux I__9460 (
            .O(N__42121),
            .I(N__42110));
    LocalMux I__9459 (
            .O(N__42118),
            .I(N__42110));
    InMux I__9458 (
            .O(N__42115),
            .I(N__42107));
    Span4Mux_h I__9457 (
            .O(N__42110),
            .I(N__42104));
    LocalMux I__9456 (
            .O(N__42107),
            .I(\nx.n2202 ));
    Odrv4 I__9455 (
            .O(N__42104),
            .I(\nx.n2202 ));
    InMux I__9454 (
            .O(N__42099),
            .I(N__42096));
    LocalMux I__9453 (
            .O(N__42096),
            .I(\nx.n2267 ));
    CascadeMux I__9452 (
            .O(N__42093),
            .I(N__42090));
    InMux I__9451 (
            .O(N__42090),
            .I(N__42086));
    CascadeMux I__9450 (
            .O(N__42089),
            .I(N__42083));
    LocalMux I__9449 (
            .O(N__42086),
            .I(N__42080));
    InMux I__9448 (
            .O(N__42083),
            .I(N__42077));
    Span4Mux_h I__9447 (
            .O(N__42080),
            .I(N__42071));
    LocalMux I__9446 (
            .O(N__42077),
            .I(N__42071));
    InMux I__9445 (
            .O(N__42076),
            .I(N__42068));
    Odrv4 I__9444 (
            .O(N__42071),
            .I(\nx.n2200 ));
    LocalMux I__9443 (
            .O(N__42068),
            .I(\nx.n2200 ));
    InMux I__9442 (
            .O(N__42063),
            .I(N__42060));
    LocalMux I__9441 (
            .O(N__42060),
            .I(\nx.n2266 ));
    InMux I__9440 (
            .O(N__42057),
            .I(N__42053));
    CascadeMux I__9439 (
            .O(N__42056),
            .I(N__42049));
    LocalMux I__9438 (
            .O(N__42053),
            .I(N__42046));
    InMux I__9437 (
            .O(N__42052),
            .I(N__42043));
    InMux I__9436 (
            .O(N__42049),
            .I(N__42040));
    Span4Mux_h I__9435 (
            .O(N__42046),
            .I(N__42035));
    LocalMux I__9434 (
            .O(N__42043),
            .I(N__42035));
    LocalMux I__9433 (
            .O(N__42040),
            .I(\nx.n2199 ));
    Odrv4 I__9432 (
            .O(N__42035),
            .I(\nx.n2199 ));
    InMux I__9431 (
            .O(N__42030),
            .I(N__42027));
    LocalMux I__9430 (
            .O(N__42027),
            .I(\nx.n2260 ));
    CascadeMux I__9429 (
            .O(N__42024),
            .I(N__42021));
    InMux I__9428 (
            .O(N__42021),
            .I(N__42017));
    CascadeMux I__9427 (
            .O(N__42020),
            .I(N__42014));
    LocalMux I__9426 (
            .O(N__42017),
            .I(N__42010));
    InMux I__9425 (
            .O(N__42014),
            .I(N__42007));
    CascadeMux I__9424 (
            .O(N__42013),
            .I(N__42004));
    Span4Mux_v I__9423 (
            .O(N__42010),
            .I(N__41999));
    LocalMux I__9422 (
            .O(N__42007),
            .I(N__41999));
    InMux I__9421 (
            .O(N__42004),
            .I(N__41996));
    Odrv4 I__9420 (
            .O(N__41999),
            .I(\nx.n2193 ));
    LocalMux I__9419 (
            .O(N__41996),
            .I(\nx.n2193 ));
    CascadeMux I__9418 (
            .O(N__41991),
            .I(N__41985));
    CascadeMux I__9417 (
            .O(N__41990),
            .I(N__41982));
    CascadeMux I__9416 (
            .O(N__41989),
            .I(N__41978));
    CascadeMux I__9415 (
            .O(N__41988),
            .I(N__41969));
    InMux I__9414 (
            .O(N__41985),
            .I(N__41958));
    InMux I__9413 (
            .O(N__41982),
            .I(N__41958));
    InMux I__9412 (
            .O(N__41981),
            .I(N__41958));
    InMux I__9411 (
            .O(N__41978),
            .I(N__41958));
    InMux I__9410 (
            .O(N__41977),
            .I(N__41958));
    CascadeMux I__9409 (
            .O(N__41976),
            .I(N__41954));
    InMux I__9408 (
            .O(N__41975),
            .I(N__41950));
    CascadeMux I__9407 (
            .O(N__41974),
            .I(N__41945));
    InMux I__9406 (
            .O(N__41973),
            .I(N__41940));
    InMux I__9405 (
            .O(N__41972),
            .I(N__41940));
    InMux I__9404 (
            .O(N__41969),
            .I(N__41937));
    LocalMux I__9403 (
            .O(N__41958),
            .I(N__41934));
    CascadeMux I__9402 (
            .O(N__41957),
            .I(N__41929));
    InMux I__9401 (
            .O(N__41954),
            .I(N__41923));
    InMux I__9400 (
            .O(N__41953),
            .I(N__41923));
    LocalMux I__9399 (
            .O(N__41950),
            .I(N__41920));
    InMux I__9398 (
            .O(N__41949),
            .I(N__41913));
    InMux I__9397 (
            .O(N__41948),
            .I(N__41913));
    InMux I__9396 (
            .O(N__41945),
            .I(N__41913));
    LocalMux I__9395 (
            .O(N__41940),
            .I(N__41910));
    LocalMux I__9394 (
            .O(N__41937),
            .I(N__41905));
    Span4Mux_h I__9393 (
            .O(N__41934),
            .I(N__41905));
    InMux I__9392 (
            .O(N__41933),
            .I(N__41896));
    InMux I__9391 (
            .O(N__41932),
            .I(N__41896));
    InMux I__9390 (
            .O(N__41929),
            .I(N__41896));
    InMux I__9389 (
            .O(N__41928),
            .I(N__41896));
    LocalMux I__9388 (
            .O(N__41923),
            .I(\nx.n2225 ));
    Odrv4 I__9387 (
            .O(N__41920),
            .I(\nx.n2225 ));
    LocalMux I__9386 (
            .O(N__41913),
            .I(\nx.n2225 ));
    Odrv4 I__9385 (
            .O(N__41910),
            .I(\nx.n2225 ));
    Odrv4 I__9384 (
            .O(N__41905),
            .I(\nx.n2225 ));
    LocalMux I__9383 (
            .O(N__41896),
            .I(\nx.n2225 ));
    InMux I__9382 (
            .O(N__41883),
            .I(N__41878));
    CascadeMux I__9381 (
            .O(N__41882),
            .I(N__41875));
    InMux I__9380 (
            .O(N__41881),
            .I(N__41872));
    LocalMux I__9379 (
            .O(N__41878),
            .I(N__41869));
    InMux I__9378 (
            .O(N__41875),
            .I(N__41866));
    LocalMux I__9377 (
            .O(N__41872),
            .I(N__41863));
    Span4Mux_h I__9376 (
            .O(N__41869),
            .I(N__41860));
    LocalMux I__9375 (
            .O(N__41866),
            .I(N__41857));
    Span4Mux_v I__9374 (
            .O(N__41863),
            .I(N__41852));
    Span4Mux_h I__9373 (
            .O(N__41860),
            .I(N__41852));
    Odrv4 I__9372 (
            .O(N__41857),
            .I(\nx.n2396 ));
    Odrv4 I__9371 (
            .O(N__41852),
            .I(\nx.n2396 ));
    CascadeMux I__9370 (
            .O(N__41847),
            .I(N__41844));
    InMux I__9369 (
            .O(N__41844),
            .I(N__41840));
    InMux I__9368 (
            .O(N__41843),
            .I(N__41837));
    LocalMux I__9367 (
            .O(N__41840),
            .I(N__41834));
    LocalMux I__9366 (
            .O(N__41837),
            .I(N__41829));
    Span4Mux_h I__9365 (
            .O(N__41834),
            .I(N__41829));
    Odrv4 I__9364 (
            .O(N__41829),
            .I(\nx.n2395 ));
    InMux I__9363 (
            .O(N__41826),
            .I(N__41823));
    LocalMux I__9362 (
            .O(N__41823),
            .I(N__41820));
    Span4Mux_h I__9361 (
            .O(N__41820),
            .I(N__41817));
    Odrv4 I__9360 (
            .O(N__41817),
            .I(\nx.n2462 ));
    InMux I__9359 (
            .O(N__41814),
            .I(\nx.n10741 ));
    CascadeMux I__9358 (
            .O(N__41811),
            .I(N__41808));
    InMux I__9357 (
            .O(N__41808),
            .I(N__41805));
    LocalMux I__9356 (
            .O(N__41805),
            .I(N__41801));
    InMux I__9355 (
            .O(N__41804),
            .I(N__41798));
    Span4Mux_v I__9354 (
            .O(N__41801),
            .I(N__41795));
    LocalMux I__9353 (
            .O(N__41798),
            .I(\nx.n2394 ));
    Odrv4 I__9352 (
            .O(N__41795),
            .I(\nx.n2394 ));
    InMux I__9351 (
            .O(N__41790),
            .I(N__41787));
    LocalMux I__9350 (
            .O(N__41787),
            .I(N__41784));
    Span4Mux_v I__9349 (
            .O(N__41784),
            .I(N__41781));
    Span4Mux_h I__9348 (
            .O(N__41781),
            .I(N__41778));
    Odrv4 I__9347 (
            .O(N__41778),
            .I(\nx.n2461 ));
    InMux I__9346 (
            .O(N__41775),
            .I(bfn_14_23_0_));
    CascadeMux I__9345 (
            .O(N__41772),
            .I(N__41769));
    InMux I__9344 (
            .O(N__41769),
            .I(N__41766));
    LocalMux I__9343 (
            .O(N__41766),
            .I(N__41761));
    InMux I__9342 (
            .O(N__41765),
            .I(N__41756));
    InMux I__9341 (
            .O(N__41764),
            .I(N__41756));
    Span4Mux_v I__9340 (
            .O(N__41761),
            .I(N__41753));
    LocalMux I__9339 (
            .O(N__41756),
            .I(\nx.n2393 ));
    Odrv4 I__9338 (
            .O(N__41753),
            .I(\nx.n2393 ));
    CascadeMux I__9337 (
            .O(N__41748),
            .I(N__41745));
    InMux I__9336 (
            .O(N__41745),
            .I(N__41742));
    LocalMux I__9335 (
            .O(N__41742),
            .I(N__41739));
    Span4Mux_h I__9334 (
            .O(N__41739),
            .I(N__41736));
    Odrv4 I__9333 (
            .O(N__41736),
            .I(\nx.n2460 ));
    InMux I__9332 (
            .O(N__41733),
            .I(\nx.n10743 ));
    CascadeMux I__9331 (
            .O(N__41730),
            .I(N__41727));
    InMux I__9330 (
            .O(N__41727),
            .I(N__41724));
    LocalMux I__9329 (
            .O(N__41724),
            .I(N__41719));
    InMux I__9328 (
            .O(N__41723),
            .I(N__41714));
    InMux I__9327 (
            .O(N__41722),
            .I(N__41714));
    Span4Mux_h I__9326 (
            .O(N__41719),
            .I(N__41711));
    LocalMux I__9325 (
            .O(N__41714),
            .I(N__41708));
    Odrv4 I__9324 (
            .O(N__41711),
            .I(\nx.n2392 ));
    Odrv4 I__9323 (
            .O(N__41708),
            .I(\nx.n2392 ));
    CascadeMux I__9322 (
            .O(N__41703),
            .I(N__41700));
    InMux I__9321 (
            .O(N__41700),
            .I(N__41697));
    LocalMux I__9320 (
            .O(N__41697),
            .I(N__41694));
    Span4Mux_v I__9319 (
            .O(N__41694),
            .I(N__41691));
    Odrv4 I__9318 (
            .O(N__41691),
            .I(\nx.n2459 ));
    InMux I__9317 (
            .O(N__41688),
            .I(\nx.n10744 ));
    InMux I__9316 (
            .O(N__41685),
            .I(N__41682));
    LocalMux I__9315 (
            .O(N__41682),
            .I(N__41679));
    Span4Mux_v I__9314 (
            .O(N__41679),
            .I(N__41676));
    Odrv4 I__9313 (
            .O(N__41676),
            .I(\nx.n2458 ));
    InMux I__9312 (
            .O(N__41673),
            .I(\nx.n10745 ));
    CascadeMux I__9311 (
            .O(N__41670),
            .I(N__41666));
    InMux I__9310 (
            .O(N__41669),
            .I(N__41657));
    InMux I__9309 (
            .O(N__41666),
            .I(N__41654));
    CascadeMux I__9308 (
            .O(N__41665),
            .I(N__41650));
    CascadeMux I__9307 (
            .O(N__41664),
            .I(N__41647));
    CascadeMux I__9306 (
            .O(N__41663),
            .I(N__41644));
    CascadeMux I__9305 (
            .O(N__41662),
            .I(N__41641));
    CascadeMux I__9304 (
            .O(N__41661),
            .I(N__41637));
    InMux I__9303 (
            .O(N__41660),
            .I(N__41632));
    LocalMux I__9302 (
            .O(N__41657),
            .I(N__41626));
    LocalMux I__9301 (
            .O(N__41654),
            .I(N__41626));
    InMux I__9300 (
            .O(N__41653),
            .I(N__41613));
    InMux I__9299 (
            .O(N__41650),
            .I(N__41613));
    InMux I__9298 (
            .O(N__41647),
            .I(N__41613));
    InMux I__9297 (
            .O(N__41644),
            .I(N__41613));
    InMux I__9296 (
            .O(N__41641),
            .I(N__41613));
    InMux I__9295 (
            .O(N__41640),
            .I(N__41613));
    InMux I__9294 (
            .O(N__41637),
            .I(N__41604));
    InMux I__9293 (
            .O(N__41636),
            .I(N__41604));
    InMux I__9292 (
            .O(N__41635),
            .I(N__41604));
    LocalMux I__9291 (
            .O(N__41632),
            .I(N__41601));
    CascadeMux I__9290 (
            .O(N__41631),
            .I(N__41595));
    Span4Mux_v I__9289 (
            .O(N__41626),
            .I(N__41588));
    LocalMux I__9288 (
            .O(N__41613),
            .I(N__41588));
    InMux I__9287 (
            .O(N__41612),
            .I(N__41585));
    InMux I__9286 (
            .O(N__41611),
            .I(N__41582));
    LocalMux I__9285 (
            .O(N__41604),
            .I(N__41577));
    Span4Mux_v I__9284 (
            .O(N__41601),
            .I(N__41577));
    InMux I__9283 (
            .O(N__41600),
            .I(N__41574));
    InMux I__9282 (
            .O(N__41599),
            .I(N__41567));
    InMux I__9281 (
            .O(N__41598),
            .I(N__41567));
    InMux I__9280 (
            .O(N__41595),
            .I(N__41567));
    InMux I__9279 (
            .O(N__41594),
            .I(N__41564));
    InMux I__9278 (
            .O(N__41593),
            .I(N__41561));
    Span4Mux_h I__9277 (
            .O(N__41588),
            .I(N__41558));
    LocalMux I__9276 (
            .O(N__41585),
            .I(\nx.n2423 ));
    LocalMux I__9275 (
            .O(N__41582),
            .I(\nx.n2423 ));
    Odrv4 I__9274 (
            .O(N__41577),
            .I(\nx.n2423 ));
    LocalMux I__9273 (
            .O(N__41574),
            .I(\nx.n2423 ));
    LocalMux I__9272 (
            .O(N__41567),
            .I(\nx.n2423 ));
    LocalMux I__9271 (
            .O(N__41564),
            .I(\nx.n2423 ));
    LocalMux I__9270 (
            .O(N__41561),
            .I(\nx.n2423 ));
    Odrv4 I__9269 (
            .O(N__41558),
            .I(\nx.n2423 ));
    InMux I__9268 (
            .O(N__41541),
            .I(\nx.n10746 ));
    InMux I__9267 (
            .O(N__41538),
            .I(N__41534));
    CascadeMux I__9266 (
            .O(N__41537),
            .I(N__41531));
    LocalMux I__9265 (
            .O(N__41534),
            .I(N__41528));
    InMux I__9264 (
            .O(N__41531),
            .I(N__41525));
    Span4Mux_h I__9263 (
            .O(N__41528),
            .I(N__41522));
    LocalMux I__9262 (
            .O(N__41525),
            .I(N__41519));
    Odrv4 I__9261 (
            .O(N__41522),
            .I(\nx.n2489 ));
    Odrv4 I__9260 (
            .O(N__41519),
            .I(\nx.n2489 ));
    InMux I__9259 (
            .O(N__41514),
            .I(N__41510));
    CascadeMux I__9258 (
            .O(N__41513),
            .I(N__41507));
    LocalMux I__9257 (
            .O(N__41510),
            .I(N__41503));
    InMux I__9256 (
            .O(N__41507),
            .I(N__41500));
    InMux I__9255 (
            .O(N__41506),
            .I(N__41497));
    Span4Mux_h I__9254 (
            .O(N__41503),
            .I(N__41492));
    LocalMux I__9253 (
            .O(N__41500),
            .I(N__41492));
    LocalMux I__9252 (
            .O(N__41497),
            .I(\nx.n2207 ));
    Odrv4 I__9251 (
            .O(N__41492),
            .I(\nx.n2207 ));
    CascadeMux I__9250 (
            .O(N__41487),
            .I(N__41484));
    InMux I__9249 (
            .O(N__41484),
            .I(N__41481));
    LocalMux I__9248 (
            .O(N__41481),
            .I(\nx.n2274 ));
    CascadeMux I__9247 (
            .O(N__41478),
            .I(N__41474));
    InMux I__9246 (
            .O(N__41477),
            .I(N__41468));
    InMux I__9245 (
            .O(N__41474),
            .I(N__41468));
    CascadeMux I__9244 (
            .O(N__41473),
            .I(N__41465));
    LocalMux I__9243 (
            .O(N__41468),
            .I(N__41462));
    InMux I__9242 (
            .O(N__41465),
            .I(N__41459));
    Span4Mux_h I__9241 (
            .O(N__41462),
            .I(N__41456));
    LocalMux I__9240 (
            .O(N__41459),
            .I(\nx.n2391 ));
    Odrv4 I__9239 (
            .O(N__41456),
            .I(\nx.n2391 ));
    InMux I__9238 (
            .O(N__41451),
            .I(N__41448));
    LocalMux I__9237 (
            .O(N__41448),
            .I(\nx.n2470 ));
    InMux I__9236 (
            .O(N__41445),
            .I(\nx.n10733 ));
    InMux I__9235 (
            .O(N__41442),
            .I(N__41439));
    LocalMux I__9234 (
            .O(N__41439),
            .I(N__41436));
    Span4Mux_v I__9233 (
            .O(N__41436),
            .I(N__41433));
    Odrv4 I__9232 (
            .O(N__41433),
            .I(\nx.n2469 ));
    InMux I__9231 (
            .O(N__41430),
            .I(bfn_14_22_0_));
    CascadeMux I__9230 (
            .O(N__41427),
            .I(N__41424));
    InMux I__9229 (
            .O(N__41424),
            .I(N__41419));
    CascadeMux I__9228 (
            .O(N__41423),
            .I(N__41416));
    CascadeMux I__9227 (
            .O(N__41422),
            .I(N__41413));
    LocalMux I__9226 (
            .O(N__41419),
            .I(N__41410));
    InMux I__9225 (
            .O(N__41416),
            .I(N__41407));
    InMux I__9224 (
            .O(N__41413),
            .I(N__41404));
    Span4Mux_h I__9223 (
            .O(N__41410),
            .I(N__41401));
    LocalMux I__9222 (
            .O(N__41407),
            .I(\nx.n2401 ));
    LocalMux I__9221 (
            .O(N__41404),
            .I(\nx.n2401 ));
    Odrv4 I__9220 (
            .O(N__41401),
            .I(\nx.n2401 ));
    InMux I__9219 (
            .O(N__41394),
            .I(N__41391));
    LocalMux I__9218 (
            .O(N__41391),
            .I(\nx.n2468 ));
    InMux I__9217 (
            .O(N__41388),
            .I(\nx.n10735 ));
    InMux I__9216 (
            .O(N__41385),
            .I(N__41382));
    LocalMux I__9215 (
            .O(N__41382),
            .I(N__41379));
    Span4Mux_h I__9214 (
            .O(N__41379),
            .I(N__41376));
    Span4Mux_h I__9213 (
            .O(N__41376),
            .I(N__41373));
    Odrv4 I__9212 (
            .O(N__41373),
            .I(\nx.n2467 ));
    InMux I__9211 (
            .O(N__41370),
            .I(\nx.n10736 ));
    CascadeMux I__9210 (
            .O(N__41367),
            .I(N__41363));
    InMux I__9209 (
            .O(N__41366),
            .I(N__41359));
    InMux I__9208 (
            .O(N__41363),
            .I(N__41356));
    InMux I__9207 (
            .O(N__41362),
            .I(N__41353));
    LocalMux I__9206 (
            .O(N__41359),
            .I(\nx.n2399 ));
    LocalMux I__9205 (
            .O(N__41356),
            .I(\nx.n2399 ));
    LocalMux I__9204 (
            .O(N__41353),
            .I(\nx.n2399 ));
    InMux I__9203 (
            .O(N__41346),
            .I(N__41343));
    LocalMux I__9202 (
            .O(N__41343),
            .I(N__41340));
    Odrv4 I__9201 (
            .O(N__41340),
            .I(\nx.n2466 ));
    InMux I__9200 (
            .O(N__41337),
            .I(\nx.n10737 ));
    CascadeMux I__9199 (
            .O(N__41334),
            .I(N__41331));
    InMux I__9198 (
            .O(N__41331),
            .I(N__41328));
    LocalMux I__9197 (
            .O(N__41328),
            .I(N__41325));
    Span4Mux_v I__9196 (
            .O(N__41325),
            .I(N__41322));
    Odrv4 I__9195 (
            .O(N__41322),
            .I(\nx.n2465 ));
    InMux I__9194 (
            .O(N__41319),
            .I(\nx.n10738 ));
    InMux I__9193 (
            .O(N__41316),
            .I(N__41313));
    LocalMux I__9192 (
            .O(N__41313),
            .I(N__41310));
    Span4Mux_h I__9191 (
            .O(N__41310),
            .I(N__41307));
    Odrv4 I__9190 (
            .O(N__41307),
            .I(\nx.n2464 ));
    InMux I__9189 (
            .O(N__41304),
            .I(\nx.n10739 ));
    CascadeMux I__9188 (
            .O(N__41301),
            .I(N__41298));
    InMux I__9187 (
            .O(N__41298),
            .I(N__41295));
    LocalMux I__9186 (
            .O(N__41295),
            .I(N__41292));
    Span4Mux_v I__9185 (
            .O(N__41292),
            .I(N__41289));
    Odrv4 I__9184 (
            .O(N__41289),
            .I(\nx.n2463 ));
    InMux I__9183 (
            .O(N__41286),
            .I(\nx.n10740 ));
    InMux I__9182 (
            .O(N__41283),
            .I(N__41280));
    LocalMux I__9181 (
            .O(N__41280),
            .I(N__41276));
    InMux I__9180 (
            .O(N__41279),
            .I(N__41272));
    Span4Mux_h I__9179 (
            .O(N__41276),
            .I(N__41269));
    InMux I__9178 (
            .O(N__41275),
            .I(N__41265));
    LocalMux I__9177 (
            .O(N__41272),
            .I(N__41262));
    Span4Mux_v I__9176 (
            .O(N__41269),
            .I(N__41259));
    CascadeMux I__9175 (
            .O(N__41268),
            .I(N__41255));
    LocalMux I__9174 (
            .O(N__41265),
            .I(N__41252));
    Span4Mux_v I__9173 (
            .O(N__41262),
            .I(N__41247));
    Span4Mux_h I__9172 (
            .O(N__41259),
            .I(N__41247));
    InMux I__9171 (
            .O(N__41258),
            .I(N__41244));
    InMux I__9170 (
            .O(N__41255),
            .I(N__41241));
    Span12Mux_v I__9169 (
            .O(N__41252),
            .I(N__41238));
    Span4Mux_h I__9168 (
            .O(N__41247),
            .I(N__41235));
    LocalMux I__9167 (
            .O(N__41244),
            .I(\nx.bit_ctr_11 ));
    LocalMux I__9166 (
            .O(N__41241),
            .I(\nx.bit_ctr_11 ));
    Odrv12 I__9165 (
            .O(N__41238),
            .I(\nx.bit_ctr_11 ));
    Odrv4 I__9164 (
            .O(N__41235),
            .I(\nx.bit_ctr_11 ));
    InMux I__9163 (
            .O(N__41226),
            .I(N__41223));
    LocalMux I__9162 (
            .O(N__41223),
            .I(N__41220));
    Sp12to4 I__9161 (
            .O(N__41220),
            .I(N__41217));
    Span12Mux_s11_v I__9160 (
            .O(N__41217),
            .I(N__41214));
    Odrv12 I__9159 (
            .O(N__41214),
            .I(\nx.n2477 ));
    InMux I__9158 (
            .O(N__41211),
            .I(bfn_14_21_0_));
    CascadeMux I__9157 (
            .O(N__41208),
            .I(N__41205));
    InMux I__9156 (
            .O(N__41205),
            .I(N__41200));
    CascadeMux I__9155 (
            .O(N__41204),
            .I(N__41197));
    CascadeMux I__9154 (
            .O(N__41203),
            .I(N__41194));
    LocalMux I__9153 (
            .O(N__41200),
            .I(N__41191));
    InMux I__9152 (
            .O(N__41197),
            .I(N__41188));
    InMux I__9151 (
            .O(N__41194),
            .I(N__41185));
    Span4Mux_h I__9150 (
            .O(N__41191),
            .I(N__41182));
    LocalMux I__9149 (
            .O(N__41188),
            .I(N__41179));
    LocalMux I__9148 (
            .O(N__41185),
            .I(N__41176));
    Span4Mux_h I__9147 (
            .O(N__41182),
            .I(N__41173));
    Span4Mux_h I__9146 (
            .O(N__41179),
            .I(N__41170));
    Odrv12 I__9145 (
            .O(N__41176),
            .I(\nx.n2409 ));
    Odrv4 I__9144 (
            .O(N__41173),
            .I(\nx.n2409 ));
    Odrv4 I__9143 (
            .O(N__41170),
            .I(\nx.n2409 ));
    InMux I__9142 (
            .O(N__41163),
            .I(N__41160));
    LocalMux I__9141 (
            .O(N__41160),
            .I(\nx.n2476 ));
    InMux I__9140 (
            .O(N__41157),
            .I(\nx.n10727 ));
    CascadeMux I__9139 (
            .O(N__41154),
            .I(N__41150));
    InMux I__9138 (
            .O(N__41153),
            .I(N__41147));
    InMux I__9137 (
            .O(N__41150),
            .I(N__41143));
    LocalMux I__9136 (
            .O(N__41147),
            .I(N__41140));
    CascadeMux I__9135 (
            .O(N__41146),
            .I(N__41137));
    LocalMux I__9134 (
            .O(N__41143),
            .I(N__41132));
    Span4Mux_h I__9133 (
            .O(N__41140),
            .I(N__41132));
    InMux I__9132 (
            .O(N__41137),
            .I(N__41129));
    Odrv4 I__9131 (
            .O(N__41132),
            .I(\nx.n2408 ));
    LocalMux I__9130 (
            .O(N__41129),
            .I(\nx.n2408 ));
    InMux I__9129 (
            .O(N__41124),
            .I(N__41121));
    LocalMux I__9128 (
            .O(N__41121),
            .I(N__41118));
    Span4Mux_h I__9127 (
            .O(N__41118),
            .I(N__41115));
    Odrv4 I__9126 (
            .O(N__41115),
            .I(\nx.n2475 ));
    InMux I__9125 (
            .O(N__41112),
            .I(\nx.n10728 ));
    InMux I__9124 (
            .O(N__41109),
            .I(N__41105));
    CascadeMux I__9123 (
            .O(N__41108),
            .I(N__41101));
    LocalMux I__9122 (
            .O(N__41105),
            .I(N__41098));
    InMux I__9121 (
            .O(N__41104),
            .I(N__41095));
    InMux I__9120 (
            .O(N__41101),
            .I(N__41092));
    Odrv4 I__9119 (
            .O(N__41098),
            .I(\nx.n2407 ));
    LocalMux I__9118 (
            .O(N__41095),
            .I(\nx.n2407 ));
    LocalMux I__9117 (
            .O(N__41092),
            .I(\nx.n2407 ));
    InMux I__9116 (
            .O(N__41085),
            .I(N__41082));
    LocalMux I__9115 (
            .O(N__41082),
            .I(\nx.n2474 ));
    InMux I__9114 (
            .O(N__41079),
            .I(\nx.n10729 ));
    InMux I__9113 (
            .O(N__41076),
            .I(N__41073));
    LocalMux I__9112 (
            .O(N__41073),
            .I(N__41070));
    Span4Mux_h I__9111 (
            .O(N__41070),
            .I(N__41067));
    Odrv4 I__9110 (
            .O(N__41067),
            .I(\nx.n2473 ));
    InMux I__9109 (
            .O(N__41064),
            .I(\nx.n10730 ));
    InMux I__9108 (
            .O(N__41061),
            .I(N__41056));
    InMux I__9107 (
            .O(N__41060),
            .I(N__41053));
    CascadeMux I__9106 (
            .O(N__41059),
            .I(N__41050));
    LocalMux I__9105 (
            .O(N__41056),
            .I(N__41047));
    LocalMux I__9104 (
            .O(N__41053),
            .I(N__41044));
    InMux I__9103 (
            .O(N__41050),
            .I(N__41041));
    Span4Mux_v I__9102 (
            .O(N__41047),
            .I(N__41036));
    Span4Mux_h I__9101 (
            .O(N__41044),
            .I(N__41036));
    LocalMux I__9100 (
            .O(N__41041),
            .I(\nx.n2405 ));
    Odrv4 I__9099 (
            .O(N__41036),
            .I(\nx.n2405 ));
    CascadeMux I__9098 (
            .O(N__41031),
            .I(N__41028));
    InMux I__9097 (
            .O(N__41028),
            .I(N__41025));
    LocalMux I__9096 (
            .O(N__41025),
            .I(N__41022));
    Span4Mux_h I__9095 (
            .O(N__41022),
            .I(N__41019));
    Odrv4 I__9094 (
            .O(N__41019),
            .I(\nx.n2472 ));
    InMux I__9093 (
            .O(N__41016),
            .I(\nx.n10731 ));
    CascadeMux I__9092 (
            .O(N__41013),
            .I(N__41009));
    InMux I__9091 (
            .O(N__41012),
            .I(N__41006));
    InMux I__9090 (
            .O(N__41009),
            .I(N__41003));
    LocalMux I__9089 (
            .O(N__41006),
            .I(\nx.n2404 ));
    LocalMux I__9088 (
            .O(N__41003),
            .I(\nx.n2404 ));
    InMux I__9087 (
            .O(N__40998),
            .I(N__40995));
    LocalMux I__9086 (
            .O(N__40995),
            .I(\nx.n2471 ));
    InMux I__9085 (
            .O(N__40992),
            .I(\nx.n10732 ));
    CascadeMux I__9084 (
            .O(N__40989),
            .I(n13474_cascade_));
    CascadeMux I__9083 (
            .O(N__40986),
            .I(N__40982));
    InMux I__9082 (
            .O(N__40985),
            .I(N__40979));
    InMux I__9081 (
            .O(N__40982),
            .I(N__40976));
    LocalMux I__9080 (
            .O(N__40979),
            .I(N__40971));
    LocalMux I__9079 (
            .O(N__40976),
            .I(N__40971));
    Span12Mux_v I__9078 (
            .O(N__40971),
            .I(N__40968));
    Span12Mux_v I__9077 (
            .O(N__40968),
            .I(N__40965));
    Span12Mux_h I__9076 (
            .O(N__40965),
            .I(N__40962));
    Odrv12 I__9075 (
            .O(N__40962),
            .I(pin_in_12));
    InMux I__9074 (
            .O(N__40959),
            .I(N__40956));
    LocalMux I__9073 (
            .O(N__40956),
            .I(n13477));
    InMux I__9072 (
            .O(N__40953),
            .I(N__40947));
    InMux I__9071 (
            .O(N__40952),
            .I(N__40947));
    LocalMux I__9070 (
            .O(N__40947),
            .I(N__40944));
    Span4Mux_v I__9069 (
            .O(N__40944),
            .I(N__40941));
    Sp12to4 I__9068 (
            .O(N__40941),
            .I(N__40938));
    Span12Mux_h I__9067 (
            .O(N__40938),
            .I(N__40935));
    Odrv12 I__9066 (
            .O(N__40935),
            .I(pin_in_13));
    CascadeMux I__9065 (
            .O(N__40932),
            .I(N__40929));
    InMux I__9064 (
            .O(N__40929),
            .I(N__40923));
    InMux I__9063 (
            .O(N__40928),
            .I(N__40923));
    LocalMux I__9062 (
            .O(N__40923),
            .I(N__40920));
    Span12Mux_v I__9061 (
            .O(N__40920),
            .I(N__40917));
    Span12Mux_h I__9060 (
            .O(N__40917),
            .I(N__40914));
    Odrv12 I__9059 (
            .O(N__40914),
            .I(pin_in_15));
    InMux I__9058 (
            .O(N__40911),
            .I(N__40908));
    LocalMux I__9057 (
            .O(N__40908),
            .I(n2367));
    InMux I__9056 (
            .O(N__40905),
            .I(N__40902));
    LocalMux I__9055 (
            .O(N__40902),
            .I(n33));
    CascadeMux I__9054 (
            .O(N__40899),
            .I(n2379_cascade_));
    InMux I__9053 (
            .O(N__40896),
            .I(N__40893));
    LocalMux I__9052 (
            .O(N__40893),
            .I(n45_adj_772));
    InMux I__9051 (
            .O(N__40890),
            .I(N__40880));
    InMux I__9050 (
            .O(N__40889),
            .I(N__40880));
    InMux I__9049 (
            .O(N__40888),
            .I(N__40880));
    InMux I__9048 (
            .O(N__40887),
            .I(N__40877));
    LocalMux I__9047 (
            .O(N__40880),
            .I(N__40874));
    LocalMux I__9046 (
            .O(N__40877),
            .I(N__40871));
    Span4Mux_h I__9045 (
            .O(N__40874),
            .I(N__40868));
    Span4Mux_v I__9044 (
            .O(N__40871),
            .I(N__40865));
    Span4Mux_h I__9043 (
            .O(N__40868),
            .I(N__40861));
    Span4Mux_v I__9042 (
            .O(N__40865),
            .I(N__40858));
    InMux I__9041 (
            .O(N__40864),
            .I(N__40855));
    Span4Mux_v I__9040 (
            .O(N__40861),
            .I(N__40852));
    Span4Mux_h I__9039 (
            .O(N__40858),
            .I(N__40849));
    LocalMux I__9038 (
            .O(N__40855),
            .I(neopxl_color_4));
    Odrv4 I__9037 (
            .O(N__40852),
            .I(neopxl_color_4));
    Odrv4 I__9036 (
            .O(N__40849),
            .I(neopxl_color_4));
    SRMux I__9035 (
            .O(N__40842),
            .I(N__40839));
    LocalMux I__9034 (
            .O(N__40839),
            .I(N__40836));
    Span4Mux_v I__9033 (
            .O(N__40836),
            .I(N__40833));
    Span4Mux_h I__9032 (
            .O(N__40833),
            .I(N__40830));
    Span4Mux_v I__9031 (
            .O(N__40830),
            .I(N__40827));
    Odrv4 I__9030 (
            .O(N__40827),
            .I(n22_adj_732));
    CEMux I__9029 (
            .O(N__40824),
            .I(N__40821));
    LocalMux I__9028 (
            .O(N__40821),
            .I(N__40817));
    CEMux I__9027 (
            .O(N__40820),
            .I(N__40814));
    Span4Mux_v I__9026 (
            .O(N__40817),
            .I(N__40807));
    LocalMux I__9025 (
            .O(N__40814),
            .I(N__40807));
    CEMux I__9024 (
            .O(N__40813),
            .I(N__40803));
    CEMux I__9023 (
            .O(N__40812),
            .I(N__40800));
    Span4Mux_v I__9022 (
            .O(N__40807),
            .I(N__40797));
    InMux I__9021 (
            .O(N__40806),
            .I(N__40794));
    LocalMux I__9020 (
            .O(N__40803),
            .I(N__40789));
    LocalMux I__9019 (
            .O(N__40800),
            .I(N__40789));
    Span4Mux_h I__9018 (
            .O(N__40797),
            .I(N__40784));
    LocalMux I__9017 (
            .O(N__40794),
            .I(N__40784));
    Span4Mux_v I__9016 (
            .O(N__40789),
            .I(N__40779));
    Span4Mux_v I__9015 (
            .O(N__40784),
            .I(N__40779));
    Span4Mux_v I__9014 (
            .O(N__40779),
            .I(N__40776));
    Odrv4 I__9013 (
            .O(N__40776),
            .I(n7232));
    InMux I__9012 (
            .O(N__40773),
            .I(N__40770));
    LocalMux I__9011 (
            .O(N__40770),
            .I(N__40767));
    Odrv4 I__9010 (
            .O(N__40767),
            .I(n43));
    InMux I__9009 (
            .O(N__40764),
            .I(N__40761));
    LocalMux I__9008 (
            .O(N__40761),
            .I(n52_adj_770));
    InMux I__9007 (
            .O(N__40758),
            .I(N__40750));
    InMux I__9006 (
            .O(N__40757),
            .I(N__40750));
    InMux I__9005 (
            .O(N__40756),
            .I(N__40747));
    InMux I__9004 (
            .O(N__40755),
            .I(N__40743));
    LocalMux I__9003 (
            .O(N__40750),
            .I(N__40740));
    LocalMux I__9002 (
            .O(N__40747),
            .I(N__40737));
    InMux I__9001 (
            .O(N__40746),
            .I(N__40734));
    LocalMux I__9000 (
            .O(N__40743),
            .I(N__40729));
    Span12Mux_v I__8999 (
            .O(N__40740),
            .I(N__40729));
    Span12Mux_s10_h I__8998 (
            .O(N__40737),
            .I(N__40726));
    LocalMux I__8997 (
            .O(N__40734),
            .I(neopxl_color_6));
    Odrv12 I__8996 (
            .O(N__40729),
            .I(neopxl_color_6));
    Odrv12 I__8995 (
            .O(N__40726),
            .I(neopxl_color_6));
    SRMux I__8994 (
            .O(N__40719),
            .I(N__40716));
    LocalMux I__8993 (
            .O(N__40716),
            .I(N__40713));
    Odrv12 I__8992 (
            .O(N__40713),
            .I(n22_adj_728));
    CascadeMux I__8991 (
            .O(N__40710),
            .I(n7150_cascade_));
    InMux I__8990 (
            .O(N__40707),
            .I(N__40704));
    LocalMux I__8989 (
            .O(N__40704),
            .I(N__40700));
    InMux I__8988 (
            .O(N__40703),
            .I(N__40697));
    Span4Mux_v I__8987 (
            .O(N__40700),
            .I(N__40694));
    LocalMux I__8986 (
            .O(N__40697),
            .I(N__40691));
    Span4Mux_h I__8985 (
            .O(N__40694),
            .I(N__40688));
    Span4Mux_v I__8984 (
            .O(N__40691),
            .I(N__40685));
    Sp12to4 I__8983 (
            .O(N__40688),
            .I(N__40680));
    Sp12to4 I__8982 (
            .O(N__40685),
            .I(N__40680));
    Span12Mux_s11_h I__8981 (
            .O(N__40680),
            .I(N__40677));
    Span12Mux_v I__8980 (
            .O(N__40677),
            .I(N__40674));
    Odrv12 I__8979 (
            .O(N__40674),
            .I(pin_in_11));
    InMux I__8978 (
            .O(N__40671),
            .I(N__40668));
    LocalMux I__8977 (
            .O(N__40668),
            .I(n2355));
    CascadeMux I__8976 (
            .O(N__40665),
            .I(N__40661));
    InMux I__8975 (
            .O(N__40664),
            .I(N__40658));
    InMux I__8974 (
            .O(N__40661),
            .I(N__40652));
    LocalMux I__8973 (
            .O(N__40658),
            .I(N__40649));
    InMux I__8972 (
            .O(N__40657),
            .I(N__40645));
    InMux I__8971 (
            .O(N__40656),
            .I(N__40642));
    InMux I__8970 (
            .O(N__40655),
            .I(N__40639));
    LocalMux I__8969 (
            .O(N__40652),
            .I(N__40636));
    Span4Mux_h I__8968 (
            .O(N__40649),
            .I(N__40633));
    InMux I__8967 (
            .O(N__40648),
            .I(N__40630));
    LocalMux I__8966 (
            .O(N__40645),
            .I(N__40627));
    LocalMux I__8965 (
            .O(N__40642),
            .I(n21_adj_714));
    LocalMux I__8964 (
            .O(N__40639),
            .I(n21_adj_714));
    Odrv4 I__8963 (
            .O(N__40636),
            .I(n21_adj_714));
    Odrv4 I__8962 (
            .O(N__40633),
            .I(n21_adj_714));
    LocalMux I__8961 (
            .O(N__40630),
            .I(n21_adj_714));
    Odrv12 I__8960 (
            .O(N__40627),
            .I(n21_adj_714));
    CascadeMux I__8959 (
            .O(N__40614),
            .I(n7_adj_719_cascade_));
    InMux I__8958 (
            .O(N__40611),
            .I(N__40606));
    InMux I__8957 (
            .O(N__40610),
            .I(N__40603));
    InMux I__8956 (
            .O(N__40609),
            .I(N__40600));
    LocalMux I__8955 (
            .O(N__40606),
            .I(n7150));
    LocalMux I__8954 (
            .O(N__40603),
            .I(n7150));
    LocalMux I__8953 (
            .O(N__40600),
            .I(n7150));
    CascadeMux I__8952 (
            .O(N__40593),
            .I(N__40590));
    InMux I__8951 (
            .O(N__40590),
            .I(N__40587));
    LocalMux I__8950 (
            .O(N__40587),
            .I(N__40584));
    Sp12to4 I__8949 (
            .O(N__40584),
            .I(N__40580));
    InMux I__8948 (
            .O(N__40583),
            .I(N__40577));
    Span12Mux_v I__8947 (
            .O(N__40580),
            .I(N__40572));
    LocalMux I__8946 (
            .O(N__40577),
            .I(N__40572));
    Span12Mux_h I__8945 (
            .O(N__40572),
            .I(N__40569));
    Span12Mux_v I__8944 (
            .O(N__40569),
            .I(N__40566));
    Odrv12 I__8943 (
            .O(N__40566),
            .I(pin_in_9));
    InMux I__8942 (
            .O(N__40563),
            .I(N__40560));
    LocalMux I__8941 (
            .O(N__40560),
            .I(n2337));
    CascadeMux I__8940 (
            .O(N__40557),
            .I(n2343_cascade_));
    InMux I__8939 (
            .O(N__40554),
            .I(N__40551));
    LocalMux I__8938 (
            .O(N__40551),
            .I(n2325));
    InMux I__8937 (
            .O(N__40548),
            .I(N__40545));
    LocalMux I__8936 (
            .O(N__40545),
            .I(N__40541));
    InMux I__8935 (
            .O(N__40544),
            .I(N__40538));
    Span4Mux_v I__8934 (
            .O(N__40541),
            .I(N__40535));
    LocalMux I__8933 (
            .O(N__40538),
            .I(N__40532));
    Span4Mux_h I__8932 (
            .O(N__40535),
            .I(N__40529));
    Span4Mux_v I__8931 (
            .O(N__40532),
            .I(N__40526));
    Sp12to4 I__8930 (
            .O(N__40529),
            .I(N__40521));
    Sp12to4 I__8929 (
            .O(N__40526),
            .I(N__40521));
    Odrv12 I__8928 (
            .O(N__40521),
            .I(pin_in_3));
    CascadeMux I__8927 (
            .O(N__40518),
            .I(N__40514));
    InMux I__8926 (
            .O(N__40517),
            .I(N__40511));
    InMux I__8925 (
            .O(N__40514),
            .I(N__40508));
    LocalMux I__8924 (
            .O(N__40511),
            .I(N__40505));
    LocalMux I__8923 (
            .O(N__40508),
            .I(N__40502));
    Span4Mux_v I__8922 (
            .O(N__40505),
            .I(N__40499));
    Span12Mux_h I__8921 (
            .O(N__40502),
            .I(N__40494));
    Sp12to4 I__8920 (
            .O(N__40499),
            .I(N__40494));
    Span12Mux_h I__8919 (
            .O(N__40494),
            .I(N__40491));
    Span12Mux_v I__8918 (
            .O(N__40491),
            .I(N__40488));
    Odrv12 I__8917 (
            .O(N__40488),
            .I(pin_in_1));
    InMux I__8916 (
            .O(N__40485),
            .I(N__40482));
    LocalMux I__8915 (
            .O(N__40482),
            .I(n2361));
    InMux I__8914 (
            .O(N__40479),
            .I(N__40475));
    InMux I__8913 (
            .O(N__40478),
            .I(N__40472));
    LocalMux I__8912 (
            .O(N__40475),
            .I(N__40469));
    LocalMux I__8911 (
            .O(N__40472),
            .I(N__40466));
    Span12Mux_v I__8910 (
            .O(N__40469),
            .I(N__40463));
    Span4Mux_v I__8909 (
            .O(N__40466),
            .I(N__40460));
    Span12Mux_h I__8908 (
            .O(N__40463),
            .I(N__40457));
    Sp12to4 I__8907 (
            .O(N__40460),
            .I(N__40454));
    Odrv12 I__8906 (
            .O(N__40457),
            .I(pin_in_2));
    Odrv12 I__8905 (
            .O(N__40454),
            .I(pin_in_2));
    InMux I__8904 (
            .O(N__40449),
            .I(N__40445));
    CascadeMux I__8903 (
            .O(N__40448),
            .I(N__40438));
    LocalMux I__8902 (
            .O(N__40445),
            .I(N__40435));
    InMux I__8901 (
            .O(N__40444),
            .I(N__40432));
    InMux I__8900 (
            .O(N__40443),
            .I(N__40429));
    InMux I__8899 (
            .O(N__40442),
            .I(N__40426));
    InMux I__8898 (
            .O(N__40441),
            .I(N__40423));
    InMux I__8897 (
            .O(N__40438),
            .I(N__40420));
    Span4Mux_v I__8896 (
            .O(N__40435),
            .I(N__40417));
    LocalMux I__8895 (
            .O(N__40432),
            .I(n22_adj_740));
    LocalMux I__8894 (
            .O(N__40429),
            .I(n22_adj_740));
    LocalMux I__8893 (
            .O(N__40426),
            .I(n22_adj_740));
    LocalMux I__8892 (
            .O(N__40423),
            .I(n22_adj_740));
    LocalMux I__8891 (
            .O(N__40420),
            .I(n22_adj_740));
    Odrv4 I__8890 (
            .O(N__40417),
            .I(n22_adj_740));
    CascadeMux I__8889 (
            .O(N__40404),
            .I(n21_adj_741_cascade_));
    InMux I__8888 (
            .O(N__40401),
            .I(N__40398));
    LocalMux I__8887 (
            .O(N__40398),
            .I(N__40394));
    InMux I__8886 (
            .O(N__40397),
            .I(N__40391));
    Span4Mux_v I__8885 (
            .O(N__40394),
            .I(N__40386));
    LocalMux I__8884 (
            .O(N__40391),
            .I(N__40386));
    Odrv4 I__8883 (
            .O(N__40386),
            .I(n7128));
    CascadeMux I__8882 (
            .O(N__40383),
            .I(N__40380));
    InMux I__8881 (
            .O(N__40380),
            .I(N__40377));
    LocalMux I__8880 (
            .O(N__40377),
            .I(N__40373));
    InMux I__8879 (
            .O(N__40376),
            .I(N__40370));
    Odrv4 I__8878 (
            .O(N__40373),
            .I(\nx.n2192 ));
    LocalMux I__8877 (
            .O(N__40370),
            .I(\nx.n2192 ));
    InMux I__8876 (
            .O(N__40365),
            .I(\nx.n10707 ));
    CascadeMux I__8875 (
            .O(N__40362),
            .I(N__40358));
    InMux I__8874 (
            .O(N__40361),
            .I(N__40355));
    InMux I__8873 (
            .O(N__40358),
            .I(N__40348));
    LocalMux I__8872 (
            .O(N__40355),
            .I(N__40343));
    InMux I__8871 (
            .O(N__40354),
            .I(N__40338));
    InMux I__8870 (
            .O(N__40353),
            .I(N__40338));
    InMux I__8869 (
            .O(N__40352),
            .I(N__40335));
    InMux I__8868 (
            .O(N__40351),
            .I(N__40331));
    LocalMux I__8867 (
            .O(N__40348),
            .I(N__40328));
    InMux I__8866 (
            .O(N__40347),
            .I(N__40323));
    InMux I__8865 (
            .O(N__40346),
            .I(N__40323));
    Span4Mux_v I__8864 (
            .O(N__40343),
            .I(N__40320));
    LocalMux I__8863 (
            .O(N__40338),
            .I(N__40317));
    LocalMux I__8862 (
            .O(N__40335),
            .I(N__40314));
    InMux I__8861 (
            .O(N__40334),
            .I(N__40311));
    LocalMux I__8860 (
            .O(N__40331),
            .I(n7155));
    Odrv4 I__8859 (
            .O(N__40328),
            .I(n7155));
    LocalMux I__8858 (
            .O(N__40323),
            .I(n7155));
    Odrv4 I__8857 (
            .O(N__40320),
            .I(n7155));
    Odrv4 I__8856 (
            .O(N__40317),
            .I(n7155));
    Odrv4 I__8855 (
            .O(N__40314),
            .I(n7155));
    LocalMux I__8854 (
            .O(N__40311),
            .I(n7155));
    InMux I__8853 (
            .O(N__40296),
            .I(N__40293));
    LocalMux I__8852 (
            .O(N__40293),
            .I(n6166));
    CascadeMux I__8851 (
            .O(N__40290),
            .I(n6166_cascade_));
    InMux I__8850 (
            .O(N__40287),
            .I(N__40284));
    LocalMux I__8849 (
            .O(N__40284),
            .I(n7286));
    CascadeMux I__8848 (
            .O(N__40281),
            .I(n7_adj_753_cascade_));
    InMux I__8847 (
            .O(N__40278),
            .I(N__40274));
    CascadeMux I__8846 (
            .O(N__40277),
            .I(N__40270));
    LocalMux I__8845 (
            .O(N__40274),
            .I(N__40267));
    InMux I__8844 (
            .O(N__40273),
            .I(N__40264));
    InMux I__8843 (
            .O(N__40270),
            .I(N__40261));
    Span4Mux_v I__8842 (
            .O(N__40267),
            .I(N__40254));
    LocalMux I__8841 (
            .O(N__40264),
            .I(N__40254));
    LocalMux I__8840 (
            .O(N__40261),
            .I(N__40254));
    Odrv4 I__8839 (
            .O(N__40254),
            .I(\nx.n2201 ));
    InMux I__8838 (
            .O(N__40251),
            .I(N__40248));
    LocalMux I__8837 (
            .O(N__40248),
            .I(N__40245));
    Odrv4 I__8836 (
            .O(N__40245),
            .I(\nx.n2268 ));
    InMux I__8835 (
            .O(N__40242),
            .I(\nx.n10698 ));
    InMux I__8834 (
            .O(N__40239),
            .I(\nx.n10699 ));
    InMux I__8833 (
            .O(N__40236),
            .I(\nx.n10700 ));
    InMux I__8832 (
            .O(N__40233),
            .I(\nx.n10701 ));
    CascadeMux I__8831 (
            .O(N__40230),
            .I(N__40225));
    InMux I__8830 (
            .O(N__40229),
            .I(N__40222));
    InMux I__8829 (
            .O(N__40228),
            .I(N__40217));
    InMux I__8828 (
            .O(N__40225),
            .I(N__40217));
    LocalMux I__8827 (
            .O(N__40222),
            .I(N__40214));
    LocalMux I__8826 (
            .O(N__40217),
            .I(N__40211));
    Odrv4 I__8825 (
            .O(N__40214),
            .I(\nx.n2197 ));
    Odrv4 I__8824 (
            .O(N__40211),
            .I(\nx.n2197 ));
    InMux I__8823 (
            .O(N__40206),
            .I(N__40203));
    LocalMux I__8822 (
            .O(N__40203),
            .I(N__40200));
    Span4Mux_v I__8821 (
            .O(N__40200),
            .I(N__40197));
    Odrv4 I__8820 (
            .O(N__40197),
            .I(\nx.n2264 ));
    InMux I__8819 (
            .O(N__40194),
            .I(\nx.n10702 ));
    InMux I__8818 (
            .O(N__40191),
            .I(N__40186));
    InMux I__8817 (
            .O(N__40190),
            .I(N__40183));
    InMux I__8816 (
            .O(N__40189),
            .I(N__40180));
    LocalMux I__8815 (
            .O(N__40186),
            .I(N__40177));
    LocalMux I__8814 (
            .O(N__40183),
            .I(N__40172));
    LocalMux I__8813 (
            .O(N__40180),
            .I(N__40172));
    Odrv4 I__8812 (
            .O(N__40177),
            .I(\nx.n2196 ));
    Odrv4 I__8811 (
            .O(N__40172),
            .I(\nx.n2196 ));
    InMux I__8810 (
            .O(N__40167),
            .I(N__40164));
    LocalMux I__8809 (
            .O(N__40164),
            .I(N__40161));
    Span4Mux_h I__8808 (
            .O(N__40161),
            .I(N__40158));
    Odrv4 I__8807 (
            .O(N__40158),
            .I(\nx.n2263 ));
    InMux I__8806 (
            .O(N__40155),
            .I(\nx.n10703 ));
    CascadeMux I__8805 (
            .O(N__40152),
            .I(N__40148));
    InMux I__8804 (
            .O(N__40151),
            .I(N__40145));
    InMux I__8803 (
            .O(N__40148),
            .I(N__40142));
    LocalMux I__8802 (
            .O(N__40145),
            .I(N__40138));
    LocalMux I__8801 (
            .O(N__40142),
            .I(N__40135));
    InMux I__8800 (
            .O(N__40141),
            .I(N__40132));
    Odrv4 I__8799 (
            .O(N__40138),
            .I(\nx.n2195 ));
    Odrv4 I__8798 (
            .O(N__40135),
            .I(\nx.n2195 ));
    LocalMux I__8797 (
            .O(N__40132),
            .I(\nx.n2195 ));
    CascadeMux I__8796 (
            .O(N__40125),
            .I(N__40122));
    InMux I__8795 (
            .O(N__40122),
            .I(N__40119));
    LocalMux I__8794 (
            .O(N__40119),
            .I(N__40116));
    Span4Mux_h I__8793 (
            .O(N__40116),
            .I(N__40113));
    Odrv4 I__8792 (
            .O(N__40113),
            .I(\nx.n2262 ));
    InMux I__8791 (
            .O(N__40110),
            .I(\nx.n10704 ));
    CascadeMux I__8790 (
            .O(N__40107),
            .I(N__40103));
    CascadeMux I__8789 (
            .O(N__40106),
            .I(N__40100));
    InMux I__8788 (
            .O(N__40103),
            .I(N__40097));
    InMux I__8787 (
            .O(N__40100),
            .I(N__40094));
    LocalMux I__8786 (
            .O(N__40097),
            .I(N__40091));
    LocalMux I__8785 (
            .O(N__40094),
            .I(N__40085));
    Span4Mux_h I__8784 (
            .O(N__40091),
            .I(N__40085));
    InMux I__8783 (
            .O(N__40090),
            .I(N__40082));
    Odrv4 I__8782 (
            .O(N__40085),
            .I(\nx.n2194 ));
    LocalMux I__8781 (
            .O(N__40082),
            .I(\nx.n2194 ));
    InMux I__8780 (
            .O(N__40077),
            .I(N__40074));
    LocalMux I__8779 (
            .O(N__40074),
            .I(N__40071));
    Span4Mux_h I__8778 (
            .O(N__40071),
            .I(N__40068));
    Odrv4 I__8777 (
            .O(N__40068),
            .I(\nx.n2261 ));
    InMux I__8776 (
            .O(N__40065),
            .I(bfn_13_25_0_));
    InMux I__8775 (
            .O(N__40062),
            .I(\nx.n10706 ));
    CascadeMux I__8774 (
            .O(N__40059),
            .I(N__40054));
    InMux I__8773 (
            .O(N__40058),
            .I(N__40051));
    InMux I__8772 (
            .O(N__40057),
            .I(N__40048));
    InMux I__8771 (
            .O(N__40054),
            .I(N__40045));
    LocalMux I__8770 (
            .O(N__40051),
            .I(N__40042));
    LocalMux I__8769 (
            .O(N__40048),
            .I(\nx.n2209 ));
    LocalMux I__8768 (
            .O(N__40045),
            .I(\nx.n2209 ));
    Odrv4 I__8767 (
            .O(N__40042),
            .I(\nx.n2209 ));
    CascadeMux I__8766 (
            .O(N__40035),
            .I(N__40032));
    InMux I__8765 (
            .O(N__40032),
            .I(N__40029));
    LocalMux I__8764 (
            .O(N__40029),
            .I(\nx.n2276 ));
    InMux I__8763 (
            .O(N__40026),
            .I(\nx.n10690 ));
    CascadeMux I__8762 (
            .O(N__40023),
            .I(N__40019));
    InMux I__8761 (
            .O(N__40022),
            .I(N__40015));
    InMux I__8760 (
            .O(N__40019),
            .I(N__40012));
    InMux I__8759 (
            .O(N__40018),
            .I(N__40009));
    LocalMux I__8758 (
            .O(N__40015),
            .I(N__40004));
    LocalMux I__8757 (
            .O(N__40012),
            .I(N__40004));
    LocalMux I__8756 (
            .O(N__40009),
            .I(\nx.n2208 ));
    Odrv4 I__8755 (
            .O(N__40004),
            .I(\nx.n2208 ));
    InMux I__8754 (
            .O(N__39999),
            .I(N__39996));
    LocalMux I__8753 (
            .O(N__39996),
            .I(\nx.n2275 ));
    InMux I__8752 (
            .O(N__39993),
            .I(\nx.n10691 ));
    InMux I__8751 (
            .O(N__39990),
            .I(\nx.n10692 ));
    CascadeMux I__8750 (
            .O(N__39987),
            .I(N__39984));
    InMux I__8749 (
            .O(N__39984),
            .I(N__39979));
    InMux I__8748 (
            .O(N__39983),
            .I(N__39976));
    InMux I__8747 (
            .O(N__39982),
            .I(N__39973));
    LocalMux I__8746 (
            .O(N__39979),
            .I(N__39970));
    LocalMux I__8745 (
            .O(N__39976),
            .I(\nx.n2206 ));
    LocalMux I__8744 (
            .O(N__39973),
            .I(\nx.n2206 ));
    Odrv4 I__8743 (
            .O(N__39970),
            .I(\nx.n2206 ));
    InMux I__8742 (
            .O(N__39963),
            .I(N__39960));
    LocalMux I__8741 (
            .O(N__39960),
            .I(\nx.n2273 ));
    InMux I__8740 (
            .O(N__39957),
            .I(\nx.n10693 ));
    CascadeMux I__8739 (
            .O(N__39954),
            .I(N__39951));
    InMux I__8738 (
            .O(N__39951),
            .I(N__39946));
    InMux I__8737 (
            .O(N__39950),
            .I(N__39941));
    InMux I__8736 (
            .O(N__39949),
            .I(N__39941));
    LocalMux I__8735 (
            .O(N__39946),
            .I(N__39938));
    LocalMux I__8734 (
            .O(N__39941),
            .I(\nx.n2205 ));
    Odrv4 I__8733 (
            .O(N__39938),
            .I(\nx.n2205 ));
    CascadeMux I__8732 (
            .O(N__39933),
            .I(N__39930));
    InMux I__8731 (
            .O(N__39930),
            .I(N__39927));
    LocalMux I__8730 (
            .O(N__39927),
            .I(\nx.n2272 ));
    InMux I__8729 (
            .O(N__39924),
            .I(\nx.n10694 ));
    InMux I__8728 (
            .O(N__39921),
            .I(\nx.n10695 ));
    CascadeMux I__8727 (
            .O(N__39918),
            .I(N__39915));
    InMux I__8726 (
            .O(N__39915),
            .I(N__39912));
    LocalMux I__8725 (
            .O(N__39912),
            .I(N__39907));
    InMux I__8724 (
            .O(N__39911),
            .I(N__39904));
    InMux I__8723 (
            .O(N__39910),
            .I(N__39901));
    Span4Mux_v I__8722 (
            .O(N__39907),
            .I(N__39896));
    LocalMux I__8721 (
            .O(N__39904),
            .I(N__39896));
    LocalMux I__8720 (
            .O(N__39901),
            .I(\nx.n2203 ));
    Odrv4 I__8719 (
            .O(N__39896),
            .I(\nx.n2203 ));
    InMux I__8718 (
            .O(N__39891),
            .I(N__39888));
    LocalMux I__8717 (
            .O(N__39888),
            .I(\nx.n2270 ));
    InMux I__8716 (
            .O(N__39885),
            .I(\nx.n10696 ));
    InMux I__8715 (
            .O(N__39882),
            .I(bfn_13_24_0_));
    CascadeMux I__8714 (
            .O(N__39879),
            .I(\nx.n2300_cascade_ ));
    InMux I__8713 (
            .O(N__39876),
            .I(N__39873));
    LocalMux I__8712 (
            .O(N__39873),
            .I(\nx.n33_adj_644 ));
    InMux I__8711 (
            .O(N__39870),
            .I(N__39867));
    LocalMux I__8710 (
            .O(N__39867),
            .I(\nx.n34_adj_641 ));
    CascadeMux I__8709 (
            .O(N__39864),
            .I(\nx.n32_cascade_ ));
    CascadeMux I__8708 (
            .O(N__39861),
            .I(\nx.n2324_cascade_ ));
    InMux I__8707 (
            .O(N__39858),
            .I(N__39853));
    InMux I__8706 (
            .O(N__39857),
            .I(N__39850));
    InMux I__8705 (
            .O(N__39856),
            .I(N__39847));
    LocalMux I__8704 (
            .O(N__39853),
            .I(N__39843));
    LocalMux I__8703 (
            .O(N__39850),
            .I(N__39838));
    LocalMux I__8702 (
            .O(N__39847),
            .I(N__39838));
    CascadeMux I__8701 (
            .O(N__39846),
            .I(N__39835));
    Span4Mux_v I__8700 (
            .O(N__39843),
            .I(N__39832));
    Span4Mux_v I__8699 (
            .O(N__39838),
            .I(N__39829));
    InMux I__8698 (
            .O(N__39835),
            .I(N__39825));
    Span4Mux_h I__8697 (
            .O(N__39832),
            .I(N__39820));
    Span4Mux_h I__8696 (
            .O(N__39829),
            .I(N__39820));
    InMux I__8695 (
            .O(N__39828),
            .I(N__39817));
    LocalMux I__8694 (
            .O(N__39825),
            .I(N__39814));
    Span4Mux_h I__8693 (
            .O(N__39820),
            .I(N__39811));
    LocalMux I__8692 (
            .O(N__39817),
            .I(\nx.bit_ctr_13 ));
    Odrv4 I__8691 (
            .O(N__39814),
            .I(\nx.bit_ctr_13 ));
    Odrv4 I__8690 (
            .O(N__39811),
            .I(\nx.bit_ctr_13 ));
    InMux I__8689 (
            .O(N__39804),
            .I(N__39801));
    LocalMux I__8688 (
            .O(N__39801),
            .I(\nx.n2277 ));
    InMux I__8687 (
            .O(N__39798),
            .I(bfn_13_23_0_));
    InMux I__8686 (
            .O(N__39795),
            .I(N__39790));
    InMux I__8685 (
            .O(N__39794),
            .I(N__39787));
    InMux I__8684 (
            .O(N__39793),
            .I(N__39784));
    LocalMux I__8683 (
            .O(N__39790),
            .I(N__39779));
    LocalMux I__8682 (
            .O(N__39787),
            .I(N__39779));
    LocalMux I__8681 (
            .O(N__39784),
            .I(N__39774));
    Span4Mux_v I__8680 (
            .O(N__39779),
            .I(N__39771));
    InMux I__8679 (
            .O(N__39778),
            .I(N__39768));
    InMux I__8678 (
            .O(N__39777),
            .I(N__39765));
    Span4Mux_h I__8677 (
            .O(N__39774),
            .I(N__39760));
    Span4Mux_h I__8676 (
            .O(N__39771),
            .I(N__39760));
    LocalMux I__8675 (
            .O(N__39768),
            .I(N__39757));
    LocalMux I__8674 (
            .O(N__39765),
            .I(N__39752));
    Span4Mux_h I__8673 (
            .O(N__39760),
            .I(N__39752));
    Span4Mux_v I__8672 (
            .O(N__39757),
            .I(N__39749));
    Odrv4 I__8671 (
            .O(N__39752),
            .I(neopxl_color_5));
    Odrv4 I__8670 (
            .O(N__39749),
            .I(neopxl_color_5));
    SRMux I__8669 (
            .O(N__39744),
            .I(N__39741));
    LocalMux I__8668 (
            .O(N__39741),
            .I(N__39738));
    Span4Mux_h I__8667 (
            .O(N__39738),
            .I(N__39735));
    Span4Mux_h I__8666 (
            .O(N__39735),
            .I(N__39732));
    Odrv4 I__8665 (
            .O(N__39732),
            .I(n22_adj_730));
    InMux I__8664 (
            .O(N__39729),
            .I(N__39725));
    CascadeMux I__8663 (
            .O(N__39728),
            .I(N__39721));
    LocalMux I__8662 (
            .O(N__39725),
            .I(N__39718));
    InMux I__8661 (
            .O(N__39724),
            .I(N__39715));
    InMux I__8660 (
            .O(N__39721),
            .I(N__39712));
    Odrv4 I__8659 (
            .O(N__39718),
            .I(\nx.n2498 ));
    LocalMux I__8658 (
            .O(N__39715),
            .I(\nx.n2498 ));
    LocalMux I__8657 (
            .O(N__39712),
            .I(\nx.n2498 ));
    CascadeMux I__8656 (
            .O(N__39705),
            .I(\nx.n2404_cascade_ ));
    InMux I__8655 (
            .O(N__39702),
            .I(N__39699));
    LocalMux I__8654 (
            .O(N__39699),
            .I(N__39696));
    Odrv4 I__8653 (
            .O(N__39696),
            .I(\nx.n34_adj_657 ));
    CascadeMux I__8652 (
            .O(N__39693),
            .I(N__39690));
    InMux I__8651 (
            .O(N__39690),
            .I(N__39687));
    LocalMux I__8650 (
            .O(N__39687),
            .I(N__39682));
    InMux I__8649 (
            .O(N__39686),
            .I(N__39679));
    InMux I__8648 (
            .O(N__39685),
            .I(N__39676));
    Span4Mux_v I__8647 (
            .O(N__39682),
            .I(N__39673));
    LocalMux I__8646 (
            .O(N__39679),
            .I(N__39670));
    LocalMux I__8645 (
            .O(N__39676),
            .I(\nx.n2490 ));
    Odrv4 I__8644 (
            .O(N__39673),
            .I(\nx.n2490 ));
    Odrv4 I__8643 (
            .O(N__39670),
            .I(\nx.n2490 ));
    InMux I__8642 (
            .O(N__39663),
            .I(N__39660));
    LocalMux I__8641 (
            .O(N__39660),
            .I(N__39656));
    CascadeMux I__8640 (
            .O(N__39659),
            .I(N__39653));
    Span4Mux_h I__8639 (
            .O(N__39656),
            .I(N__39650));
    InMux I__8638 (
            .O(N__39653),
            .I(N__39647));
    Odrv4 I__8637 (
            .O(N__39650),
            .I(\nx.n2504 ));
    LocalMux I__8636 (
            .O(N__39647),
            .I(\nx.n2504 ));
    CascadeMux I__8635 (
            .O(N__39642),
            .I(\nx.n22_adj_637_cascade_ ));
    InMux I__8634 (
            .O(N__39639),
            .I(N__39634));
    CascadeMux I__8633 (
            .O(N__39638),
            .I(N__39631));
    InMux I__8632 (
            .O(N__39637),
            .I(N__39628));
    LocalMux I__8631 (
            .O(N__39634),
            .I(N__39625));
    InMux I__8630 (
            .O(N__39631),
            .I(N__39622));
    LocalMux I__8629 (
            .O(N__39628),
            .I(N__39619));
    Span4Mux_v I__8628 (
            .O(N__39625),
            .I(N__39616));
    LocalMux I__8627 (
            .O(N__39622),
            .I(N__39613));
    Odrv4 I__8626 (
            .O(N__39619),
            .I(\nx.n2507 ));
    Odrv4 I__8625 (
            .O(N__39616),
            .I(\nx.n2507 ));
    Odrv4 I__8624 (
            .O(N__39613),
            .I(\nx.n2507 ));
    InMux I__8623 (
            .O(N__39606),
            .I(N__39603));
    LocalMux I__8622 (
            .O(N__39603),
            .I(N__39600));
    Odrv4 I__8621 (
            .O(N__39600),
            .I(\nx.n37_adj_638 ));
    InMux I__8620 (
            .O(N__39597),
            .I(N__39594));
    LocalMux I__8619 (
            .O(N__39594),
            .I(N__39590));
    CascadeMux I__8618 (
            .O(N__39593),
            .I(N__39587));
    Span4Mux_h I__8617 (
            .O(N__39590),
            .I(N__39583));
    InMux I__8616 (
            .O(N__39587),
            .I(N__39580));
    InMux I__8615 (
            .O(N__39586),
            .I(N__39577));
    Odrv4 I__8614 (
            .O(N__39583),
            .I(\nx.n2500 ));
    LocalMux I__8613 (
            .O(N__39580),
            .I(\nx.n2500 ));
    LocalMux I__8612 (
            .O(N__39577),
            .I(\nx.n2500 ));
    InMux I__8611 (
            .O(N__39570),
            .I(N__39567));
    LocalMux I__8610 (
            .O(N__39567),
            .I(N__39564));
    Odrv4 I__8609 (
            .O(N__39564),
            .I(n13483));
    InMux I__8608 (
            .O(N__39561),
            .I(N__39558));
    LocalMux I__8607 (
            .O(N__39558),
            .I(n13360));
    InMux I__8606 (
            .O(N__39555),
            .I(N__39552));
    LocalMux I__8605 (
            .O(N__39552),
            .I(\nx.n2575 ));
    CascadeMux I__8604 (
            .O(N__39549),
            .I(N__39545));
    CascadeMux I__8603 (
            .O(N__39548),
            .I(N__39541));
    InMux I__8602 (
            .O(N__39545),
            .I(N__39533));
    InMux I__8601 (
            .O(N__39544),
            .I(N__39530));
    InMux I__8600 (
            .O(N__39541),
            .I(N__39527));
    CascadeMux I__8599 (
            .O(N__39540),
            .I(N__39520));
    CascadeMux I__8598 (
            .O(N__39539),
            .I(N__39514));
    CascadeMux I__8597 (
            .O(N__39538),
            .I(N__39510));
    CascadeMux I__8596 (
            .O(N__39537),
            .I(N__39504));
    CascadeMux I__8595 (
            .O(N__39536),
            .I(N__39500));
    LocalMux I__8594 (
            .O(N__39533),
            .I(N__39496));
    LocalMux I__8593 (
            .O(N__39530),
            .I(N__39491));
    LocalMux I__8592 (
            .O(N__39527),
            .I(N__39491));
    InMux I__8591 (
            .O(N__39526),
            .I(N__39488));
    InMux I__8590 (
            .O(N__39525),
            .I(N__39483));
    InMux I__8589 (
            .O(N__39524),
            .I(N__39483));
    InMux I__8588 (
            .O(N__39523),
            .I(N__39474));
    InMux I__8587 (
            .O(N__39520),
            .I(N__39474));
    InMux I__8586 (
            .O(N__39519),
            .I(N__39474));
    InMux I__8585 (
            .O(N__39518),
            .I(N__39474));
    InMux I__8584 (
            .O(N__39517),
            .I(N__39463));
    InMux I__8583 (
            .O(N__39514),
            .I(N__39463));
    InMux I__8582 (
            .O(N__39513),
            .I(N__39463));
    InMux I__8581 (
            .O(N__39510),
            .I(N__39463));
    InMux I__8580 (
            .O(N__39509),
            .I(N__39463));
    InMux I__8579 (
            .O(N__39508),
            .I(N__39460));
    InMux I__8578 (
            .O(N__39507),
            .I(N__39457));
    InMux I__8577 (
            .O(N__39504),
            .I(N__39448));
    InMux I__8576 (
            .O(N__39503),
            .I(N__39448));
    InMux I__8575 (
            .O(N__39500),
            .I(N__39448));
    InMux I__8574 (
            .O(N__39499),
            .I(N__39448));
    Span4Mux_v I__8573 (
            .O(N__39496),
            .I(N__39443));
    Span4Mux_v I__8572 (
            .O(N__39491),
            .I(N__39443));
    LocalMux I__8571 (
            .O(N__39488),
            .I(N__39440));
    LocalMux I__8570 (
            .O(N__39483),
            .I(\nx.n2522 ));
    LocalMux I__8569 (
            .O(N__39474),
            .I(\nx.n2522 ));
    LocalMux I__8568 (
            .O(N__39463),
            .I(\nx.n2522 ));
    LocalMux I__8567 (
            .O(N__39460),
            .I(\nx.n2522 ));
    LocalMux I__8566 (
            .O(N__39457),
            .I(\nx.n2522 ));
    LocalMux I__8565 (
            .O(N__39448),
            .I(\nx.n2522 ));
    Odrv4 I__8564 (
            .O(N__39443),
            .I(\nx.n2522 ));
    Odrv4 I__8563 (
            .O(N__39440),
            .I(\nx.n2522 ));
    InMux I__8562 (
            .O(N__39423),
            .I(N__39419));
    CascadeMux I__8561 (
            .O(N__39422),
            .I(N__39416));
    LocalMux I__8560 (
            .O(N__39419),
            .I(N__39413));
    InMux I__8559 (
            .O(N__39416),
            .I(N__39409));
    Span4Mux_v I__8558 (
            .O(N__39413),
            .I(N__39406));
    InMux I__8557 (
            .O(N__39412),
            .I(N__39403));
    LocalMux I__8556 (
            .O(N__39409),
            .I(N__39400));
    Span4Mux_h I__8555 (
            .O(N__39406),
            .I(N__39395));
    LocalMux I__8554 (
            .O(N__39403),
            .I(N__39395));
    Span4Mux_h I__8553 (
            .O(N__39400),
            .I(N__39392));
    Odrv4 I__8552 (
            .O(N__39395),
            .I(\nx.n2607 ));
    Odrv4 I__8551 (
            .O(N__39392),
            .I(\nx.n2607 ));
    CascadeMux I__8550 (
            .O(N__39387),
            .I(N__39384));
    InMux I__8549 (
            .O(N__39384),
            .I(N__39381));
    LocalMux I__8548 (
            .O(N__39381),
            .I(N__39377));
    CascadeMux I__8547 (
            .O(N__39380),
            .I(N__39373));
    Span4Mux_v I__8546 (
            .O(N__39377),
            .I(N__39370));
    InMux I__8545 (
            .O(N__39376),
            .I(N__39367));
    InMux I__8544 (
            .O(N__39373),
            .I(N__39364));
    Odrv4 I__8543 (
            .O(N__39370),
            .I(\nx.n2495 ));
    LocalMux I__8542 (
            .O(N__39367),
            .I(\nx.n2495 ));
    LocalMux I__8541 (
            .O(N__39364),
            .I(\nx.n2495 ));
    CascadeMux I__8540 (
            .O(N__39357),
            .I(N__39354));
    InMux I__8539 (
            .O(N__39354),
            .I(N__39351));
    LocalMux I__8538 (
            .O(N__39351),
            .I(N__39347));
    CascadeMux I__8537 (
            .O(N__39350),
            .I(N__39344));
    Span4Mux_v I__8536 (
            .O(N__39347),
            .I(N__39341));
    InMux I__8535 (
            .O(N__39344),
            .I(N__39338));
    Odrv4 I__8534 (
            .O(N__39341),
            .I(\nx.n2503 ));
    LocalMux I__8533 (
            .O(N__39338),
            .I(\nx.n2503 ));
    CascadeMux I__8532 (
            .O(N__39333),
            .I(\nx.n2503_cascade_ ));
    InMux I__8531 (
            .O(N__39330),
            .I(N__39327));
    LocalMux I__8530 (
            .O(N__39327),
            .I(\nx.n36_adj_636 ));
    CascadeMux I__8529 (
            .O(N__39324),
            .I(N__39321));
    InMux I__8528 (
            .O(N__39321),
            .I(N__39317));
    CascadeMux I__8527 (
            .O(N__39320),
            .I(N__39313));
    LocalMux I__8526 (
            .O(N__39317),
            .I(N__39310));
    InMux I__8525 (
            .O(N__39316),
            .I(N__39307));
    InMux I__8524 (
            .O(N__39313),
            .I(N__39304));
    Odrv4 I__8523 (
            .O(N__39310),
            .I(\nx.n2502 ));
    LocalMux I__8522 (
            .O(N__39307),
            .I(\nx.n2502 ));
    LocalMux I__8521 (
            .O(N__39304),
            .I(\nx.n2502 ));
    CascadeMux I__8520 (
            .O(N__39297),
            .I(N__39293));
    CascadeMux I__8519 (
            .O(N__39296),
            .I(N__39289));
    InMux I__8518 (
            .O(N__39293),
            .I(N__39286));
    InMux I__8517 (
            .O(N__39292),
            .I(N__39283));
    InMux I__8516 (
            .O(N__39289),
            .I(N__39280));
    LocalMux I__8515 (
            .O(N__39286),
            .I(\nx.n2508 ));
    LocalMux I__8514 (
            .O(N__39283),
            .I(\nx.n2508 ));
    LocalMux I__8513 (
            .O(N__39280),
            .I(\nx.n2508 ));
    CascadeMux I__8512 (
            .O(N__39273),
            .I(N__39269));
    CascadeMux I__8511 (
            .O(N__39272),
            .I(N__39265));
    InMux I__8510 (
            .O(N__39269),
            .I(N__39262));
    InMux I__8509 (
            .O(N__39268),
            .I(N__39259));
    InMux I__8508 (
            .O(N__39265),
            .I(N__39256));
    LocalMux I__8507 (
            .O(N__39262),
            .I(\nx.n2506 ));
    LocalMux I__8506 (
            .O(N__39259),
            .I(\nx.n2506 ));
    LocalMux I__8505 (
            .O(N__39256),
            .I(\nx.n2506 ));
    InMux I__8504 (
            .O(N__39249),
            .I(N__39243));
    InMux I__8503 (
            .O(N__39248),
            .I(N__39243));
    LocalMux I__8502 (
            .O(N__39243),
            .I(N__39240));
    Span12Mux_h I__8501 (
            .O(N__39240),
            .I(N__39237));
    Span12Mux_v I__8500 (
            .O(N__39237),
            .I(N__39234));
    Odrv12 I__8499 (
            .O(N__39234),
            .I(pin_in_8));
    CascadeMux I__8498 (
            .O(N__39231),
            .I(n13480_cascade_));
    CascadeMux I__8497 (
            .O(N__39228),
            .I(current_pin_7__N_157_cascade_));
    InMux I__8496 (
            .O(N__39225),
            .I(N__39222));
    LocalMux I__8495 (
            .O(N__39222),
            .I(N__39218));
    InMux I__8494 (
            .O(N__39221),
            .I(N__39215));
    Span4Mux_v I__8493 (
            .O(N__39218),
            .I(N__39212));
    LocalMux I__8492 (
            .O(N__39215),
            .I(N__39209));
    Span4Mux_h I__8491 (
            .O(N__39212),
            .I(N__39204));
    Span4Mux_v I__8490 (
            .O(N__39209),
            .I(N__39204));
    Span4Mux_h I__8489 (
            .O(N__39204),
            .I(N__39201));
    Sp12to4 I__8488 (
            .O(N__39201),
            .I(N__39198));
    Odrv12 I__8487 (
            .O(N__39198),
            .I(pin_in_0));
    InMux I__8486 (
            .O(N__39195),
            .I(N__39191));
    CascadeMux I__8485 (
            .O(N__39194),
            .I(N__39188));
    LocalMux I__8484 (
            .O(N__39191),
            .I(N__39185));
    InMux I__8483 (
            .O(N__39188),
            .I(N__39182));
    Span4Mux_v I__8482 (
            .O(N__39185),
            .I(N__39179));
    LocalMux I__8481 (
            .O(N__39182),
            .I(N__39176));
    Span4Mux_v I__8480 (
            .O(N__39179),
            .I(N__39173));
    Span4Mux_h I__8479 (
            .O(N__39176),
            .I(N__39170));
    Span4Mux_v I__8478 (
            .O(N__39173),
            .I(N__39167));
    Sp12to4 I__8477 (
            .O(N__39170),
            .I(N__39164));
    Sp12to4 I__8476 (
            .O(N__39167),
            .I(N__39159));
    Span12Mux_v I__8475 (
            .O(N__39164),
            .I(N__39159));
    Span12Mux_h I__8474 (
            .O(N__39159),
            .I(N__39156));
    Odrv12 I__8473 (
            .O(N__39156),
            .I(pin_in_10));
    CascadeMux I__8472 (
            .O(N__39153),
            .I(n2289_cascade_));
    CascadeMux I__8471 (
            .O(N__39150),
            .I(N__39146));
    InMux I__8470 (
            .O(N__39149),
            .I(N__39143));
    InMux I__8469 (
            .O(N__39146),
            .I(N__39140));
    LocalMux I__8468 (
            .O(N__39143),
            .I(N__39137));
    LocalMux I__8467 (
            .O(N__39140),
            .I(N__39134));
    Span4Mux_v I__8466 (
            .O(N__39137),
            .I(N__39131));
    Span4Mux_h I__8465 (
            .O(N__39134),
            .I(N__39128));
    Span4Mux_v I__8464 (
            .O(N__39131),
            .I(N__39125));
    Sp12to4 I__8463 (
            .O(N__39128),
            .I(N__39122));
    Span4Mux_v I__8462 (
            .O(N__39125),
            .I(N__39119));
    Span12Mux_v I__8461 (
            .O(N__39122),
            .I(N__39116));
    Span4Mux_h I__8460 (
            .O(N__39119),
            .I(N__39113));
    Odrv12 I__8459 (
            .O(N__39116),
            .I(pin_in_6));
    Odrv4 I__8458 (
            .O(N__39113),
            .I(pin_in_6));
    InMux I__8457 (
            .O(N__39108),
            .I(N__39105));
    LocalMux I__8456 (
            .O(N__39105),
            .I(N__39102));
    Span4Mux_h I__8455 (
            .O(N__39102),
            .I(N__39099));
    Odrv4 I__8454 (
            .O(N__39099),
            .I(n13453));
    CascadeMux I__8453 (
            .O(N__39096),
            .I(n13364_cascade_));
    InMux I__8452 (
            .O(N__39093),
            .I(N__39090));
    LocalMux I__8451 (
            .O(N__39090),
            .I(n150));
    CascadeMux I__8450 (
            .O(N__39087),
            .I(n7155_cascade_));
    InMux I__8449 (
            .O(N__39084),
            .I(N__39081));
    LocalMux I__8448 (
            .O(N__39081),
            .I(N__39078));
    Odrv4 I__8447 (
            .O(N__39078),
            .I(n6190));
    CascadeMux I__8446 (
            .O(N__39075),
            .I(n6190_cascade_));
    InMux I__8445 (
            .O(N__39072),
            .I(N__39069));
    LocalMux I__8444 (
            .O(N__39069),
            .I(N__39066));
    Odrv4 I__8443 (
            .O(N__39066),
            .I(n7334));
    InMux I__8442 (
            .O(N__39063),
            .I(N__39057));
    InMux I__8441 (
            .O(N__39062),
            .I(N__39057));
    LocalMux I__8440 (
            .O(N__39057),
            .I(n6170));
    InMux I__8439 (
            .O(N__39054),
            .I(N__39050));
    InMux I__8438 (
            .O(N__39053),
            .I(N__39047));
    LocalMux I__8437 (
            .O(N__39050),
            .I(n9415));
    LocalMux I__8436 (
            .O(N__39047),
            .I(n9415));
    InMux I__8435 (
            .O(N__39042),
            .I(N__39038));
    InMux I__8434 (
            .O(N__39041),
            .I(N__39035));
    LocalMux I__8433 (
            .O(N__39038),
            .I(delay_counter_28));
    LocalMux I__8432 (
            .O(N__39035),
            .I(delay_counter_28));
    InMux I__8431 (
            .O(N__39030),
            .I(n10544));
    InMux I__8430 (
            .O(N__39027),
            .I(N__39023));
    InMux I__8429 (
            .O(N__39026),
            .I(N__39020));
    LocalMux I__8428 (
            .O(N__39023),
            .I(delay_counter_29));
    LocalMux I__8427 (
            .O(N__39020),
            .I(delay_counter_29));
    InMux I__8426 (
            .O(N__39015),
            .I(n10545));
    InMux I__8425 (
            .O(N__39012),
            .I(N__39008));
    InMux I__8424 (
            .O(N__39011),
            .I(N__39005));
    LocalMux I__8423 (
            .O(N__39008),
            .I(delay_counter_30));
    LocalMux I__8422 (
            .O(N__39005),
            .I(delay_counter_30));
    InMux I__8421 (
            .O(N__39000),
            .I(n10546));
    InMux I__8420 (
            .O(N__38997),
            .I(n10547));
    SRMux I__8419 (
            .O(N__38994),
            .I(N__38990));
    SRMux I__8418 (
            .O(N__38993),
            .I(N__38986));
    LocalMux I__8417 (
            .O(N__38990),
            .I(N__38983));
    SRMux I__8416 (
            .O(N__38989),
            .I(N__38980));
    LocalMux I__8415 (
            .O(N__38986),
            .I(N__38977));
    Span4Mux_v I__8414 (
            .O(N__38983),
            .I(N__38973));
    LocalMux I__8413 (
            .O(N__38980),
            .I(N__38970));
    Span4Mux_h I__8412 (
            .O(N__38977),
            .I(N__38967));
    SRMux I__8411 (
            .O(N__38976),
            .I(N__38964));
    Odrv4 I__8410 (
            .O(N__38973),
            .I(n7442));
    Odrv12 I__8409 (
            .O(N__38970),
            .I(n7442));
    Odrv4 I__8408 (
            .O(N__38967),
            .I(n7442));
    LocalMux I__8407 (
            .O(N__38964),
            .I(n7442));
    CascadeMux I__8406 (
            .O(N__38955),
            .I(n10_adj_779_cascade_));
    InMux I__8405 (
            .O(N__38952),
            .I(N__38949));
    LocalMux I__8404 (
            .O(N__38949),
            .I(n10_adj_779));
    CascadeMux I__8403 (
            .O(N__38946),
            .I(n7290_cascade_));
    IoInMux I__8402 (
            .O(N__38943),
            .I(N__38940));
    LocalMux I__8401 (
            .O(N__38940),
            .I(N__38937));
    Span4Mux_s3_v I__8400 (
            .O(N__38937),
            .I(N__38934));
    Span4Mux_h I__8399 (
            .O(N__38934),
            .I(N__38931));
    Sp12to4 I__8398 (
            .O(N__38931),
            .I(N__38928));
    Span12Mux_v I__8397 (
            .O(N__38928),
            .I(N__38923));
    InMux I__8396 (
            .O(N__38927),
            .I(N__38920));
    InMux I__8395 (
            .O(N__38926),
            .I(N__38917));
    Odrv12 I__8394 (
            .O(N__38923),
            .I(pin_out_10));
    LocalMux I__8393 (
            .O(N__38920),
            .I(pin_out_10));
    LocalMux I__8392 (
            .O(N__38917),
            .I(pin_out_10));
    InMux I__8391 (
            .O(N__38910),
            .I(N__38907));
    LocalMux I__8390 (
            .O(N__38907),
            .I(N__38903));
    InMux I__8389 (
            .O(N__38906),
            .I(N__38900));
    Span4Mux_h I__8388 (
            .O(N__38903),
            .I(N__38897));
    LocalMux I__8387 (
            .O(N__38900),
            .I(N__38894));
    Odrv4 I__8386 (
            .O(N__38897),
            .I(n7135));
    Odrv4 I__8385 (
            .O(N__38894),
            .I(n7135));
    InMux I__8384 (
            .O(N__38889),
            .I(N__38885));
    InMux I__8383 (
            .O(N__38888),
            .I(N__38882));
    LocalMux I__8382 (
            .O(N__38885),
            .I(N__38879));
    LocalMux I__8381 (
            .O(N__38882),
            .I(delay_counter_20));
    Odrv4 I__8380 (
            .O(N__38879),
            .I(delay_counter_20));
    InMux I__8379 (
            .O(N__38874),
            .I(n10536));
    InMux I__8378 (
            .O(N__38871),
            .I(N__38867));
    InMux I__8377 (
            .O(N__38870),
            .I(N__38864));
    LocalMux I__8376 (
            .O(N__38867),
            .I(delay_counter_21));
    LocalMux I__8375 (
            .O(N__38864),
            .I(delay_counter_21));
    InMux I__8374 (
            .O(N__38859),
            .I(n10537));
    CascadeMux I__8373 (
            .O(N__38856),
            .I(N__38852));
    InMux I__8372 (
            .O(N__38855),
            .I(N__38849));
    InMux I__8371 (
            .O(N__38852),
            .I(N__38846));
    LocalMux I__8370 (
            .O(N__38849),
            .I(delay_counter_22));
    LocalMux I__8369 (
            .O(N__38846),
            .I(delay_counter_22));
    InMux I__8368 (
            .O(N__38841),
            .I(n10538));
    InMux I__8367 (
            .O(N__38838),
            .I(N__38834));
    InMux I__8366 (
            .O(N__38837),
            .I(N__38831));
    LocalMux I__8365 (
            .O(N__38834),
            .I(delay_counter_23));
    LocalMux I__8364 (
            .O(N__38831),
            .I(delay_counter_23));
    InMux I__8363 (
            .O(N__38826),
            .I(n10539));
    InMux I__8362 (
            .O(N__38823),
            .I(N__38819));
    InMux I__8361 (
            .O(N__38822),
            .I(N__38816));
    LocalMux I__8360 (
            .O(N__38819),
            .I(delay_counter_24));
    LocalMux I__8359 (
            .O(N__38816),
            .I(delay_counter_24));
    InMux I__8358 (
            .O(N__38811),
            .I(bfn_12_29_0_));
    InMux I__8357 (
            .O(N__38808),
            .I(N__38804));
    InMux I__8356 (
            .O(N__38807),
            .I(N__38801));
    LocalMux I__8355 (
            .O(N__38804),
            .I(delay_counter_25));
    LocalMux I__8354 (
            .O(N__38801),
            .I(delay_counter_25));
    InMux I__8353 (
            .O(N__38796),
            .I(n10541));
    InMux I__8352 (
            .O(N__38793),
            .I(N__38789));
    InMux I__8351 (
            .O(N__38792),
            .I(N__38786));
    LocalMux I__8350 (
            .O(N__38789),
            .I(delay_counter_26));
    LocalMux I__8349 (
            .O(N__38786),
            .I(delay_counter_26));
    InMux I__8348 (
            .O(N__38781),
            .I(n10542));
    CascadeMux I__8347 (
            .O(N__38778),
            .I(N__38774));
    InMux I__8346 (
            .O(N__38777),
            .I(N__38771));
    InMux I__8345 (
            .O(N__38774),
            .I(N__38768));
    LocalMux I__8344 (
            .O(N__38771),
            .I(delay_counter_27));
    LocalMux I__8343 (
            .O(N__38768),
            .I(delay_counter_27));
    InMux I__8342 (
            .O(N__38763),
            .I(n10543));
    InMux I__8341 (
            .O(N__38760),
            .I(N__38756));
    InMux I__8340 (
            .O(N__38759),
            .I(N__38753));
    LocalMux I__8339 (
            .O(N__38756),
            .I(delay_counter_12));
    LocalMux I__8338 (
            .O(N__38753),
            .I(delay_counter_12));
    InMux I__8337 (
            .O(N__38748),
            .I(n10528));
    InMux I__8336 (
            .O(N__38745),
            .I(N__38741));
    InMux I__8335 (
            .O(N__38744),
            .I(N__38738));
    LocalMux I__8334 (
            .O(N__38741),
            .I(delay_counter_13));
    LocalMux I__8333 (
            .O(N__38738),
            .I(delay_counter_13));
    InMux I__8332 (
            .O(N__38733),
            .I(n10529));
    InMux I__8331 (
            .O(N__38730),
            .I(N__38726));
    InMux I__8330 (
            .O(N__38729),
            .I(N__38723));
    LocalMux I__8329 (
            .O(N__38726),
            .I(delay_counter_14));
    LocalMux I__8328 (
            .O(N__38723),
            .I(delay_counter_14));
    InMux I__8327 (
            .O(N__38718),
            .I(n10530));
    CascadeMux I__8326 (
            .O(N__38715),
            .I(N__38712));
    InMux I__8325 (
            .O(N__38712),
            .I(N__38709));
    LocalMux I__8324 (
            .O(N__38709),
            .I(N__38705));
    InMux I__8323 (
            .O(N__38708),
            .I(N__38702));
    Span4Mux_h I__8322 (
            .O(N__38705),
            .I(N__38699));
    LocalMux I__8321 (
            .O(N__38702),
            .I(delay_counter_15));
    Odrv4 I__8320 (
            .O(N__38699),
            .I(delay_counter_15));
    InMux I__8319 (
            .O(N__38694),
            .I(n10531));
    InMux I__8318 (
            .O(N__38691),
            .I(N__38687));
    InMux I__8317 (
            .O(N__38690),
            .I(N__38684));
    LocalMux I__8316 (
            .O(N__38687),
            .I(N__38681));
    LocalMux I__8315 (
            .O(N__38684),
            .I(delay_counter_16));
    Odrv4 I__8314 (
            .O(N__38681),
            .I(delay_counter_16));
    InMux I__8313 (
            .O(N__38676),
            .I(bfn_12_28_0_));
    InMux I__8312 (
            .O(N__38673),
            .I(N__38670));
    LocalMux I__8311 (
            .O(N__38670),
            .I(N__38666));
    InMux I__8310 (
            .O(N__38669),
            .I(N__38663));
    Span4Mux_h I__8309 (
            .O(N__38666),
            .I(N__38660));
    LocalMux I__8308 (
            .O(N__38663),
            .I(delay_counter_17));
    Odrv4 I__8307 (
            .O(N__38660),
            .I(delay_counter_17));
    InMux I__8306 (
            .O(N__38655),
            .I(n10533));
    InMux I__8305 (
            .O(N__38652),
            .I(N__38649));
    LocalMux I__8304 (
            .O(N__38649),
            .I(N__38645));
    InMux I__8303 (
            .O(N__38648),
            .I(N__38642));
    Span4Mux_h I__8302 (
            .O(N__38645),
            .I(N__38639));
    LocalMux I__8301 (
            .O(N__38642),
            .I(delay_counter_18));
    Odrv4 I__8300 (
            .O(N__38639),
            .I(delay_counter_18));
    InMux I__8299 (
            .O(N__38634),
            .I(n10534));
    InMux I__8298 (
            .O(N__38631),
            .I(N__38627));
    InMux I__8297 (
            .O(N__38630),
            .I(N__38624));
    LocalMux I__8296 (
            .O(N__38627),
            .I(N__38621));
    LocalMux I__8295 (
            .O(N__38624),
            .I(delay_counter_19));
    Odrv4 I__8294 (
            .O(N__38621),
            .I(delay_counter_19));
    InMux I__8293 (
            .O(N__38616),
            .I(n10535));
    InMux I__8292 (
            .O(N__38613),
            .I(N__38609));
    InMux I__8291 (
            .O(N__38612),
            .I(N__38606));
    LocalMux I__8290 (
            .O(N__38609),
            .I(delay_counter_3));
    LocalMux I__8289 (
            .O(N__38606),
            .I(delay_counter_3));
    InMux I__8288 (
            .O(N__38601),
            .I(n10519));
    InMux I__8287 (
            .O(N__38598),
            .I(N__38594));
    InMux I__8286 (
            .O(N__38597),
            .I(N__38591));
    LocalMux I__8285 (
            .O(N__38594),
            .I(delay_counter_4));
    LocalMux I__8284 (
            .O(N__38591),
            .I(delay_counter_4));
    InMux I__8283 (
            .O(N__38586),
            .I(n10520));
    InMux I__8282 (
            .O(N__38583),
            .I(N__38579));
    InMux I__8281 (
            .O(N__38582),
            .I(N__38576));
    LocalMux I__8280 (
            .O(N__38579),
            .I(delay_counter_5));
    LocalMux I__8279 (
            .O(N__38576),
            .I(delay_counter_5));
    InMux I__8278 (
            .O(N__38571),
            .I(n10521));
    InMux I__8277 (
            .O(N__38568),
            .I(N__38564));
    InMux I__8276 (
            .O(N__38567),
            .I(N__38561));
    LocalMux I__8275 (
            .O(N__38564),
            .I(delay_counter_6));
    LocalMux I__8274 (
            .O(N__38561),
            .I(delay_counter_6));
    InMux I__8273 (
            .O(N__38556),
            .I(n10522));
    InMux I__8272 (
            .O(N__38553),
            .I(N__38549));
    InMux I__8271 (
            .O(N__38552),
            .I(N__38546));
    LocalMux I__8270 (
            .O(N__38549),
            .I(delay_counter_7));
    LocalMux I__8269 (
            .O(N__38546),
            .I(delay_counter_7));
    InMux I__8268 (
            .O(N__38541),
            .I(n10523));
    InMux I__8267 (
            .O(N__38538),
            .I(N__38534));
    InMux I__8266 (
            .O(N__38537),
            .I(N__38531));
    LocalMux I__8265 (
            .O(N__38534),
            .I(delay_counter_8));
    LocalMux I__8264 (
            .O(N__38531),
            .I(delay_counter_8));
    InMux I__8263 (
            .O(N__38526),
            .I(bfn_12_27_0_));
    CascadeMux I__8262 (
            .O(N__38523),
            .I(N__38519));
    InMux I__8261 (
            .O(N__38522),
            .I(N__38516));
    InMux I__8260 (
            .O(N__38519),
            .I(N__38513));
    LocalMux I__8259 (
            .O(N__38516),
            .I(delay_counter_9));
    LocalMux I__8258 (
            .O(N__38513),
            .I(delay_counter_9));
    InMux I__8257 (
            .O(N__38508),
            .I(n10525));
    InMux I__8256 (
            .O(N__38505),
            .I(N__38501));
    InMux I__8255 (
            .O(N__38504),
            .I(N__38498));
    LocalMux I__8254 (
            .O(N__38501),
            .I(delay_counter_10));
    LocalMux I__8253 (
            .O(N__38498),
            .I(delay_counter_10));
    InMux I__8252 (
            .O(N__38493),
            .I(n10526));
    InMux I__8251 (
            .O(N__38490),
            .I(N__38486));
    InMux I__8250 (
            .O(N__38489),
            .I(N__38483));
    LocalMux I__8249 (
            .O(N__38486),
            .I(delay_counter_11));
    LocalMux I__8248 (
            .O(N__38483),
            .I(delay_counter_11));
    InMux I__8247 (
            .O(N__38478),
            .I(n10527));
    CascadeMux I__8246 (
            .O(N__38475),
            .I(N__38472));
    InMux I__8245 (
            .O(N__38472),
            .I(N__38469));
    LocalMux I__8244 (
            .O(N__38469),
            .I(\nx.n31 ));
    InMux I__8243 (
            .O(N__38466),
            .I(N__38463));
    LocalMux I__8242 (
            .O(N__38463),
            .I(\nx.n28_adj_601 ));
    InMux I__8241 (
            .O(N__38460),
            .I(N__38457));
    LocalMux I__8240 (
            .O(N__38457),
            .I(N__38454));
    Sp12to4 I__8239 (
            .O(N__38454),
            .I(N__38450));
    InMux I__8238 (
            .O(N__38453),
            .I(N__38447));
    Span12Mux_s10_v I__8237 (
            .O(N__38450),
            .I(N__38442));
    LocalMux I__8236 (
            .O(N__38447),
            .I(N__38439));
    InMux I__8235 (
            .O(N__38446),
            .I(N__38434));
    InMux I__8234 (
            .O(N__38445),
            .I(N__38434));
    Odrv12 I__8233 (
            .O(N__38442),
            .I(neopxl_color_12));
    Odrv4 I__8232 (
            .O(N__38439),
            .I(neopxl_color_12));
    LocalMux I__8231 (
            .O(N__38434),
            .I(neopxl_color_12));
    InMux I__8230 (
            .O(N__38427),
            .I(N__38424));
    LocalMux I__8229 (
            .O(N__38424),
            .I(N__38421));
    Span4Mux_h I__8228 (
            .O(N__38421),
            .I(N__38418));
    Span4Mux_h I__8227 (
            .O(N__38418),
            .I(N__38415));
    Span4Mux_h I__8226 (
            .O(N__38415),
            .I(N__38412));
    Odrv4 I__8225 (
            .O(N__38412),
            .I(neopxl_color_prev_12));
    InMux I__8224 (
            .O(N__38409),
            .I(N__38406));
    LocalMux I__8223 (
            .O(N__38406),
            .I(\nx.n30 ));
    InMux I__8222 (
            .O(N__38403),
            .I(N__38400));
    LocalMux I__8221 (
            .O(N__38400),
            .I(\nx.n22_adj_604 ));
    CascadeMux I__8220 (
            .O(N__38397),
            .I(N__38393));
    InMux I__8219 (
            .O(N__38396),
            .I(N__38390));
    InMux I__8218 (
            .O(N__38393),
            .I(N__38387));
    LocalMux I__8217 (
            .O(N__38390),
            .I(delay_counter_0));
    LocalMux I__8216 (
            .O(N__38387),
            .I(delay_counter_0));
    InMux I__8215 (
            .O(N__38382),
            .I(bfn_12_26_0_));
    InMux I__8214 (
            .O(N__38379),
            .I(N__38375));
    InMux I__8213 (
            .O(N__38378),
            .I(N__38372));
    LocalMux I__8212 (
            .O(N__38375),
            .I(delay_counter_1));
    LocalMux I__8211 (
            .O(N__38372),
            .I(delay_counter_1));
    InMux I__8210 (
            .O(N__38367),
            .I(n10517));
    InMux I__8209 (
            .O(N__38364),
            .I(N__38360));
    InMux I__8208 (
            .O(N__38363),
            .I(N__38357));
    LocalMux I__8207 (
            .O(N__38360),
            .I(delay_counter_2));
    LocalMux I__8206 (
            .O(N__38357),
            .I(delay_counter_2));
    InMux I__8205 (
            .O(N__38352),
            .I(n10518));
    InMux I__8204 (
            .O(N__38349),
            .I(N__38346));
    LocalMux I__8203 (
            .O(N__38346),
            .I(\nx.n30_adj_640 ));
    CascadeMux I__8202 (
            .O(N__38343),
            .I(\nx.n34_cascade_ ));
    InMux I__8201 (
            .O(N__38340),
            .I(N__38337));
    LocalMux I__8200 (
            .O(N__38337),
            .I(N__38334));
    Odrv4 I__8199 (
            .O(N__38334),
            .I(\nx.n21 ));
    CascadeMux I__8198 (
            .O(N__38331),
            .I(\nx.n2225_cascade_ ));
    InMux I__8197 (
            .O(N__38328),
            .I(N__38325));
    LocalMux I__8196 (
            .O(N__38325),
            .I(N__38322));
    Odrv4 I__8195 (
            .O(N__38322),
            .I(\nx.n2562 ));
    InMux I__8194 (
            .O(N__38319),
            .I(\nx.n10761 ));
    InMux I__8193 (
            .O(N__38316),
            .I(N__38312));
    InMux I__8192 (
            .O(N__38315),
            .I(N__38309));
    LocalMux I__8191 (
            .O(N__38312),
            .I(\nx.n2494 ));
    LocalMux I__8190 (
            .O(N__38309),
            .I(\nx.n2494 ));
    InMux I__8189 (
            .O(N__38304),
            .I(N__38301));
    LocalMux I__8188 (
            .O(N__38301),
            .I(\nx.n2561 ));
    InMux I__8187 (
            .O(N__38298),
            .I(bfn_12_22_0_));
    InMux I__8186 (
            .O(N__38295),
            .I(N__38292));
    LocalMux I__8185 (
            .O(N__38292),
            .I(N__38288));
    InMux I__8184 (
            .O(N__38291),
            .I(N__38285));
    Span4Mux_v I__8183 (
            .O(N__38288),
            .I(N__38279));
    LocalMux I__8182 (
            .O(N__38285),
            .I(N__38279));
    InMux I__8181 (
            .O(N__38284),
            .I(N__38276));
    Odrv4 I__8180 (
            .O(N__38279),
            .I(\nx.n2493 ));
    LocalMux I__8179 (
            .O(N__38276),
            .I(\nx.n2493 ));
    InMux I__8178 (
            .O(N__38271),
            .I(N__38268));
    LocalMux I__8177 (
            .O(N__38268),
            .I(N__38265));
    Span4Mux_h I__8176 (
            .O(N__38265),
            .I(N__38262));
    Odrv4 I__8175 (
            .O(N__38262),
            .I(\nx.n2560 ));
    InMux I__8174 (
            .O(N__38259),
            .I(\nx.n10763 ));
    InMux I__8173 (
            .O(N__38256),
            .I(N__38253));
    LocalMux I__8172 (
            .O(N__38253),
            .I(N__38249));
    InMux I__8171 (
            .O(N__38252),
            .I(N__38245));
    Span4Mux_v I__8170 (
            .O(N__38249),
            .I(N__38242));
    InMux I__8169 (
            .O(N__38248),
            .I(N__38239));
    LocalMux I__8168 (
            .O(N__38245),
            .I(\nx.n2492 ));
    Odrv4 I__8167 (
            .O(N__38242),
            .I(\nx.n2492 ));
    LocalMux I__8166 (
            .O(N__38239),
            .I(\nx.n2492 ));
    InMux I__8165 (
            .O(N__38232),
            .I(N__38229));
    LocalMux I__8164 (
            .O(N__38229),
            .I(N__38226));
    Odrv4 I__8163 (
            .O(N__38226),
            .I(\nx.n2559 ));
    InMux I__8162 (
            .O(N__38223),
            .I(\nx.n10764 ));
    CascadeMux I__8161 (
            .O(N__38220),
            .I(N__38217));
    InMux I__8160 (
            .O(N__38217),
            .I(N__38214));
    LocalMux I__8159 (
            .O(N__38214),
            .I(N__38210));
    InMux I__8158 (
            .O(N__38213),
            .I(N__38207));
    Span4Mux_v I__8157 (
            .O(N__38210),
            .I(N__38204));
    LocalMux I__8156 (
            .O(N__38207),
            .I(\nx.n2491 ));
    Odrv4 I__8155 (
            .O(N__38204),
            .I(\nx.n2491 ));
    InMux I__8154 (
            .O(N__38199),
            .I(N__38196));
    LocalMux I__8153 (
            .O(N__38196),
            .I(N__38193));
    Odrv4 I__8152 (
            .O(N__38193),
            .I(\nx.n2558 ));
    InMux I__8151 (
            .O(N__38190),
            .I(\nx.n10765 ));
    CascadeMux I__8150 (
            .O(N__38187),
            .I(N__38184));
    InMux I__8149 (
            .O(N__38184),
            .I(N__38181));
    LocalMux I__8148 (
            .O(N__38181),
            .I(N__38178));
    Odrv4 I__8147 (
            .O(N__38178),
            .I(\nx.n2557 ));
    InMux I__8146 (
            .O(N__38175),
            .I(\nx.n10766 ));
    InMux I__8145 (
            .O(N__38172),
            .I(\nx.n10767 ));
    InMux I__8144 (
            .O(N__38169),
            .I(N__38165));
    InMux I__8143 (
            .O(N__38168),
            .I(N__38162));
    LocalMux I__8142 (
            .O(N__38165),
            .I(N__38159));
    LocalMux I__8141 (
            .O(N__38162),
            .I(N__38156));
    Span4Mux_v I__8140 (
            .O(N__38159),
            .I(N__38153));
    Span4Mux_h I__8139 (
            .O(N__38156),
            .I(N__38150));
    Odrv4 I__8138 (
            .O(N__38153),
            .I(\nx.n2588 ));
    Odrv4 I__8137 (
            .O(N__38150),
            .I(\nx.n2588 ));
    InMux I__8136 (
            .O(N__38145),
            .I(\nx.n10752 ));
    InMux I__8135 (
            .O(N__38142),
            .I(N__38139));
    LocalMux I__8134 (
            .O(N__38139),
            .I(\nx.n2570 ));
    InMux I__8133 (
            .O(N__38136),
            .I(\nx.n10753 ));
    InMux I__8132 (
            .O(N__38133),
            .I(N__38130));
    LocalMux I__8131 (
            .O(N__38130),
            .I(N__38127));
    Odrv4 I__8130 (
            .O(N__38127),
            .I(\nx.n2569 ));
    InMux I__8129 (
            .O(N__38124),
            .I(bfn_12_21_0_));
    InMux I__8128 (
            .O(N__38121),
            .I(N__38115));
    InMux I__8127 (
            .O(N__38120),
            .I(N__38115));
    LocalMux I__8126 (
            .O(N__38115),
            .I(N__38111));
    CascadeMux I__8125 (
            .O(N__38114),
            .I(N__38108));
    Span4Mux_h I__8124 (
            .O(N__38111),
            .I(N__38105));
    InMux I__8123 (
            .O(N__38108),
            .I(N__38102));
    Odrv4 I__8122 (
            .O(N__38105),
            .I(\nx.n2501 ));
    LocalMux I__8121 (
            .O(N__38102),
            .I(\nx.n2501 ));
    InMux I__8120 (
            .O(N__38097),
            .I(N__38094));
    LocalMux I__8119 (
            .O(N__38094),
            .I(N__38091));
    Odrv4 I__8118 (
            .O(N__38091),
            .I(\nx.n2568 ));
    InMux I__8117 (
            .O(N__38088),
            .I(\nx.n10755 ));
    InMux I__8116 (
            .O(N__38085),
            .I(N__38082));
    LocalMux I__8115 (
            .O(N__38082),
            .I(N__38079));
    Span4Mux_h I__8114 (
            .O(N__38079),
            .I(N__38076));
    Odrv4 I__8113 (
            .O(N__38076),
            .I(\nx.n2567 ));
    InMux I__8112 (
            .O(N__38073),
            .I(\nx.n10756 ));
    CascadeMux I__8111 (
            .O(N__38070),
            .I(N__38067));
    InMux I__8110 (
            .O(N__38067),
            .I(N__38062));
    CascadeMux I__8109 (
            .O(N__38066),
            .I(N__38059));
    InMux I__8108 (
            .O(N__38065),
            .I(N__38056));
    LocalMux I__8107 (
            .O(N__38062),
            .I(N__38053));
    InMux I__8106 (
            .O(N__38059),
            .I(N__38050));
    LocalMux I__8105 (
            .O(N__38056),
            .I(N__38047));
    Span4Mux_v I__8104 (
            .O(N__38053),
            .I(N__38044));
    LocalMux I__8103 (
            .O(N__38050),
            .I(N__38039));
    Span4Mux_v I__8102 (
            .O(N__38047),
            .I(N__38039));
    Odrv4 I__8101 (
            .O(N__38044),
            .I(\nx.n2499 ));
    Odrv4 I__8100 (
            .O(N__38039),
            .I(\nx.n2499 ));
    InMux I__8099 (
            .O(N__38034),
            .I(N__38031));
    LocalMux I__8098 (
            .O(N__38031),
            .I(N__38028));
    Odrv4 I__8097 (
            .O(N__38028),
            .I(\nx.n2566 ));
    InMux I__8096 (
            .O(N__38025),
            .I(\nx.n10757 ));
    CascadeMux I__8095 (
            .O(N__38022),
            .I(N__38019));
    InMux I__8094 (
            .O(N__38019),
            .I(N__38016));
    LocalMux I__8093 (
            .O(N__38016),
            .I(N__38013));
    Odrv4 I__8092 (
            .O(N__38013),
            .I(\nx.n2565 ));
    InMux I__8091 (
            .O(N__38010),
            .I(\nx.n10758 ));
    CascadeMux I__8090 (
            .O(N__38007),
            .I(N__38004));
    InMux I__8089 (
            .O(N__38004),
            .I(N__38000));
    InMux I__8088 (
            .O(N__38003),
            .I(N__37997));
    LocalMux I__8087 (
            .O(N__38000),
            .I(N__37994));
    LocalMux I__8086 (
            .O(N__37997),
            .I(\nx.n2497 ));
    Odrv4 I__8085 (
            .O(N__37994),
            .I(\nx.n2497 ));
    InMux I__8084 (
            .O(N__37989),
            .I(N__37986));
    LocalMux I__8083 (
            .O(N__37986),
            .I(N__37983));
    Span4Mux_h I__8082 (
            .O(N__37983),
            .I(N__37980));
    Odrv4 I__8081 (
            .O(N__37980),
            .I(\nx.n2564 ));
    InMux I__8080 (
            .O(N__37977),
            .I(\nx.n10759 ));
    InMux I__8079 (
            .O(N__37974),
            .I(N__37969));
    CascadeMux I__8078 (
            .O(N__37973),
            .I(N__37966));
    InMux I__8077 (
            .O(N__37972),
            .I(N__37963));
    LocalMux I__8076 (
            .O(N__37969),
            .I(N__37960));
    InMux I__8075 (
            .O(N__37966),
            .I(N__37957));
    LocalMux I__8074 (
            .O(N__37963),
            .I(N__37950));
    Span4Mux_v I__8073 (
            .O(N__37960),
            .I(N__37950));
    LocalMux I__8072 (
            .O(N__37957),
            .I(N__37950));
    Odrv4 I__8071 (
            .O(N__37950),
            .I(\nx.n2496 ));
    CascadeMux I__8070 (
            .O(N__37947),
            .I(N__37944));
    InMux I__8069 (
            .O(N__37944),
            .I(N__37941));
    LocalMux I__8068 (
            .O(N__37941),
            .I(N__37938));
    Odrv4 I__8067 (
            .O(N__37938),
            .I(\nx.n2563 ));
    InMux I__8066 (
            .O(N__37935),
            .I(\nx.n10760 ));
    CascadeMux I__8065 (
            .O(N__37932),
            .I(N__37929));
    InMux I__8064 (
            .O(N__37929),
            .I(N__37925));
    InMux I__8063 (
            .O(N__37928),
            .I(N__37922));
    LocalMux I__8062 (
            .O(N__37925),
            .I(N__37918));
    LocalMux I__8061 (
            .O(N__37922),
            .I(N__37915));
    InMux I__8060 (
            .O(N__37921),
            .I(N__37912));
    Span4Mux_h I__8059 (
            .O(N__37918),
            .I(N__37909));
    Odrv4 I__8058 (
            .O(N__37915),
            .I(\nx.n2605 ));
    LocalMux I__8057 (
            .O(N__37912),
            .I(\nx.n2605 ));
    Odrv4 I__8056 (
            .O(N__37909),
            .I(\nx.n2605 ));
    InMux I__8055 (
            .O(N__37902),
            .I(N__37899));
    LocalMux I__8054 (
            .O(N__37899),
            .I(\nx.n35_adj_639 ));
    InMux I__8053 (
            .O(N__37896),
            .I(N__37893));
    LocalMux I__8052 (
            .O(N__37893),
            .I(N__37888));
    InMux I__8051 (
            .O(N__37892),
            .I(N__37885));
    InMux I__8050 (
            .O(N__37891),
            .I(N__37882));
    Span4Mux_h I__8049 (
            .O(N__37888),
            .I(N__37878));
    LocalMux I__8048 (
            .O(N__37885),
            .I(N__37875));
    LocalMux I__8047 (
            .O(N__37882),
            .I(N__37872));
    InMux I__8046 (
            .O(N__37881),
            .I(N__37869));
    Span4Mux_v I__8045 (
            .O(N__37878),
            .I(N__37866));
    Span4Mux_h I__8044 (
            .O(N__37875),
            .I(N__37863));
    Span4Mux_h I__8043 (
            .O(N__37872),
            .I(N__37860));
    LocalMux I__8042 (
            .O(N__37869),
            .I(N__37854));
    Span4Mux_v I__8041 (
            .O(N__37866),
            .I(N__37854));
    Sp12to4 I__8040 (
            .O(N__37863),
            .I(N__37849));
    Sp12to4 I__8039 (
            .O(N__37860),
            .I(N__37849));
    InMux I__8038 (
            .O(N__37859),
            .I(N__37846));
    Span4Mux_h I__8037 (
            .O(N__37854),
            .I(N__37843));
    Span12Mux_v I__8036 (
            .O(N__37849),
            .I(N__37840));
    LocalMux I__8035 (
            .O(N__37846),
            .I(\nx.bit_ctr_10 ));
    Odrv4 I__8034 (
            .O(N__37843),
            .I(\nx.bit_ctr_10 ));
    Odrv12 I__8033 (
            .O(N__37840),
            .I(\nx.bit_ctr_10 ));
    InMux I__8032 (
            .O(N__37833),
            .I(N__37830));
    LocalMux I__8031 (
            .O(N__37830),
            .I(N__37827));
    Odrv4 I__8030 (
            .O(N__37827),
            .I(\nx.n2577 ));
    InMux I__8029 (
            .O(N__37824),
            .I(bfn_12_20_0_));
    InMux I__8028 (
            .O(N__37821),
            .I(N__37816));
    InMux I__8027 (
            .O(N__37820),
            .I(N__37813));
    CascadeMux I__8026 (
            .O(N__37819),
            .I(N__37810));
    LocalMux I__8025 (
            .O(N__37816),
            .I(N__37807));
    LocalMux I__8024 (
            .O(N__37813),
            .I(N__37804));
    InMux I__8023 (
            .O(N__37810),
            .I(N__37801));
    Span4Mux_h I__8022 (
            .O(N__37807),
            .I(N__37798));
    Span4Mux_v I__8021 (
            .O(N__37804),
            .I(N__37793));
    LocalMux I__8020 (
            .O(N__37801),
            .I(N__37793));
    Odrv4 I__8019 (
            .O(N__37798),
            .I(\nx.n2509 ));
    Odrv4 I__8018 (
            .O(N__37793),
            .I(\nx.n2509 ));
    InMux I__8017 (
            .O(N__37788),
            .I(N__37785));
    LocalMux I__8016 (
            .O(N__37785),
            .I(N__37782));
    Odrv4 I__8015 (
            .O(N__37782),
            .I(\nx.n2576 ));
    InMux I__8014 (
            .O(N__37779),
            .I(\nx.n10747 ));
    InMux I__8013 (
            .O(N__37776),
            .I(\nx.n10748 ));
    InMux I__8012 (
            .O(N__37773),
            .I(N__37770));
    LocalMux I__8011 (
            .O(N__37770),
            .I(\nx.n2574 ));
    InMux I__8010 (
            .O(N__37767),
            .I(\nx.n10749 ));
    InMux I__8009 (
            .O(N__37764),
            .I(N__37761));
    LocalMux I__8008 (
            .O(N__37761),
            .I(\nx.n2573 ));
    InMux I__8007 (
            .O(N__37758),
            .I(\nx.n10750 ));
    CascadeMux I__8006 (
            .O(N__37755),
            .I(N__37751));
    InMux I__8005 (
            .O(N__37754),
            .I(N__37748));
    InMux I__8004 (
            .O(N__37751),
            .I(N__37745));
    LocalMux I__8003 (
            .O(N__37748),
            .I(N__37739));
    LocalMux I__8002 (
            .O(N__37745),
            .I(N__37739));
    CascadeMux I__8001 (
            .O(N__37744),
            .I(N__37736));
    Span4Mux_v I__8000 (
            .O(N__37739),
            .I(N__37733));
    InMux I__7999 (
            .O(N__37736),
            .I(N__37730));
    Odrv4 I__7998 (
            .O(N__37733),
            .I(\nx.n2505 ));
    LocalMux I__7997 (
            .O(N__37730),
            .I(\nx.n2505 ));
    CascadeMux I__7996 (
            .O(N__37725),
            .I(N__37722));
    InMux I__7995 (
            .O(N__37722),
            .I(N__37719));
    LocalMux I__7994 (
            .O(N__37719),
            .I(N__37716));
    Odrv4 I__7993 (
            .O(N__37716),
            .I(\nx.n2572 ));
    InMux I__7992 (
            .O(N__37713),
            .I(\nx.n10751 ));
    InMux I__7991 (
            .O(N__37710),
            .I(N__37707));
    LocalMux I__7990 (
            .O(N__37707),
            .I(\nx.n2571 ));
    CascadeMux I__7989 (
            .O(N__37704),
            .I(N__37701));
    InMux I__7988 (
            .O(N__37701),
            .I(N__37698));
    LocalMux I__7987 (
            .O(N__37698),
            .I(N__37695));
    Span4Mux_v I__7986 (
            .O(N__37695),
            .I(N__37691));
    CascadeMux I__7985 (
            .O(N__37694),
            .I(N__37688));
    Span4Mux_h I__7984 (
            .O(N__37691),
            .I(N__37685));
    InMux I__7983 (
            .O(N__37688),
            .I(N__37682));
    Span4Mux_v I__7982 (
            .O(N__37685),
            .I(N__37676));
    LocalMux I__7981 (
            .O(N__37682),
            .I(N__37676));
    InMux I__7980 (
            .O(N__37681),
            .I(N__37673));
    Odrv4 I__7979 (
            .O(N__37676),
            .I(\nx.n2597 ));
    LocalMux I__7978 (
            .O(N__37673),
            .I(\nx.n2597 ));
    InMux I__7977 (
            .O(N__37668),
            .I(N__37664));
    CascadeMux I__7976 (
            .O(N__37667),
            .I(N__37661));
    LocalMux I__7975 (
            .O(N__37664),
            .I(N__37657));
    InMux I__7974 (
            .O(N__37661),
            .I(N__37654));
    InMux I__7973 (
            .O(N__37660),
            .I(N__37651));
    Span4Mux_h I__7972 (
            .O(N__37657),
            .I(N__37646));
    LocalMux I__7971 (
            .O(N__37654),
            .I(N__37646));
    LocalMux I__7970 (
            .O(N__37651),
            .I(\nx.n2601 ));
    Odrv4 I__7969 (
            .O(N__37646),
            .I(\nx.n2601 ));
    CascadeMux I__7968 (
            .O(N__37641),
            .I(\nx.n2497_cascade_ ));
    CascadeMux I__7967 (
            .O(N__37638),
            .I(\nx.n26_adj_611_cascade_ ));
    InMux I__7966 (
            .O(N__37635),
            .I(N__37632));
    LocalMux I__7965 (
            .O(N__37632),
            .I(N__37629));
    Span4Mux_h I__7964 (
            .O(N__37629),
            .I(N__37626));
    Odrv4 I__7963 (
            .O(N__37626),
            .I(\nx.n33 ));
    CascadeMux I__7962 (
            .O(N__37623),
            .I(\nx.n38_adj_612_cascade_ ));
    CascadeMux I__7961 (
            .O(N__37620),
            .I(\nx.n2522_cascade_ ));
    CascadeMux I__7960 (
            .O(N__37617),
            .I(N__37612));
    InMux I__7959 (
            .O(N__37616),
            .I(N__37607));
    InMux I__7958 (
            .O(N__37615),
            .I(N__37607));
    InMux I__7957 (
            .O(N__37612),
            .I(N__37604));
    LocalMux I__7956 (
            .O(N__37607),
            .I(N__37601));
    LocalMux I__7955 (
            .O(N__37604),
            .I(N__37598));
    Span4Mux_v I__7954 (
            .O(N__37601),
            .I(N__37595));
    Span4Mux_h I__7953 (
            .O(N__37598),
            .I(N__37592));
    Odrv4 I__7952 (
            .O(N__37595),
            .I(\nx.n2600 ));
    Odrv4 I__7951 (
            .O(N__37592),
            .I(\nx.n2600 ));
    CascadeMux I__7950 (
            .O(N__37587),
            .I(n7166_cascade_));
    CascadeMux I__7949 (
            .O(N__37584),
            .I(N__37580));
    InMux I__7948 (
            .O(N__37583),
            .I(N__37577));
    InMux I__7947 (
            .O(N__37580),
            .I(N__37574));
    LocalMux I__7946 (
            .O(N__37577),
            .I(N__37569));
    LocalMux I__7945 (
            .O(N__37574),
            .I(N__37569));
    Odrv4 I__7944 (
            .O(N__37569),
            .I(n6152));
    CascadeMux I__7943 (
            .O(N__37566),
            .I(n8_adj_751_cascade_));
    CascadeMux I__7942 (
            .O(N__37563),
            .I(n7294_cascade_));
    IoInMux I__7941 (
            .O(N__37560),
            .I(N__37557));
    LocalMux I__7940 (
            .O(N__37557),
            .I(N__37554));
    IoSpan4Mux I__7939 (
            .O(N__37554),
            .I(N__37551));
    Span4Mux_s0_h I__7938 (
            .O(N__37551),
            .I(N__37548));
    Sp12to4 I__7937 (
            .O(N__37548),
            .I(N__37545));
    Span12Mux_s11_h I__7936 (
            .O(N__37545),
            .I(N__37541));
    InMux I__7935 (
            .O(N__37544),
            .I(N__37537));
    Span12Mux_v I__7934 (
            .O(N__37541),
            .I(N__37534));
    InMux I__7933 (
            .O(N__37540),
            .I(N__37531));
    LocalMux I__7932 (
            .O(N__37537),
            .I(N__37528));
    Odrv12 I__7931 (
            .O(N__37534),
            .I(pin_out_11));
    LocalMux I__7930 (
            .O(N__37531),
            .I(pin_out_11));
    Odrv4 I__7929 (
            .O(N__37528),
            .I(pin_out_11));
    CascadeMux I__7928 (
            .O(N__37521),
            .I(N__37518));
    InMux I__7927 (
            .O(N__37518),
            .I(N__37514));
    InMux I__7926 (
            .O(N__37517),
            .I(N__37511));
    LocalMux I__7925 (
            .O(N__37514),
            .I(N__37508));
    LocalMux I__7924 (
            .O(N__37511),
            .I(N__37505));
    Span4Mux_h I__7923 (
            .O(N__37508),
            .I(N__37502));
    Span4Mux_h I__7922 (
            .O(N__37505),
            .I(N__37499));
    Odrv4 I__7921 (
            .O(N__37502),
            .I(n6154));
    Odrv4 I__7920 (
            .O(N__37499),
            .I(n6154));
    InMux I__7919 (
            .O(N__37494),
            .I(N__37490));
    InMux I__7918 (
            .O(N__37493),
            .I(N__37487));
    LocalMux I__7917 (
            .O(N__37490),
            .I(N__37482));
    LocalMux I__7916 (
            .O(N__37487),
            .I(N__37482));
    Span4Mux_v I__7915 (
            .O(N__37482),
            .I(N__37477));
    InMux I__7914 (
            .O(N__37481),
            .I(N__37474));
    InMux I__7913 (
            .O(N__37480),
            .I(N__37471));
    Odrv4 I__7912 (
            .O(N__37477),
            .I(n8_adj_744));
    LocalMux I__7911 (
            .O(N__37474),
            .I(n8_adj_744));
    LocalMux I__7910 (
            .O(N__37471),
            .I(n8_adj_744));
    CascadeMux I__7909 (
            .O(N__37464),
            .I(n13048_cascade_));
    InMux I__7908 (
            .O(N__37461),
            .I(N__37458));
    LocalMux I__7907 (
            .O(N__37458),
            .I(N__37455));
    Odrv4 I__7906 (
            .O(N__37455),
            .I(n13264));
    InMux I__7905 (
            .O(N__37452),
            .I(N__37449));
    LocalMux I__7904 (
            .O(N__37449),
            .I(n12091));
    CascadeMux I__7903 (
            .O(N__37446),
            .I(n24_adj_720_cascade_));
    InMux I__7902 (
            .O(N__37443),
            .I(N__37440));
    LocalMux I__7901 (
            .O(N__37440),
            .I(N__37437));
    Odrv4 I__7900 (
            .O(N__37437),
            .I(n11898));
    InMux I__7899 (
            .O(N__37434),
            .I(N__37431));
    LocalMux I__7898 (
            .O(N__37431),
            .I(N__37427));
    CascadeMux I__7897 (
            .O(N__37430),
            .I(N__37424));
    Span4Mux_v I__7896 (
            .O(N__37427),
            .I(N__37420));
    InMux I__7895 (
            .O(N__37424),
            .I(N__37417));
    InMux I__7894 (
            .O(N__37423),
            .I(N__37413));
    IoSpan4Mux I__7893 (
            .O(N__37420),
            .I(N__37408));
    LocalMux I__7892 (
            .O(N__37417),
            .I(N__37408));
    InMux I__7891 (
            .O(N__37416),
            .I(N__37405));
    LocalMux I__7890 (
            .O(N__37413),
            .I(N__37402));
    Span4Mux_s2_h I__7889 (
            .O(N__37408),
            .I(N__37399));
    LocalMux I__7888 (
            .O(N__37405),
            .I(N__37396));
    Span4Mux_v I__7887 (
            .O(N__37402),
            .I(N__37390));
    Span4Mux_v I__7886 (
            .O(N__37399),
            .I(N__37390));
    Span4Mux_v I__7885 (
            .O(N__37396),
            .I(N__37387));
    InMux I__7884 (
            .O(N__37395),
            .I(N__37384));
    Span4Mux_h I__7883 (
            .O(N__37390),
            .I(N__37381));
    Span4Mux_h I__7882 (
            .O(N__37387),
            .I(N__37378));
    LocalMux I__7881 (
            .O(N__37384),
            .I(neopxl_color_7));
    Odrv4 I__7880 (
            .O(N__37381),
            .I(neopxl_color_7));
    Odrv4 I__7879 (
            .O(N__37378),
            .I(neopxl_color_7));
    SRMux I__7878 (
            .O(N__37371),
            .I(N__37368));
    LocalMux I__7877 (
            .O(N__37368),
            .I(N__37365));
    Span4Mux_v I__7876 (
            .O(N__37365),
            .I(N__37362));
    Span4Mux_h I__7875 (
            .O(N__37362),
            .I(N__37359));
    Odrv4 I__7874 (
            .O(N__37359),
            .I(n22_adj_724));
    InMux I__7873 (
            .O(N__37356),
            .I(N__37353));
    LocalMux I__7872 (
            .O(N__37353),
            .I(n17_adj_765));
    CascadeMux I__7871 (
            .O(N__37350),
            .I(n16_adj_764_cascade_));
    InMux I__7870 (
            .O(N__37347),
            .I(N__37344));
    LocalMux I__7869 (
            .O(N__37344),
            .I(N__37341));
    Odrv12 I__7868 (
            .O(N__37341),
            .I(n10978));
    CEMux I__7867 (
            .O(N__37338),
            .I(N__37335));
    LocalMux I__7866 (
            .O(N__37335),
            .I(N__37332));
    Odrv4 I__7865 (
            .O(N__37332),
            .I(n36));
    InMux I__7864 (
            .O(N__37329),
            .I(N__37325));
    InMux I__7863 (
            .O(N__37328),
            .I(N__37322));
    LocalMux I__7862 (
            .O(N__37325),
            .I(N__37317));
    LocalMux I__7861 (
            .O(N__37322),
            .I(N__37317));
    Span4Mux_h I__7860 (
            .O(N__37317),
            .I(N__37313));
    InMux I__7859 (
            .O(N__37316),
            .I(N__37310));
    Odrv4 I__7858 (
            .O(N__37313),
            .I(\nx.n2095 ));
    LocalMux I__7857 (
            .O(N__37310),
            .I(\nx.n2095 ));
    InMux I__7856 (
            .O(N__37305),
            .I(\nx.n10687 ));
    InMux I__7855 (
            .O(N__37302),
            .I(N__37298));
    InMux I__7854 (
            .O(N__37301),
            .I(N__37295));
    LocalMux I__7853 (
            .O(N__37298),
            .I(N__37289));
    LocalMux I__7852 (
            .O(N__37295),
            .I(N__37289));
    InMux I__7851 (
            .O(N__37294),
            .I(N__37286));
    Odrv4 I__7850 (
            .O(N__37289),
            .I(\nx.n2094 ));
    LocalMux I__7849 (
            .O(N__37286),
            .I(\nx.n2094 ));
    InMux I__7848 (
            .O(N__37281),
            .I(bfn_11_25_0_));
    InMux I__7847 (
            .O(N__37278),
            .I(N__37274));
    InMux I__7846 (
            .O(N__37277),
            .I(N__37271));
    LocalMux I__7845 (
            .O(N__37274),
            .I(N__37265));
    LocalMux I__7844 (
            .O(N__37271),
            .I(N__37265));
    InMux I__7843 (
            .O(N__37270),
            .I(N__37262));
    Odrv4 I__7842 (
            .O(N__37265),
            .I(\nx.n2093 ));
    LocalMux I__7841 (
            .O(N__37262),
            .I(\nx.n2093 ));
    CascadeMux I__7840 (
            .O(N__37257),
            .I(N__37239));
    CascadeMux I__7839 (
            .O(N__37256),
            .I(N__37236));
    CascadeMux I__7838 (
            .O(N__37255),
            .I(N__37233));
    CascadeMux I__7837 (
            .O(N__37254),
            .I(N__37230));
    CascadeMux I__7836 (
            .O(N__37253),
            .I(N__37227));
    CascadeMux I__7835 (
            .O(N__37252),
            .I(N__37224));
    CascadeMux I__7834 (
            .O(N__37251),
            .I(N__37221));
    CascadeMux I__7833 (
            .O(N__37250),
            .I(N__37218));
    CascadeMux I__7832 (
            .O(N__37249),
            .I(N__37215));
    CascadeMux I__7831 (
            .O(N__37248),
            .I(N__37212));
    CascadeMux I__7830 (
            .O(N__37247),
            .I(N__37209));
    CascadeMux I__7829 (
            .O(N__37246),
            .I(N__37206));
    CascadeMux I__7828 (
            .O(N__37245),
            .I(N__37203));
    CascadeMux I__7827 (
            .O(N__37244),
            .I(N__37200));
    CascadeMux I__7826 (
            .O(N__37243),
            .I(N__37197));
    CascadeMux I__7825 (
            .O(N__37242),
            .I(N__37194));
    InMux I__7824 (
            .O(N__37239),
            .I(N__37190));
    InMux I__7823 (
            .O(N__37236),
            .I(N__37187));
    InMux I__7822 (
            .O(N__37233),
            .I(N__37178));
    InMux I__7821 (
            .O(N__37230),
            .I(N__37178));
    InMux I__7820 (
            .O(N__37227),
            .I(N__37178));
    InMux I__7819 (
            .O(N__37224),
            .I(N__37178));
    InMux I__7818 (
            .O(N__37221),
            .I(N__37169));
    InMux I__7817 (
            .O(N__37218),
            .I(N__37169));
    InMux I__7816 (
            .O(N__37215),
            .I(N__37169));
    InMux I__7815 (
            .O(N__37212),
            .I(N__37169));
    InMux I__7814 (
            .O(N__37209),
            .I(N__37162));
    InMux I__7813 (
            .O(N__37206),
            .I(N__37162));
    InMux I__7812 (
            .O(N__37203),
            .I(N__37162));
    InMux I__7811 (
            .O(N__37200),
            .I(N__37155));
    InMux I__7810 (
            .O(N__37197),
            .I(N__37155));
    InMux I__7809 (
            .O(N__37194),
            .I(N__37155));
    InMux I__7808 (
            .O(N__37193),
            .I(N__37152));
    LocalMux I__7807 (
            .O(N__37190),
            .I(\nx.n2126 ));
    LocalMux I__7806 (
            .O(N__37187),
            .I(\nx.n2126 ));
    LocalMux I__7805 (
            .O(N__37178),
            .I(\nx.n2126 ));
    LocalMux I__7804 (
            .O(N__37169),
            .I(\nx.n2126 ));
    LocalMux I__7803 (
            .O(N__37162),
            .I(\nx.n2126 ));
    LocalMux I__7802 (
            .O(N__37155),
            .I(\nx.n2126 ));
    LocalMux I__7801 (
            .O(N__37152),
            .I(\nx.n2126 ));
    InMux I__7800 (
            .O(N__37137),
            .I(\nx.n10689 ));
    CascadeMux I__7799 (
            .O(N__37134),
            .I(N__37131));
    InMux I__7798 (
            .O(N__37131),
            .I(N__37128));
    LocalMux I__7797 (
            .O(N__37128),
            .I(n12171));
    InMux I__7796 (
            .O(N__37125),
            .I(N__37122));
    LocalMux I__7795 (
            .O(N__37122),
            .I(n6_adj_761));
    CascadeMux I__7794 (
            .O(N__37119),
            .I(n15_cascade_));
    InMux I__7793 (
            .O(N__37116),
            .I(N__37113));
    LocalMux I__7792 (
            .O(N__37113),
            .I(n14));
    InMux I__7791 (
            .O(N__37110),
            .I(N__37106));
    InMux I__7790 (
            .O(N__37109),
            .I(N__37103));
    LocalMux I__7789 (
            .O(N__37106),
            .I(N__37098));
    LocalMux I__7788 (
            .O(N__37103),
            .I(N__37098));
    Span4Mux_h I__7787 (
            .O(N__37098),
            .I(N__37094));
    InMux I__7786 (
            .O(N__37097),
            .I(N__37091));
    Odrv4 I__7785 (
            .O(N__37094),
            .I(\nx.n2103 ));
    LocalMux I__7784 (
            .O(N__37091),
            .I(\nx.n2103 ));
    InMux I__7783 (
            .O(N__37086),
            .I(\nx.n10679 ));
    InMux I__7782 (
            .O(N__37083),
            .I(N__37078));
    InMux I__7781 (
            .O(N__37082),
            .I(N__37075));
    InMux I__7780 (
            .O(N__37081),
            .I(N__37072));
    LocalMux I__7779 (
            .O(N__37078),
            .I(\nx.n2102 ));
    LocalMux I__7778 (
            .O(N__37075),
            .I(\nx.n2102 ));
    LocalMux I__7777 (
            .O(N__37072),
            .I(\nx.n2102 ));
    InMux I__7776 (
            .O(N__37065),
            .I(bfn_11_24_0_));
    InMux I__7775 (
            .O(N__37062),
            .I(N__37057));
    InMux I__7774 (
            .O(N__37061),
            .I(N__37054));
    InMux I__7773 (
            .O(N__37060),
            .I(N__37051));
    LocalMux I__7772 (
            .O(N__37057),
            .I(\nx.n2101 ));
    LocalMux I__7771 (
            .O(N__37054),
            .I(\nx.n2101 ));
    LocalMux I__7770 (
            .O(N__37051),
            .I(\nx.n2101 ));
    InMux I__7769 (
            .O(N__37044),
            .I(\nx.n10681 ));
    InMux I__7768 (
            .O(N__37041),
            .I(N__37037));
    InMux I__7767 (
            .O(N__37040),
            .I(N__37034));
    LocalMux I__7766 (
            .O(N__37037),
            .I(N__37031));
    LocalMux I__7765 (
            .O(N__37034),
            .I(N__37028));
    Span4Mux_v I__7764 (
            .O(N__37031),
            .I(N__37022));
    Span4Mux_v I__7763 (
            .O(N__37028),
            .I(N__37022));
    InMux I__7762 (
            .O(N__37027),
            .I(N__37019));
    Odrv4 I__7761 (
            .O(N__37022),
            .I(\nx.n2100 ));
    LocalMux I__7760 (
            .O(N__37019),
            .I(\nx.n2100 ));
    InMux I__7759 (
            .O(N__37014),
            .I(\nx.n10682 ));
    InMux I__7758 (
            .O(N__37011),
            .I(N__37007));
    InMux I__7757 (
            .O(N__37010),
            .I(N__37004));
    LocalMux I__7756 (
            .O(N__37007),
            .I(N__36999));
    LocalMux I__7755 (
            .O(N__37004),
            .I(N__36999));
    Span4Mux_h I__7754 (
            .O(N__36999),
            .I(N__36996));
    Odrv4 I__7753 (
            .O(N__36996),
            .I(\nx.n2099 ));
    InMux I__7752 (
            .O(N__36993),
            .I(\nx.n10683 ));
    InMux I__7751 (
            .O(N__36990),
            .I(N__36986));
    InMux I__7750 (
            .O(N__36989),
            .I(N__36983));
    LocalMux I__7749 (
            .O(N__36986),
            .I(N__36980));
    LocalMux I__7748 (
            .O(N__36983),
            .I(N__36977));
    Span4Mux_v I__7747 (
            .O(N__36980),
            .I(N__36971));
    Span4Mux_v I__7746 (
            .O(N__36977),
            .I(N__36971));
    InMux I__7745 (
            .O(N__36976),
            .I(N__36968));
    Odrv4 I__7744 (
            .O(N__36971),
            .I(\nx.n2098 ));
    LocalMux I__7743 (
            .O(N__36968),
            .I(\nx.n2098 ));
    InMux I__7742 (
            .O(N__36963),
            .I(\nx.n10684 ));
    InMux I__7741 (
            .O(N__36960),
            .I(N__36957));
    LocalMux I__7740 (
            .O(N__36957),
            .I(N__36953));
    InMux I__7739 (
            .O(N__36956),
            .I(N__36950));
    Odrv4 I__7738 (
            .O(N__36953),
            .I(\nx.n2097 ));
    LocalMux I__7737 (
            .O(N__36950),
            .I(\nx.n2097 ));
    InMux I__7736 (
            .O(N__36945),
            .I(\nx.n10685 ));
    InMux I__7735 (
            .O(N__36942),
            .I(N__36937));
    InMux I__7734 (
            .O(N__36941),
            .I(N__36934));
    InMux I__7733 (
            .O(N__36940),
            .I(N__36931));
    LocalMux I__7732 (
            .O(N__36937),
            .I(\nx.n2096 ));
    LocalMux I__7731 (
            .O(N__36934),
            .I(\nx.n2096 ));
    LocalMux I__7730 (
            .O(N__36931),
            .I(\nx.n2096 ));
    InMux I__7729 (
            .O(N__36924),
            .I(\nx.n10686 ));
    CascadeMux I__7728 (
            .O(N__36921),
            .I(\nx.n2293_cascade_ ));
    InMux I__7727 (
            .O(N__36918),
            .I(N__36914));
    InMux I__7726 (
            .O(N__36917),
            .I(N__36911));
    LocalMux I__7725 (
            .O(N__36914),
            .I(N__36905));
    LocalMux I__7724 (
            .O(N__36911),
            .I(N__36905));
    InMux I__7723 (
            .O(N__36910),
            .I(N__36902));
    Span4Mux_v I__7722 (
            .O(N__36905),
            .I(N__36896));
    LocalMux I__7721 (
            .O(N__36902),
            .I(N__36896));
    InMux I__7720 (
            .O(N__36901),
            .I(N__36892));
    Span4Mux_h I__7719 (
            .O(N__36896),
            .I(N__36889));
    InMux I__7718 (
            .O(N__36895),
            .I(N__36886));
    LocalMux I__7717 (
            .O(N__36892),
            .I(N__36881));
    Span4Mux_v I__7716 (
            .O(N__36889),
            .I(N__36881));
    LocalMux I__7715 (
            .O(N__36886),
            .I(\nx.bit_ctr_14 ));
    Odrv4 I__7714 (
            .O(N__36881),
            .I(\nx.bit_ctr_14 ));
    InMux I__7713 (
            .O(N__36876),
            .I(bfn_11_23_0_));
    CascadeMux I__7712 (
            .O(N__36873),
            .I(N__36870));
    InMux I__7711 (
            .O(N__36870),
            .I(N__36865));
    InMux I__7710 (
            .O(N__36869),
            .I(N__36862));
    InMux I__7709 (
            .O(N__36868),
            .I(N__36859));
    LocalMux I__7708 (
            .O(N__36865),
            .I(N__36856));
    LocalMux I__7707 (
            .O(N__36862),
            .I(\nx.n2109 ));
    LocalMux I__7706 (
            .O(N__36859),
            .I(\nx.n2109 ));
    Odrv4 I__7705 (
            .O(N__36856),
            .I(\nx.n2109 ));
    CascadeMux I__7704 (
            .O(N__36849),
            .I(N__36845));
    CascadeMux I__7703 (
            .O(N__36848),
            .I(N__36842));
    InMux I__7702 (
            .O(N__36845),
            .I(N__36839));
    InMux I__7701 (
            .O(N__36842),
            .I(N__36836));
    LocalMux I__7700 (
            .O(N__36839),
            .I(\nx.n13436 ));
    LocalMux I__7699 (
            .O(N__36836),
            .I(\nx.n13436 ));
    InMux I__7698 (
            .O(N__36831),
            .I(\nx.n10673 ));
    InMux I__7697 (
            .O(N__36828),
            .I(N__36823));
    InMux I__7696 (
            .O(N__36827),
            .I(N__36820));
    InMux I__7695 (
            .O(N__36826),
            .I(N__36817));
    LocalMux I__7694 (
            .O(N__36823),
            .I(\nx.n2108 ));
    LocalMux I__7693 (
            .O(N__36820),
            .I(\nx.n2108 ));
    LocalMux I__7692 (
            .O(N__36817),
            .I(\nx.n2108 ));
    InMux I__7691 (
            .O(N__36810),
            .I(\nx.n10674 ));
    InMux I__7690 (
            .O(N__36807),
            .I(N__36803));
    InMux I__7689 (
            .O(N__36806),
            .I(N__36800));
    LocalMux I__7688 (
            .O(N__36803),
            .I(\nx.n2107 ));
    LocalMux I__7687 (
            .O(N__36800),
            .I(\nx.n2107 ));
    InMux I__7686 (
            .O(N__36795),
            .I(\nx.n10675 ));
    InMux I__7685 (
            .O(N__36792),
            .I(N__36787));
    InMux I__7684 (
            .O(N__36791),
            .I(N__36784));
    InMux I__7683 (
            .O(N__36790),
            .I(N__36781));
    LocalMux I__7682 (
            .O(N__36787),
            .I(\nx.n2106 ));
    LocalMux I__7681 (
            .O(N__36784),
            .I(\nx.n2106 ));
    LocalMux I__7680 (
            .O(N__36781),
            .I(\nx.n2106 ));
    InMux I__7679 (
            .O(N__36774),
            .I(\nx.n10676 ));
    InMux I__7678 (
            .O(N__36771),
            .I(N__36767));
    InMux I__7677 (
            .O(N__36770),
            .I(N__36764));
    LocalMux I__7676 (
            .O(N__36767),
            .I(N__36759));
    LocalMux I__7675 (
            .O(N__36764),
            .I(N__36759));
    Span4Mux_h I__7674 (
            .O(N__36759),
            .I(N__36756));
    Odrv4 I__7673 (
            .O(N__36756),
            .I(\nx.n2105 ));
    InMux I__7672 (
            .O(N__36753),
            .I(\nx.n10677 ));
    InMux I__7671 (
            .O(N__36750),
            .I(N__36746));
    InMux I__7670 (
            .O(N__36749),
            .I(N__36743));
    LocalMux I__7669 (
            .O(N__36746),
            .I(N__36738));
    LocalMux I__7668 (
            .O(N__36743),
            .I(N__36738));
    Span4Mux_h I__7667 (
            .O(N__36738),
            .I(N__36734));
    InMux I__7666 (
            .O(N__36737),
            .I(N__36731));
    Odrv4 I__7665 (
            .O(N__36734),
            .I(\nx.n2104 ));
    LocalMux I__7664 (
            .O(N__36731),
            .I(\nx.n2104 ));
    InMux I__7663 (
            .O(N__36726),
            .I(\nx.n10678 ));
    CascadeMux I__7662 (
            .O(N__36723),
            .I(\nx.n2296_cascade_ ));
    CascadeMux I__7661 (
            .O(N__36720),
            .I(\nx.n2395_cascade_ ));
    CascadeMux I__7660 (
            .O(N__36717),
            .I(\nx.n2494_cascade_ ));
    InMux I__7659 (
            .O(N__36714),
            .I(N__36709));
    InMux I__7658 (
            .O(N__36713),
            .I(N__36706));
    InMux I__7657 (
            .O(N__36712),
            .I(N__36703));
    LocalMux I__7656 (
            .O(N__36709),
            .I(N__36700));
    LocalMux I__7655 (
            .O(N__36706),
            .I(N__36697));
    LocalMux I__7654 (
            .O(N__36703),
            .I(\nx.n2593 ));
    Odrv4 I__7653 (
            .O(N__36700),
            .I(\nx.n2593 ));
    Odrv4 I__7652 (
            .O(N__36697),
            .I(\nx.n2593 ));
    CascadeMux I__7651 (
            .O(N__36690),
            .I(\nx.n2504_cascade_ ));
    InMux I__7650 (
            .O(N__36687),
            .I(N__36683));
    CascadeMux I__7649 (
            .O(N__36686),
            .I(N__36680));
    LocalMux I__7648 (
            .O(N__36683),
            .I(N__36677));
    InMux I__7647 (
            .O(N__36680),
            .I(N__36673));
    Span4Mux_h I__7646 (
            .O(N__36677),
            .I(N__36670));
    InMux I__7645 (
            .O(N__36676),
            .I(N__36667));
    LocalMux I__7644 (
            .O(N__36673),
            .I(N__36664));
    Odrv4 I__7643 (
            .O(N__36670),
            .I(\nx.n2603 ));
    LocalMux I__7642 (
            .O(N__36667),
            .I(\nx.n2603 ));
    Odrv4 I__7641 (
            .O(N__36664),
            .I(\nx.n2603 ));
    CascadeMux I__7640 (
            .O(N__36657),
            .I(N__36653));
    CascadeMux I__7639 (
            .O(N__36656),
            .I(N__36649));
    InMux I__7638 (
            .O(N__36653),
            .I(N__36646));
    InMux I__7637 (
            .O(N__36652),
            .I(N__36641));
    InMux I__7636 (
            .O(N__36649),
            .I(N__36641));
    LocalMux I__7635 (
            .O(N__36646),
            .I(\nx.n2589 ));
    LocalMux I__7634 (
            .O(N__36641),
            .I(\nx.n2589 ));
    CascadeMux I__7633 (
            .O(N__36636),
            .I(N__36633));
    InMux I__7632 (
            .O(N__36633),
            .I(N__36630));
    LocalMux I__7631 (
            .O(N__36630),
            .I(N__36626));
    InMux I__7630 (
            .O(N__36629),
            .I(N__36622));
    Span4Mux_h I__7629 (
            .O(N__36626),
            .I(N__36619));
    InMux I__7628 (
            .O(N__36625),
            .I(N__36616));
    LocalMux I__7627 (
            .O(N__36622),
            .I(\nx.n2688 ));
    Odrv4 I__7626 (
            .O(N__36619),
            .I(\nx.n2688 ));
    LocalMux I__7625 (
            .O(N__36616),
            .I(\nx.n2688 ));
    CascadeMux I__7624 (
            .O(N__36609),
            .I(N__36606));
    InMux I__7623 (
            .O(N__36606),
            .I(N__36602));
    CascadeMux I__7622 (
            .O(N__36605),
            .I(N__36597));
    LocalMux I__7621 (
            .O(N__36602),
            .I(N__36587));
    InMux I__7620 (
            .O(N__36601),
            .I(N__36583));
    InMux I__7619 (
            .O(N__36600),
            .I(N__36576));
    InMux I__7618 (
            .O(N__36597),
            .I(N__36576));
    InMux I__7617 (
            .O(N__36596),
            .I(N__36576));
    InMux I__7616 (
            .O(N__36595),
            .I(N__36570));
    InMux I__7615 (
            .O(N__36594),
            .I(N__36570));
    CascadeMux I__7614 (
            .O(N__36593),
            .I(N__36566));
    CascadeMux I__7613 (
            .O(N__36592),
            .I(N__36561));
    CascadeMux I__7612 (
            .O(N__36591),
            .I(N__36557));
    CascadeMux I__7611 (
            .O(N__36590),
            .I(N__36551));
    Span4Mux_v I__7610 (
            .O(N__36587),
            .I(N__36545));
    InMux I__7609 (
            .O(N__36586),
            .I(N__36542));
    LocalMux I__7608 (
            .O(N__36583),
            .I(N__36537));
    LocalMux I__7607 (
            .O(N__36576),
            .I(N__36537));
    InMux I__7606 (
            .O(N__36575),
            .I(N__36534));
    LocalMux I__7605 (
            .O(N__36570),
            .I(N__36531));
    InMux I__7604 (
            .O(N__36569),
            .I(N__36528));
    InMux I__7603 (
            .O(N__36566),
            .I(N__36523));
    InMux I__7602 (
            .O(N__36565),
            .I(N__36523));
    InMux I__7601 (
            .O(N__36564),
            .I(N__36508));
    InMux I__7600 (
            .O(N__36561),
            .I(N__36508));
    InMux I__7599 (
            .O(N__36560),
            .I(N__36508));
    InMux I__7598 (
            .O(N__36557),
            .I(N__36508));
    InMux I__7597 (
            .O(N__36556),
            .I(N__36508));
    InMux I__7596 (
            .O(N__36555),
            .I(N__36508));
    InMux I__7595 (
            .O(N__36554),
            .I(N__36508));
    InMux I__7594 (
            .O(N__36551),
            .I(N__36499));
    InMux I__7593 (
            .O(N__36550),
            .I(N__36499));
    InMux I__7592 (
            .O(N__36549),
            .I(N__36499));
    InMux I__7591 (
            .O(N__36548),
            .I(N__36499));
    Sp12to4 I__7590 (
            .O(N__36545),
            .I(N__36494));
    LocalMux I__7589 (
            .O(N__36542),
            .I(N__36494));
    Odrv4 I__7588 (
            .O(N__36537),
            .I(\nx.n2720 ));
    LocalMux I__7587 (
            .O(N__36534),
            .I(\nx.n2720 ));
    Odrv12 I__7586 (
            .O(N__36531),
            .I(\nx.n2720 ));
    LocalMux I__7585 (
            .O(N__36528),
            .I(\nx.n2720 ));
    LocalMux I__7584 (
            .O(N__36523),
            .I(\nx.n2720 ));
    LocalMux I__7583 (
            .O(N__36508),
            .I(\nx.n2720 ));
    LocalMux I__7582 (
            .O(N__36499),
            .I(\nx.n2720 ));
    Odrv12 I__7581 (
            .O(N__36494),
            .I(\nx.n2720 ));
    InMux I__7580 (
            .O(N__36477),
            .I(N__36474));
    LocalMux I__7579 (
            .O(N__36474),
            .I(N__36471));
    Span4Mux_h I__7578 (
            .O(N__36471),
            .I(N__36468));
    Odrv4 I__7577 (
            .O(N__36468),
            .I(\nx.n2755 ));
    CascadeMux I__7576 (
            .O(N__36465),
            .I(N__36462));
    InMux I__7575 (
            .O(N__36462),
            .I(N__36459));
    LocalMux I__7574 (
            .O(N__36459),
            .I(N__36454));
    InMux I__7573 (
            .O(N__36458),
            .I(N__36449));
    InMux I__7572 (
            .O(N__36457),
            .I(N__36449));
    Span4Mux_h I__7571 (
            .O(N__36454),
            .I(N__36444));
    LocalMux I__7570 (
            .O(N__36449),
            .I(N__36444));
    Span4Mux_h I__7569 (
            .O(N__36444),
            .I(N__36441));
    Odrv4 I__7568 (
            .O(N__36441),
            .I(\nx.n2787 ));
    CascadeMux I__7567 (
            .O(N__36438),
            .I(N__36435));
    InMux I__7566 (
            .O(N__36435),
            .I(N__36431));
    CascadeMux I__7565 (
            .O(N__36434),
            .I(N__36428));
    LocalMux I__7564 (
            .O(N__36431),
            .I(N__36424));
    InMux I__7563 (
            .O(N__36428),
            .I(N__36421));
    InMux I__7562 (
            .O(N__36427),
            .I(N__36418));
    Odrv12 I__7561 (
            .O(N__36424),
            .I(\nx.n2590 ));
    LocalMux I__7560 (
            .O(N__36421),
            .I(\nx.n2590 ));
    LocalMux I__7559 (
            .O(N__36418),
            .I(\nx.n2590 ));
    InMux I__7558 (
            .O(N__36411),
            .I(N__36407));
    CascadeMux I__7557 (
            .O(N__36410),
            .I(N__36404));
    LocalMux I__7556 (
            .O(N__36407),
            .I(N__36400));
    InMux I__7555 (
            .O(N__36404),
            .I(N__36397));
    InMux I__7554 (
            .O(N__36403),
            .I(N__36394));
    Odrv4 I__7553 (
            .O(N__36400),
            .I(\nx.n2591 ));
    LocalMux I__7552 (
            .O(N__36397),
            .I(\nx.n2591 ));
    LocalMux I__7551 (
            .O(N__36394),
            .I(\nx.n2591 ));
    InMux I__7550 (
            .O(N__36387),
            .I(N__36383));
    CascadeMux I__7549 (
            .O(N__36386),
            .I(N__36380));
    LocalMux I__7548 (
            .O(N__36383),
            .I(N__36377));
    InMux I__7547 (
            .O(N__36380),
            .I(N__36374));
    Odrv4 I__7546 (
            .O(N__36377),
            .I(\nx.n2596 ));
    LocalMux I__7545 (
            .O(N__36374),
            .I(\nx.n2596 ));
    InMux I__7544 (
            .O(N__36369),
            .I(N__36366));
    LocalMux I__7543 (
            .O(N__36366),
            .I(N__36362));
    CascadeMux I__7542 (
            .O(N__36365),
            .I(N__36358));
    Span4Mux_h I__7541 (
            .O(N__36362),
            .I(N__36355));
    InMux I__7540 (
            .O(N__36361),
            .I(N__36352));
    InMux I__7539 (
            .O(N__36358),
            .I(N__36349));
    Odrv4 I__7538 (
            .O(N__36355),
            .I(\nx.n2599 ));
    LocalMux I__7537 (
            .O(N__36352),
            .I(\nx.n2599 ));
    LocalMux I__7536 (
            .O(N__36349),
            .I(\nx.n2599 ));
    CascadeMux I__7535 (
            .O(N__36342),
            .I(\nx.n2596_cascade_ ));
    InMux I__7534 (
            .O(N__36339),
            .I(N__36336));
    LocalMux I__7533 (
            .O(N__36336),
            .I(N__36332));
    CascadeMux I__7532 (
            .O(N__36335),
            .I(N__36328));
    Span4Mux_h I__7531 (
            .O(N__36332),
            .I(N__36325));
    InMux I__7530 (
            .O(N__36331),
            .I(N__36322));
    InMux I__7529 (
            .O(N__36328),
            .I(N__36319));
    Odrv4 I__7528 (
            .O(N__36325),
            .I(\nx.n2604 ));
    LocalMux I__7527 (
            .O(N__36322),
            .I(\nx.n2604 ));
    LocalMux I__7526 (
            .O(N__36319),
            .I(\nx.n2604 ));
    InMux I__7525 (
            .O(N__36312),
            .I(N__36309));
    LocalMux I__7524 (
            .O(N__36309),
            .I(\nx.n37 ));
    InMux I__7523 (
            .O(N__36306),
            .I(N__36303));
    LocalMux I__7522 (
            .O(N__36303),
            .I(N__36298));
    CascadeMux I__7521 (
            .O(N__36302),
            .I(N__36295));
    CascadeMux I__7520 (
            .O(N__36301),
            .I(N__36292));
    Span4Mux_v I__7519 (
            .O(N__36298),
            .I(N__36289));
    InMux I__7518 (
            .O(N__36295),
            .I(N__36286));
    InMux I__7517 (
            .O(N__36292),
            .I(N__36283));
    Odrv4 I__7516 (
            .O(N__36289),
            .I(\nx.n2598 ));
    LocalMux I__7515 (
            .O(N__36286),
            .I(\nx.n2598 ));
    LocalMux I__7514 (
            .O(N__36283),
            .I(\nx.n2598 ));
    InMux I__7513 (
            .O(N__36276),
            .I(N__36273));
    LocalMux I__7512 (
            .O(N__36273),
            .I(\nx.n38 ));
    CascadeMux I__7511 (
            .O(N__36270),
            .I(N__36267));
    InMux I__7510 (
            .O(N__36267),
            .I(N__36264));
    LocalMux I__7509 (
            .O(N__36264),
            .I(N__36260));
    CascadeMux I__7508 (
            .O(N__36263),
            .I(N__36256));
    Span4Mux_h I__7507 (
            .O(N__36260),
            .I(N__36253));
    InMux I__7506 (
            .O(N__36259),
            .I(N__36250));
    InMux I__7505 (
            .O(N__36256),
            .I(N__36247));
    Odrv4 I__7504 (
            .O(N__36253),
            .I(\nx.n2602 ));
    LocalMux I__7503 (
            .O(N__36250),
            .I(\nx.n2602 ));
    LocalMux I__7502 (
            .O(N__36247),
            .I(\nx.n2602 ));
    CascadeMux I__7501 (
            .O(N__36240),
            .I(N__36237));
    InMux I__7500 (
            .O(N__36237),
            .I(N__36233));
    InMux I__7499 (
            .O(N__36236),
            .I(N__36230));
    LocalMux I__7498 (
            .O(N__36233),
            .I(N__36227));
    LocalMux I__7497 (
            .O(N__36230),
            .I(\nx.n2606 ));
    Odrv4 I__7496 (
            .O(N__36227),
            .I(\nx.n2606 ));
    InMux I__7495 (
            .O(N__36222),
            .I(N__36219));
    LocalMux I__7494 (
            .O(N__36219),
            .I(N__36216));
    Odrv4 I__7493 (
            .O(N__36216),
            .I(\nx.n2673 ));
    CascadeMux I__7492 (
            .O(N__36213),
            .I(\nx.n2606_cascade_ ));
    CascadeMux I__7491 (
            .O(N__36210),
            .I(N__36203));
    CascadeMux I__7490 (
            .O(N__36209),
            .I(N__36200));
    InMux I__7489 (
            .O(N__36208),
            .I(N__36188));
    InMux I__7488 (
            .O(N__36207),
            .I(N__36185));
    InMux I__7487 (
            .O(N__36206),
            .I(N__36176));
    InMux I__7486 (
            .O(N__36203),
            .I(N__36176));
    InMux I__7485 (
            .O(N__36200),
            .I(N__36176));
    InMux I__7484 (
            .O(N__36199),
            .I(N__36176));
    CascadeMux I__7483 (
            .O(N__36198),
            .I(N__36173));
    CascadeMux I__7482 (
            .O(N__36197),
            .I(N__36167));
    CascadeMux I__7481 (
            .O(N__36196),
            .I(N__36163));
    CascadeMux I__7480 (
            .O(N__36195),
            .I(N__36160));
    CascadeMux I__7479 (
            .O(N__36194),
            .I(N__36155));
    CascadeMux I__7478 (
            .O(N__36193),
            .I(N__36152));
    CascadeMux I__7477 (
            .O(N__36192),
            .I(N__36148));
    CascadeMux I__7476 (
            .O(N__36191),
            .I(N__36145));
    LocalMux I__7475 (
            .O(N__36188),
            .I(N__36141));
    LocalMux I__7474 (
            .O(N__36185),
            .I(N__36136));
    LocalMux I__7473 (
            .O(N__36176),
            .I(N__36136));
    InMux I__7472 (
            .O(N__36173),
            .I(N__36133));
    InMux I__7471 (
            .O(N__36172),
            .I(N__36130));
    InMux I__7470 (
            .O(N__36171),
            .I(N__36121));
    InMux I__7469 (
            .O(N__36170),
            .I(N__36121));
    InMux I__7468 (
            .O(N__36167),
            .I(N__36121));
    InMux I__7467 (
            .O(N__36166),
            .I(N__36121));
    InMux I__7466 (
            .O(N__36163),
            .I(N__36114));
    InMux I__7465 (
            .O(N__36160),
            .I(N__36114));
    InMux I__7464 (
            .O(N__36159),
            .I(N__36114));
    InMux I__7463 (
            .O(N__36158),
            .I(N__36099));
    InMux I__7462 (
            .O(N__36155),
            .I(N__36099));
    InMux I__7461 (
            .O(N__36152),
            .I(N__36099));
    InMux I__7460 (
            .O(N__36151),
            .I(N__36099));
    InMux I__7459 (
            .O(N__36148),
            .I(N__36099));
    InMux I__7458 (
            .O(N__36145),
            .I(N__36099));
    InMux I__7457 (
            .O(N__36144),
            .I(N__36099));
    Span4Mux_v I__7456 (
            .O(N__36141),
            .I(N__36094));
    Span4Mux_v I__7455 (
            .O(N__36136),
            .I(N__36094));
    LocalMux I__7454 (
            .O(N__36133),
            .I(\nx.n2621 ));
    LocalMux I__7453 (
            .O(N__36130),
            .I(\nx.n2621 ));
    LocalMux I__7452 (
            .O(N__36121),
            .I(\nx.n2621 ));
    LocalMux I__7451 (
            .O(N__36114),
            .I(\nx.n2621 ));
    LocalMux I__7450 (
            .O(N__36099),
            .I(\nx.n2621 ));
    Odrv4 I__7449 (
            .O(N__36094),
            .I(\nx.n2621 ));
    CascadeMux I__7448 (
            .O(N__36081),
            .I(N__36077));
    InMux I__7447 (
            .O(N__36080),
            .I(N__36074));
    InMux I__7446 (
            .O(N__36077),
            .I(N__36071));
    LocalMux I__7445 (
            .O(N__36074),
            .I(N__36068));
    LocalMux I__7444 (
            .O(N__36071),
            .I(N__36065));
    Odrv4 I__7443 (
            .O(N__36068),
            .I(\nx.n2705 ));
    Odrv12 I__7442 (
            .O(N__36065),
            .I(\nx.n2705 ));
    InMux I__7441 (
            .O(N__36060),
            .I(N__36057));
    LocalMux I__7440 (
            .O(N__36057),
            .I(N__36054));
    Odrv12 I__7439 (
            .O(N__36054),
            .I(\nx.n2772 ));
    CascadeMux I__7438 (
            .O(N__36051),
            .I(\nx.n2705_cascade_ ));
    CascadeMux I__7437 (
            .O(N__36048),
            .I(N__36044));
    CascadeMux I__7436 (
            .O(N__36047),
            .I(N__36040));
    InMux I__7435 (
            .O(N__36044),
            .I(N__36037));
    InMux I__7434 (
            .O(N__36043),
            .I(N__36034));
    InMux I__7433 (
            .O(N__36040),
            .I(N__36031));
    LocalMux I__7432 (
            .O(N__36037),
            .I(N__36028));
    LocalMux I__7431 (
            .O(N__36034),
            .I(N__36025));
    LocalMux I__7430 (
            .O(N__36031),
            .I(N__36022));
    Span4Mux_v I__7429 (
            .O(N__36028),
            .I(N__36015));
    Span4Mux_v I__7428 (
            .O(N__36025),
            .I(N__36015));
    Span4Mux_h I__7427 (
            .O(N__36022),
            .I(N__36015));
    Span4Mux_h I__7426 (
            .O(N__36015),
            .I(N__36012));
    Odrv4 I__7425 (
            .O(N__36012),
            .I(\nx.n2804 ));
    InMux I__7424 (
            .O(N__36009),
            .I(N__36005));
    CascadeMux I__7423 (
            .O(N__36008),
            .I(N__36001));
    LocalMux I__7422 (
            .O(N__36005),
            .I(N__35998));
    InMux I__7421 (
            .O(N__36004),
            .I(N__35995));
    InMux I__7420 (
            .O(N__36001),
            .I(N__35992));
    Span4Mux_h I__7419 (
            .O(N__35998),
            .I(N__35989));
    LocalMux I__7418 (
            .O(N__35995),
            .I(\nx.n2594 ));
    LocalMux I__7417 (
            .O(N__35992),
            .I(\nx.n2594 ));
    Odrv4 I__7416 (
            .O(N__35989),
            .I(\nx.n2594 ));
    CascadeMux I__7415 (
            .O(N__35982),
            .I(N__35978));
    InMux I__7414 (
            .O(N__35981),
            .I(N__35975));
    InMux I__7413 (
            .O(N__35978),
            .I(N__35972));
    LocalMux I__7412 (
            .O(N__35975),
            .I(n6156));
    LocalMux I__7411 (
            .O(N__35972),
            .I(n6156));
    CascadeMux I__7410 (
            .O(N__35967),
            .I(n7266_cascade_));
    IoInMux I__7409 (
            .O(N__35964),
            .I(N__35961));
    LocalMux I__7408 (
            .O(N__35961),
            .I(N__35958));
    Span4Mux_s2_h I__7407 (
            .O(N__35958),
            .I(N__35955));
    Span4Mux_h I__7406 (
            .O(N__35955),
            .I(N__35952));
    Span4Mux_h I__7405 (
            .O(N__35952),
            .I(N__35948));
    InMux I__7404 (
            .O(N__35951),
            .I(N__35944));
    Sp12to4 I__7403 (
            .O(N__35948),
            .I(N__35941));
    InMux I__7402 (
            .O(N__35947),
            .I(N__35938));
    LocalMux I__7401 (
            .O(N__35944),
            .I(N__35935));
    Odrv12 I__7400 (
            .O(N__35941),
            .I(pin_out_4));
    LocalMux I__7399 (
            .O(N__35938),
            .I(pin_out_4));
    Odrv4 I__7398 (
            .O(N__35935),
            .I(pin_out_4));
    InMux I__7397 (
            .O(N__35928),
            .I(N__35925));
    LocalMux I__7396 (
            .O(N__35925),
            .I(N__35921));
    CascadeMux I__7395 (
            .O(N__35924),
            .I(N__35918));
    Span4Mux_h I__7394 (
            .O(N__35921),
            .I(N__35915));
    InMux I__7393 (
            .O(N__35918),
            .I(N__35912));
    Odrv4 I__7392 (
            .O(N__35915),
            .I(\nx.n2609 ));
    LocalMux I__7391 (
            .O(N__35912),
            .I(\nx.n2609 ));
    InMux I__7390 (
            .O(N__35907),
            .I(N__35903));
    InMux I__7389 (
            .O(N__35906),
            .I(N__35900));
    LocalMux I__7388 (
            .O(N__35903),
            .I(N__35896));
    LocalMux I__7387 (
            .O(N__35900),
            .I(N__35893));
    InMux I__7386 (
            .O(N__35899),
            .I(N__35890));
    Span4Mux_v I__7385 (
            .O(N__35896),
            .I(N__35887));
    Span4Mux_h I__7384 (
            .O(N__35893),
            .I(N__35882));
    LocalMux I__7383 (
            .O(N__35890),
            .I(N__35882));
    Sp12to4 I__7382 (
            .O(N__35887),
            .I(N__35877));
    Sp12to4 I__7381 (
            .O(N__35882),
            .I(N__35874));
    InMux I__7380 (
            .O(N__35881),
            .I(N__35871));
    InMux I__7379 (
            .O(N__35880),
            .I(N__35868));
    Span12Mux_h I__7378 (
            .O(N__35877),
            .I(N__35865));
    Span12Mux_v I__7377 (
            .O(N__35874),
            .I(N__35862));
    LocalMux I__7376 (
            .O(N__35871),
            .I(\nx.bit_ctr_9 ));
    LocalMux I__7375 (
            .O(N__35868),
            .I(\nx.bit_ctr_9 ));
    Odrv12 I__7374 (
            .O(N__35865),
            .I(\nx.bit_ctr_9 ));
    Odrv12 I__7373 (
            .O(N__35862),
            .I(\nx.bit_ctr_9 ));
    CascadeMux I__7372 (
            .O(N__35853),
            .I(\nx.n2609_cascade_ ));
    CascadeMux I__7371 (
            .O(N__35850),
            .I(\nx.n28_adj_599_cascade_ ));
    InMux I__7370 (
            .O(N__35847),
            .I(N__35844));
    LocalMux I__7369 (
            .O(N__35844),
            .I(N__35841));
    Span4Mux_h I__7368 (
            .O(N__35841),
            .I(N__35838));
    Odrv4 I__7367 (
            .O(N__35838),
            .I(\nx.n35 ));
    InMux I__7366 (
            .O(N__35835),
            .I(N__35832));
    LocalMux I__7365 (
            .O(N__35832),
            .I(N__35829));
    Odrv4 I__7364 (
            .O(N__35829),
            .I(\nx.n40 ));
    InMux I__7363 (
            .O(N__35826),
            .I(N__35822));
    CascadeMux I__7362 (
            .O(N__35825),
            .I(N__35818));
    LocalMux I__7361 (
            .O(N__35822),
            .I(N__35815));
    InMux I__7360 (
            .O(N__35821),
            .I(N__35812));
    InMux I__7359 (
            .O(N__35818),
            .I(N__35809));
    Odrv12 I__7358 (
            .O(N__35815),
            .I(\nx.n2608 ));
    LocalMux I__7357 (
            .O(N__35812),
            .I(\nx.n2608 ));
    LocalMux I__7356 (
            .O(N__35809),
            .I(\nx.n2608 ));
    IoInMux I__7355 (
            .O(N__35802),
            .I(N__35797));
    IoInMux I__7354 (
            .O(N__35801),
            .I(N__35790));
    IoInMux I__7353 (
            .O(N__35800),
            .I(N__35787));
    LocalMux I__7352 (
            .O(N__35797),
            .I(N__35784));
    IoInMux I__7351 (
            .O(N__35796),
            .I(N__35779));
    IoInMux I__7350 (
            .O(N__35795),
            .I(N__35776));
    IoInMux I__7349 (
            .O(N__35794),
            .I(N__35773));
    IoInMux I__7348 (
            .O(N__35793),
            .I(N__35769));
    LocalMux I__7347 (
            .O(N__35790),
            .I(N__35761));
    LocalMux I__7346 (
            .O(N__35787),
            .I(N__35761));
    IoSpan4Mux I__7345 (
            .O(N__35784),
            .I(N__35761));
    IoInMux I__7344 (
            .O(N__35783),
            .I(N__35758));
    IoInMux I__7343 (
            .O(N__35782),
            .I(N__35755));
    LocalMux I__7342 (
            .O(N__35779),
            .I(N__35750));
    LocalMux I__7341 (
            .O(N__35776),
            .I(N__35750));
    LocalMux I__7340 (
            .O(N__35773),
            .I(N__35747));
    IoInMux I__7339 (
            .O(N__35772),
            .I(N__35744));
    LocalMux I__7338 (
            .O(N__35769),
            .I(N__35741));
    IoInMux I__7337 (
            .O(N__35768),
            .I(N__35738));
    IoSpan4Mux I__7336 (
            .O(N__35761),
            .I(N__35726));
    LocalMux I__7335 (
            .O(N__35758),
            .I(N__35726));
    LocalMux I__7334 (
            .O(N__35755),
            .I(N__35726));
    IoSpan4Mux I__7333 (
            .O(N__35750),
            .I(N__35716));
    IoSpan4Mux I__7332 (
            .O(N__35747),
            .I(N__35716));
    LocalMux I__7331 (
            .O(N__35744),
            .I(N__35716));
    IoSpan4Mux I__7330 (
            .O(N__35741),
            .I(N__35713));
    LocalMux I__7329 (
            .O(N__35738),
            .I(N__35710));
    IoInMux I__7328 (
            .O(N__35737),
            .I(N__35707));
    IoInMux I__7327 (
            .O(N__35736),
            .I(N__35704));
    IoInMux I__7326 (
            .O(N__35735),
            .I(N__35701));
    IoInMux I__7325 (
            .O(N__35734),
            .I(N__35698));
    IoInMux I__7324 (
            .O(N__35733),
            .I(N__35695));
    IoSpan4Mux I__7323 (
            .O(N__35726),
            .I(N__35692));
    IoInMux I__7322 (
            .O(N__35725),
            .I(N__35689));
    IoInMux I__7321 (
            .O(N__35724),
            .I(N__35686));
    IoInMux I__7320 (
            .O(N__35723),
            .I(N__35683));
    IoSpan4Mux I__7319 (
            .O(N__35716),
            .I(N__35680));
    IoSpan4Mux I__7318 (
            .O(N__35713),
            .I(N__35676));
    IoSpan4Mux I__7317 (
            .O(N__35710),
            .I(N__35671));
    LocalMux I__7316 (
            .O(N__35707),
            .I(N__35671));
    LocalMux I__7315 (
            .O(N__35704),
            .I(N__35665));
    LocalMux I__7314 (
            .O(N__35701),
            .I(N__35662));
    LocalMux I__7313 (
            .O(N__35698),
            .I(N__35657));
    LocalMux I__7312 (
            .O(N__35695),
            .I(N__35657));
    IoSpan4Mux I__7311 (
            .O(N__35692),
            .I(N__35650));
    LocalMux I__7310 (
            .O(N__35689),
            .I(N__35650));
    LocalMux I__7309 (
            .O(N__35686),
            .I(N__35650));
    LocalMux I__7308 (
            .O(N__35683),
            .I(N__35647));
    Span4Mux_s2_v I__7307 (
            .O(N__35680),
            .I(N__35644));
    IoInMux I__7306 (
            .O(N__35679),
            .I(N__35641));
    IoSpan4Mux I__7305 (
            .O(N__35676),
            .I(N__35636));
    IoSpan4Mux I__7304 (
            .O(N__35671),
            .I(N__35636));
    IoInMux I__7303 (
            .O(N__35670),
            .I(N__35633));
    IoInMux I__7302 (
            .O(N__35669),
            .I(N__35630));
    IoInMux I__7301 (
            .O(N__35668),
            .I(N__35627));
    Span4Mux_s2_v I__7300 (
            .O(N__35665),
            .I(N__35624));
    Span4Mux_s2_v I__7299 (
            .O(N__35662),
            .I(N__35621));
    IoSpan4Mux I__7298 (
            .O(N__35657),
            .I(N__35618));
    IoSpan4Mux I__7297 (
            .O(N__35650),
            .I(N__35615));
    Span12Mux_s9_h I__7296 (
            .O(N__35647),
            .I(N__35612));
    Span4Mux_v I__7295 (
            .O(N__35644),
            .I(N__35609));
    LocalMux I__7294 (
            .O(N__35641),
            .I(N__35606));
    Span4Mux_s2_h I__7293 (
            .O(N__35636),
            .I(N__35603));
    LocalMux I__7292 (
            .O(N__35633),
            .I(N__35598));
    LocalMux I__7291 (
            .O(N__35630),
            .I(N__35598));
    LocalMux I__7290 (
            .O(N__35627),
            .I(N__35595));
    Sp12to4 I__7289 (
            .O(N__35624),
            .I(N__35592));
    Sp12to4 I__7288 (
            .O(N__35621),
            .I(N__35589));
    Span4Mux_s3_h I__7287 (
            .O(N__35618),
            .I(N__35586));
    Span4Mux_s2_h I__7286 (
            .O(N__35615),
            .I(N__35583));
    Span12Mux_h I__7285 (
            .O(N__35612),
            .I(N__35580));
    Sp12to4 I__7284 (
            .O(N__35609),
            .I(N__35575));
    Span12Mux_s6_v I__7283 (
            .O(N__35606),
            .I(N__35575));
    Sp12to4 I__7282 (
            .O(N__35603),
            .I(N__35572));
    Sp12to4 I__7281 (
            .O(N__35598),
            .I(N__35569));
    Span12Mux_s9_h I__7280 (
            .O(N__35595),
            .I(N__35566));
    Span12Mux_h I__7279 (
            .O(N__35592),
            .I(N__35561));
    Span12Mux_s10_h I__7278 (
            .O(N__35589),
            .I(N__35561));
    Sp12to4 I__7277 (
            .O(N__35586),
            .I(N__35558));
    Span4Mux_h I__7276 (
            .O(N__35583),
            .I(N__35555));
    Span12Mux_v I__7275 (
            .O(N__35580),
            .I(N__35548));
    Span12Mux_v I__7274 (
            .O(N__35575),
            .I(N__35548));
    Span12Mux_s9_h I__7273 (
            .O(N__35572),
            .I(N__35548));
    Span12Mux_v I__7272 (
            .O(N__35569),
            .I(N__35545));
    Span12Mux_h I__7271 (
            .O(N__35566),
            .I(N__35538));
    Span12Mux_v I__7270 (
            .O(N__35561),
            .I(N__35538));
    Span12Mux_s10_h I__7269 (
            .O(N__35558),
            .I(N__35538));
    Span4Mux_h I__7268 (
            .O(N__35555),
            .I(N__35535));
    Odrv12 I__7267 (
            .O(N__35548),
            .I(pin_oe_22));
    Odrv12 I__7266 (
            .O(N__35545),
            .I(pin_oe_22));
    Odrv12 I__7265 (
            .O(N__35538),
            .I(pin_oe_22));
    Odrv4 I__7264 (
            .O(N__35535),
            .I(pin_oe_22));
    InMux I__7263 (
            .O(N__35526),
            .I(N__35522));
    InMux I__7262 (
            .O(N__35525),
            .I(N__35519));
    LocalMux I__7261 (
            .O(N__35522),
            .I(N__35514));
    LocalMux I__7260 (
            .O(N__35519),
            .I(N__35514));
    Span4Mux_h I__7259 (
            .O(N__35514),
            .I(N__35511));
    Odrv4 I__7258 (
            .O(N__35511),
            .I(n6158));
    CascadeMux I__7257 (
            .O(N__35508),
            .I(N__35505));
    InMux I__7256 (
            .O(N__35505),
            .I(N__35499));
    InMux I__7255 (
            .O(N__35504),
            .I(N__35494));
    InMux I__7254 (
            .O(N__35503),
            .I(N__35494));
    InMux I__7253 (
            .O(N__35502),
            .I(N__35491));
    LocalMux I__7252 (
            .O(N__35499),
            .I(N__35486));
    LocalMux I__7251 (
            .O(N__35494),
            .I(N__35486));
    LocalMux I__7250 (
            .O(N__35491),
            .I(N__35483));
    Span4Mux_h I__7249 (
            .O(N__35486),
            .I(N__35480));
    Odrv4 I__7248 (
            .O(N__35483),
            .I(n8));
    Odrv4 I__7247 (
            .O(N__35480),
            .I(n8));
    CascadeMux I__7246 (
            .O(N__35475),
            .I(n22_adj_740_cascade_));
    InMux I__7245 (
            .O(N__35472),
            .I(N__35468));
    InMux I__7244 (
            .O(N__35471),
            .I(N__35465));
    LocalMux I__7243 (
            .O(N__35468),
            .I(N__35460));
    LocalMux I__7242 (
            .O(N__35465),
            .I(N__35460));
    Span4Mux_h I__7241 (
            .O(N__35460),
            .I(N__35457));
    Odrv4 I__7240 (
            .O(N__35457),
            .I(n5907));
    InMux I__7239 (
            .O(N__35454),
            .I(N__35451));
    LocalMux I__7238 (
            .O(N__35451),
            .I(n6162));
    CascadeMux I__7237 (
            .O(N__35448),
            .I(n6162_cascade_));
    InMux I__7236 (
            .O(N__35445),
            .I(N__35442));
    LocalMux I__7235 (
            .O(N__35442),
            .I(n7278));
    InMux I__7234 (
            .O(N__35439),
            .I(N__35435));
    CascadeMux I__7233 (
            .O(N__35438),
            .I(N__35432));
    LocalMux I__7232 (
            .O(N__35435),
            .I(N__35429));
    InMux I__7231 (
            .O(N__35432),
            .I(N__35426));
    Span4Mux_v I__7230 (
            .O(N__35429),
            .I(N__35422));
    LocalMux I__7229 (
            .O(N__35426),
            .I(N__35419));
    CascadeMux I__7228 (
            .O(N__35425),
            .I(N__35416));
    Span4Mux_h I__7227 (
            .O(N__35422),
            .I(N__35411));
    Span4Mux_h I__7226 (
            .O(N__35419),
            .I(N__35411));
    InMux I__7225 (
            .O(N__35416),
            .I(N__35408));
    Odrv4 I__7224 (
            .O(N__35411),
            .I(\nx.n1704 ));
    LocalMux I__7223 (
            .O(N__35408),
            .I(\nx.n1704 ));
    InMux I__7222 (
            .O(N__35403),
            .I(N__35400));
    LocalMux I__7221 (
            .O(N__35400),
            .I(\nx.n1771 ));
    InMux I__7220 (
            .O(N__35397),
            .I(\nx.n10620 ));
    InMux I__7219 (
            .O(N__35394),
            .I(N__35387));
    InMux I__7218 (
            .O(N__35393),
            .I(N__35387));
    CascadeMux I__7217 (
            .O(N__35392),
            .I(N__35384));
    LocalMux I__7216 (
            .O(N__35387),
            .I(N__35381));
    InMux I__7215 (
            .O(N__35384),
            .I(N__35378));
    Odrv4 I__7214 (
            .O(N__35381),
            .I(\nx.n1703 ));
    LocalMux I__7213 (
            .O(N__35378),
            .I(\nx.n1703 ));
    InMux I__7212 (
            .O(N__35373),
            .I(N__35370));
    LocalMux I__7211 (
            .O(N__35370),
            .I(\nx.n1770 ));
    InMux I__7210 (
            .O(N__35367),
            .I(\nx.n10621 ));
    CascadeMux I__7209 (
            .O(N__35364),
            .I(N__35361));
    InMux I__7208 (
            .O(N__35361),
            .I(N__35358));
    LocalMux I__7207 (
            .O(N__35358),
            .I(N__35353));
    InMux I__7206 (
            .O(N__35357),
            .I(N__35348));
    InMux I__7205 (
            .O(N__35356),
            .I(N__35348));
    Odrv4 I__7204 (
            .O(N__35353),
            .I(\nx.n1702 ));
    LocalMux I__7203 (
            .O(N__35348),
            .I(\nx.n1702 ));
    CascadeMux I__7202 (
            .O(N__35343),
            .I(N__35340));
    InMux I__7201 (
            .O(N__35340),
            .I(N__35337));
    LocalMux I__7200 (
            .O(N__35337),
            .I(N__35334));
    Span4Mux_v I__7199 (
            .O(N__35334),
            .I(N__35331));
    Span4Mux_h I__7198 (
            .O(N__35331),
            .I(N__35328));
    Odrv4 I__7197 (
            .O(N__35328),
            .I(\nx.n1769 ));
    InMux I__7196 (
            .O(N__35325),
            .I(bfn_10_29_0_));
    CascadeMux I__7195 (
            .O(N__35322),
            .I(N__35319));
    InMux I__7194 (
            .O(N__35319),
            .I(N__35315));
    InMux I__7193 (
            .O(N__35318),
            .I(N__35312));
    LocalMux I__7192 (
            .O(N__35315),
            .I(N__35309));
    LocalMux I__7191 (
            .O(N__35312),
            .I(N__35306));
    Span4Mux_v I__7190 (
            .O(N__35309),
            .I(N__35301));
    Span4Mux_v I__7189 (
            .O(N__35306),
            .I(N__35301));
    Odrv4 I__7188 (
            .O(N__35301),
            .I(\nx.n1701 ));
    InMux I__7187 (
            .O(N__35298),
            .I(N__35295));
    LocalMux I__7186 (
            .O(N__35295),
            .I(N__35292));
    Span4Mux_v I__7185 (
            .O(N__35292),
            .I(N__35289));
    Odrv4 I__7184 (
            .O(N__35289),
            .I(\nx.n1768 ));
    InMux I__7183 (
            .O(N__35286),
            .I(\nx.n10623 ));
    InMux I__7182 (
            .O(N__35283),
            .I(N__35280));
    LocalMux I__7181 (
            .O(N__35280),
            .I(N__35275));
    InMux I__7180 (
            .O(N__35279),
            .I(N__35272));
    InMux I__7179 (
            .O(N__35278),
            .I(N__35269));
    Odrv4 I__7178 (
            .O(N__35275),
            .I(\nx.n1700 ));
    LocalMux I__7177 (
            .O(N__35272),
            .I(\nx.n1700 ));
    LocalMux I__7176 (
            .O(N__35269),
            .I(\nx.n1700 ));
    InMux I__7175 (
            .O(N__35262),
            .I(N__35259));
    LocalMux I__7174 (
            .O(N__35259),
            .I(N__35256));
    Odrv4 I__7173 (
            .O(N__35256),
            .I(\nx.n1767 ));
    InMux I__7172 (
            .O(N__35253),
            .I(\nx.n10624 ));
    CascadeMux I__7171 (
            .O(N__35250),
            .I(N__35246));
    CascadeMux I__7170 (
            .O(N__35249),
            .I(N__35243));
    InMux I__7169 (
            .O(N__35246),
            .I(N__35239));
    InMux I__7168 (
            .O(N__35243),
            .I(N__35234));
    InMux I__7167 (
            .O(N__35242),
            .I(N__35234));
    LocalMux I__7166 (
            .O(N__35239),
            .I(N__35231));
    LocalMux I__7165 (
            .O(N__35234),
            .I(N__35228));
    Span4Mux_h I__7164 (
            .O(N__35231),
            .I(N__35225));
    Span4Mux_h I__7163 (
            .O(N__35228),
            .I(N__35222));
    Odrv4 I__7162 (
            .O(N__35225),
            .I(\nx.n1699 ));
    Odrv4 I__7161 (
            .O(N__35222),
            .I(\nx.n1699 ));
    InMux I__7160 (
            .O(N__35217),
            .I(N__35214));
    LocalMux I__7159 (
            .O(N__35214),
            .I(N__35211));
    Odrv4 I__7158 (
            .O(N__35211),
            .I(\nx.n1766 ));
    InMux I__7157 (
            .O(N__35208),
            .I(\nx.n10625 ));
    InMux I__7156 (
            .O(N__35205),
            .I(N__35201));
    CascadeMux I__7155 (
            .O(N__35204),
            .I(N__35198));
    LocalMux I__7154 (
            .O(N__35201),
            .I(N__35195));
    InMux I__7153 (
            .O(N__35198),
            .I(N__35192));
    Span4Mux_h I__7152 (
            .O(N__35195),
            .I(N__35189));
    LocalMux I__7151 (
            .O(N__35192),
            .I(N__35186));
    Span4Mux_v I__7150 (
            .O(N__35189),
            .I(N__35182));
    Span4Mux_h I__7149 (
            .O(N__35186),
            .I(N__35179));
    InMux I__7148 (
            .O(N__35185),
            .I(N__35176));
    Odrv4 I__7147 (
            .O(N__35182),
            .I(\nx.n1698 ));
    Odrv4 I__7146 (
            .O(N__35179),
            .I(\nx.n1698 ));
    LocalMux I__7145 (
            .O(N__35176),
            .I(\nx.n1698 ));
    CascadeMux I__7144 (
            .O(N__35169),
            .I(N__35166));
    InMux I__7143 (
            .O(N__35166),
            .I(N__35163));
    LocalMux I__7142 (
            .O(N__35163),
            .I(N__35160));
    Span4Mux_v I__7141 (
            .O(N__35160),
            .I(N__35157));
    Odrv4 I__7140 (
            .O(N__35157),
            .I(\nx.n1765 ));
    InMux I__7139 (
            .O(N__35154),
            .I(\nx.n10626 ));
    InMux I__7138 (
            .O(N__35151),
            .I(N__35142));
    InMux I__7137 (
            .O(N__35150),
            .I(N__35137));
    InMux I__7136 (
            .O(N__35149),
            .I(N__35137));
    InMux I__7135 (
            .O(N__35148),
            .I(N__35134));
    InMux I__7134 (
            .O(N__35147),
            .I(N__35129));
    InMux I__7133 (
            .O(N__35146),
            .I(N__35129));
    InMux I__7132 (
            .O(N__35145),
            .I(N__35122));
    LocalMux I__7131 (
            .O(N__35142),
            .I(N__35115));
    LocalMux I__7130 (
            .O(N__35137),
            .I(N__35115));
    LocalMux I__7129 (
            .O(N__35134),
            .I(N__35115));
    LocalMux I__7128 (
            .O(N__35129),
            .I(N__35112));
    CascadeMux I__7127 (
            .O(N__35128),
            .I(N__35109));
    InMux I__7126 (
            .O(N__35127),
            .I(N__35100));
    InMux I__7125 (
            .O(N__35126),
            .I(N__35100));
    InMux I__7124 (
            .O(N__35125),
            .I(N__35100));
    LocalMux I__7123 (
            .O(N__35122),
            .I(N__35097));
    Span4Mux_h I__7122 (
            .O(N__35115),
            .I(N__35094));
    Span4Mux_h I__7121 (
            .O(N__35112),
            .I(N__35091));
    InMux I__7120 (
            .O(N__35109),
            .I(N__35084));
    InMux I__7119 (
            .O(N__35108),
            .I(N__35084));
    InMux I__7118 (
            .O(N__35107),
            .I(N__35084));
    LocalMux I__7117 (
            .O(N__35100),
            .I(\nx.n1730 ));
    Odrv4 I__7116 (
            .O(N__35097),
            .I(\nx.n1730 ));
    Odrv4 I__7115 (
            .O(N__35094),
            .I(\nx.n1730 ));
    Odrv4 I__7114 (
            .O(N__35091),
            .I(\nx.n1730 ));
    LocalMux I__7113 (
            .O(N__35084),
            .I(\nx.n1730 ));
    CascadeMux I__7112 (
            .O(N__35073),
            .I(N__35070));
    InMux I__7111 (
            .O(N__35070),
            .I(N__35067));
    LocalMux I__7110 (
            .O(N__35067),
            .I(N__35064));
    Span4Mux_h I__7109 (
            .O(N__35064),
            .I(N__35060));
    InMux I__7108 (
            .O(N__35063),
            .I(N__35057));
    Odrv4 I__7107 (
            .O(N__35060),
            .I(\nx.n1697 ));
    LocalMux I__7106 (
            .O(N__35057),
            .I(\nx.n1697 ));
    InMux I__7105 (
            .O(N__35052),
            .I(\nx.n10627 ));
    CascadeMux I__7104 (
            .O(N__35049),
            .I(N__35046));
    InMux I__7103 (
            .O(N__35046),
            .I(N__35042));
    InMux I__7102 (
            .O(N__35045),
            .I(N__35039));
    LocalMux I__7101 (
            .O(N__35042),
            .I(N__35036));
    LocalMux I__7100 (
            .O(N__35039),
            .I(\nx.n1796 ));
    Odrv4 I__7099 (
            .O(N__35036),
            .I(\nx.n1796 ));
    CascadeMux I__7098 (
            .O(N__35031),
            .I(N__35028));
    InMux I__7097 (
            .O(N__35028),
            .I(N__35025));
    LocalMux I__7096 (
            .O(N__35025),
            .I(N__35022));
    Span4Mux_v I__7095 (
            .O(N__35022),
            .I(N__35019));
    Odrv4 I__7094 (
            .O(N__35019),
            .I(\nx.n20_adj_680 ));
    InMux I__7093 (
            .O(N__35016),
            .I(N__35013));
    LocalMux I__7092 (
            .O(N__35013),
            .I(\nx.n24_adj_685 ));
    CascadeMux I__7091 (
            .O(N__35010),
            .I(\nx.n1730_cascade_ ));
    CascadeMux I__7090 (
            .O(N__35007),
            .I(N__35002));
    InMux I__7089 (
            .O(N__35006),
            .I(N__34999));
    CascadeMux I__7088 (
            .O(N__35005),
            .I(N__34996));
    InMux I__7087 (
            .O(N__35002),
            .I(N__34993));
    LocalMux I__7086 (
            .O(N__34999),
            .I(N__34990));
    InMux I__7085 (
            .O(N__34996),
            .I(N__34987));
    LocalMux I__7084 (
            .O(N__34993),
            .I(N__34982));
    Span4Mux_h I__7083 (
            .O(N__34990),
            .I(N__34982));
    LocalMux I__7082 (
            .O(N__34987),
            .I(\nx.n1802 ));
    Odrv4 I__7081 (
            .O(N__34982),
            .I(\nx.n1802 ));
    InMux I__7080 (
            .O(N__34977),
            .I(N__34972));
    InMux I__7079 (
            .O(N__34976),
            .I(N__34969));
    InMux I__7078 (
            .O(N__34975),
            .I(N__34966));
    LocalMux I__7077 (
            .O(N__34972),
            .I(N__34962));
    LocalMux I__7076 (
            .O(N__34969),
            .I(N__34959));
    LocalMux I__7075 (
            .O(N__34966),
            .I(N__34956));
    InMux I__7074 (
            .O(N__34965),
            .I(N__34953));
    Span4Mux_s3_h I__7073 (
            .O(N__34962),
            .I(N__34943));
    Span4Mux_v I__7072 (
            .O(N__34959),
            .I(N__34943));
    Span4Mux_h I__7071 (
            .O(N__34956),
            .I(N__34943));
    LocalMux I__7070 (
            .O(N__34953),
            .I(N__34943));
    InMux I__7069 (
            .O(N__34952),
            .I(N__34940));
    Span4Mux_h I__7068 (
            .O(N__34943),
            .I(N__34937));
    LocalMux I__7067 (
            .O(N__34940),
            .I(\nx.bit_ctr_18 ));
    Odrv4 I__7066 (
            .O(N__34937),
            .I(\nx.bit_ctr_18 ));
    InMux I__7065 (
            .O(N__34932),
            .I(N__34929));
    LocalMux I__7064 (
            .O(N__34929),
            .I(N__34926));
    Span4Mux_v I__7063 (
            .O(N__34926),
            .I(N__34923));
    Odrv4 I__7062 (
            .O(N__34923),
            .I(\nx.n1777 ));
    InMux I__7061 (
            .O(N__34920),
            .I(bfn_10_28_0_));
    CascadeMux I__7060 (
            .O(N__34917),
            .I(N__34913));
    CascadeMux I__7059 (
            .O(N__34916),
            .I(N__34909));
    InMux I__7058 (
            .O(N__34913),
            .I(N__34906));
    CascadeMux I__7057 (
            .O(N__34912),
            .I(N__34903));
    InMux I__7056 (
            .O(N__34909),
            .I(N__34900));
    LocalMux I__7055 (
            .O(N__34906),
            .I(N__34897));
    InMux I__7054 (
            .O(N__34903),
            .I(N__34894));
    LocalMux I__7053 (
            .O(N__34900),
            .I(\nx.n1709 ));
    Odrv12 I__7052 (
            .O(N__34897),
            .I(\nx.n1709 ));
    LocalMux I__7051 (
            .O(N__34894),
            .I(\nx.n1709 ));
    InMux I__7050 (
            .O(N__34887),
            .I(N__34884));
    LocalMux I__7049 (
            .O(N__34884),
            .I(N__34881));
    Span4Mux_v I__7048 (
            .O(N__34881),
            .I(N__34878));
    Span4Mux_h I__7047 (
            .O(N__34878),
            .I(N__34875));
    Odrv4 I__7046 (
            .O(N__34875),
            .I(\nx.n1776 ));
    InMux I__7045 (
            .O(N__34872),
            .I(\nx.n10615 ));
    CascadeMux I__7044 (
            .O(N__34869),
            .I(N__34864));
    InMux I__7043 (
            .O(N__34868),
            .I(N__34861));
    CascadeMux I__7042 (
            .O(N__34867),
            .I(N__34858));
    InMux I__7041 (
            .O(N__34864),
            .I(N__34855));
    LocalMux I__7040 (
            .O(N__34861),
            .I(N__34852));
    InMux I__7039 (
            .O(N__34858),
            .I(N__34849));
    LocalMux I__7038 (
            .O(N__34855),
            .I(N__34846));
    Span4Mux_v I__7037 (
            .O(N__34852),
            .I(N__34841));
    LocalMux I__7036 (
            .O(N__34849),
            .I(N__34841));
    Span4Mux_v I__7035 (
            .O(N__34846),
            .I(N__34838));
    Span4Mux_h I__7034 (
            .O(N__34841),
            .I(N__34835));
    Odrv4 I__7033 (
            .O(N__34838),
            .I(\nx.n1708 ));
    Odrv4 I__7032 (
            .O(N__34835),
            .I(\nx.n1708 ));
    InMux I__7031 (
            .O(N__34830),
            .I(N__34827));
    LocalMux I__7030 (
            .O(N__34827),
            .I(N__34824));
    Odrv4 I__7029 (
            .O(N__34824),
            .I(\nx.n1775 ));
    InMux I__7028 (
            .O(N__34821),
            .I(\nx.n10616 ));
    CascadeMux I__7027 (
            .O(N__34818),
            .I(N__34815));
    InMux I__7026 (
            .O(N__34815),
            .I(N__34811));
    InMux I__7025 (
            .O(N__34814),
            .I(N__34808));
    LocalMux I__7024 (
            .O(N__34811),
            .I(\nx.n1707 ));
    LocalMux I__7023 (
            .O(N__34808),
            .I(\nx.n1707 ));
    InMux I__7022 (
            .O(N__34803),
            .I(N__34800));
    LocalMux I__7021 (
            .O(N__34800),
            .I(\nx.n1774 ));
    InMux I__7020 (
            .O(N__34797),
            .I(\nx.n10617 ));
    CascadeMux I__7019 (
            .O(N__34794),
            .I(N__34791));
    InMux I__7018 (
            .O(N__34791),
            .I(N__34788));
    LocalMux I__7017 (
            .O(N__34788),
            .I(N__34784));
    InMux I__7016 (
            .O(N__34787),
            .I(N__34781));
    Span4Mux_v I__7015 (
            .O(N__34784),
            .I(N__34775));
    LocalMux I__7014 (
            .O(N__34781),
            .I(N__34775));
    InMux I__7013 (
            .O(N__34780),
            .I(N__34772));
    Span4Mux_h I__7012 (
            .O(N__34775),
            .I(N__34769));
    LocalMux I__7011 (
            .O(N__34772),
            .I(\nx.n1706 ));
    Odrv4 I__7010 (
            .O(N__34769),
            .I(\nx.n1706 ));
    InMux I__7009 (
            .O(N__34764),
            .I(N__34761));
    LocalMux I__7008 (
            .O(N__34761),
            .I(N__34758));
    Span4Mux_h I__7007 (
            .O(N__34758),
            .I(N__34755));
    Odrv4 I__7006 (
            .O(N__34755),
            .I(\nx.n1773 ));
    InMux I__7005 (
            .O(N__34752),
            .I(\nx.n10618 ));
    CascadeMux I__7004 (
            .O(N__34749),
            .I(N__34746));
    InMux I__7003 (
            .O(N__34746),
            .I(N__34743));
    LocalMux I__7002 (
            .O(N__34743),
            .I(N__34738));
    CascadeMux I__7001 (
            .O(N__34742),
            .I(N__34735));
    InMux I__7000 (
            .O(N__34741),
            .I(N__34732));
    Span4Mux_h I__6999 (
            .O(N__34738),
            .I(N__34729));
    InMux I__6998 (
            .O(N__34735),
            .I(N__34726));
    LocalMux I__6997 (
            .O(N__34732),
            .I(N__34723));
    Odrv4 I__6996 (
            .O(N__34729),
            .I(\nx.n1705 ));
    LocalMux I__6995 (
            .O(N__34726),
            .I(\nx.n1705 ));
    Odrv4 I__6994 (
            .O(N__34723),
            .I(\nx.n1705 ));
    InMux I__6993 (
            .O(N__34716),
            .I(N__34713));
    LocalMux I__6992 (
            .O(N__34713),
            .I(N__34710));
    Span4Mux_h I__6991 (
            .O(N__34710),
            .I(N__34707));
    Odrv4 I__6990 (
            .O(N__34707),
            .I(\nx.n1772 ));
    InMux I__6989 (
            .O(N__34704),
            .I(\nx.n10619 ));
    CascadeMux I__6988 (
            .O(N__34701),
            .I(\nx.n2097_cascade_ ));
    InMux I__6987 (
            .O(N__34698),
            .I(N__34695));
    LocalMux I__6986 (
            .O(N__34695),
            .I(\nx.n27_adj_671 ));
    CascadeMux I__6985 (
            .O(N__34692),
            .I(N__34688));
    CascadeMux I__6984 (
            .O(N__34691),
            .I(N__34684));
    InMux I__6983 (
            .O(N__34688),
            .I(N__34681));
    InMux I__6982 (
            .O(N__34687),
            .I(N__34678));
    InMux I__6981 (
            .O(N__34684),
            .I(N__34675));
    LocalMux I__6980 (
            .O(N__34681),
            .I(N__34672));
    LocalMux I__6979 (
            .O(N__34678),
            .I(N__34667));
    LocalMux I__6978 (
            .O(N__34675),
            .I(N__34667));
    Span4Mux_h I__6977 (
            .O(N__34672),
            .I(N__34662));
    Span4Mux_v I__6976 (
            .O(N__34667),
            .I(N__34662));
    Odrv4 I__6975 (
            .O(N__34662),
            .I(\nx.n2007 ));
    InMux I__6974 (
            .O(N__34659),
            .I(N__34655));
    CascadeMux I__6973 (
            .O(N__34658),
            .I(N__34652));
    LocalMux I__6972 (
            .O(N__34655),
            .I(N__34649));
    InMux I__6971 (
            .O(N__34652),
            .I(N__34646));
    Span4Mux_v I__6970 (
            .O(N__34649),
            .I(N__34640));
    LocalMux I__6969 (
            .O(N__34646),
            .I(N__34640));
    InMux I__6968 (
            .O(N__34645),
            .I(N__34637));
    Span4Mux_h I__6967 (
            .O(N__34640),
            .I(N__34634));
    LocalMux I__6966 (
            .O(N__34637),
            .I(N__34631));
    Odrv4 I__6965 (
            .O(N__34634),
            .I(\nx.n2002 ));
    Odrv12 I__6964 (
            .O(N__34631),
            .I(\nx.n2002 ));
    InMux I__6963 (
            .O(N__34626),
            .I(N__34623));
    LocalMux I__6962 (
            .O(N__34623),
            .I(N__34620));
    Odrv4 I__6961 (
            .O(N__34620),
            .I(\nx.n22_adj_662 ));
    CascadeMux I__6960 (
            .O(N__34617),
            .I(N__34614));
    InMux I__6959 (
            .O(N__34614),
            .I(N__34609));
    InMux I__6958 (
            .O(N__34613),
            .I(N__34606));
    InMux I__6957 (
            .O(N__34612),
            .I(N__34603));
    LocalMux I__6956 (
            .O(N__34609),
            .I(N__34598));
    LocalMux I__6955 (
            .O(N__34606),
            .I(N__34598));
    LocalMux I__6954 (
            .O(N__34603),
            .I(\nx.n1803 ));
    Odrv12 I__6953 (
            .O(N__34598),
            .I(\nx.n1803 ));
    CascadeMux I__6952 (
            .O(N__34593),
            .I(\nx.n22_adj_673_cascade_ ));
    InMux I__6951 (
            .O(N__34590),
            .I(N__34587));
    LocalMux I__6950 (
            .O(N__34587),
            .I(N__34584));
    Span4Mux_h I__6949 (
            .O(N__34584),
            .I(N__34581));
    Odrv4 I__6948 (
            .O(N__34581),
            .I(\nx.n16_adj_672 ));
    InMux I__6947 (
            .O(N__34578),
            .I(N__34574));
    CascadeMux I__6946 (
            .O(N__34577),
            .I(N__34571));
    LocalMux I__6945 (
            .O(N__34574),
            .I(N__34567));
    InMux I__6944 (
            .O(N__34571),
            .I(N__34564));
    InMux I__6943 (
            .O(N__34570),
            .I(N__34561));
    Odrv4 I__6942 (
            .O(N__34567),
            .I(\nx.n1798 ));
    LocalMux I__6941 (
            .O(N__34564),
            .I(\nx.n1798 ));
    LocalMux I__6940 (
            .O(N__34561),
            .I(\nx.n1798 ));
    CascadeMux I__6939 (
            .O(N__34554),
            .I(N__34551));
    InMux I__6938 (
            .O(N__34551),
            .I(N__34547));
    InMux I__6937 (
            .O(N__34550),
            .I(N__34544));
    LocalMux I__6936 (
            .O(N__34547),
            .I(N__34541));
    LocalMux I__6935 (
            .O(N__34544),
            .I(N__34536));
    Span4Mux_h I__6934 (
            .O(N__34541),
            .I(N__34536));
    Odrv4 I__6933 (
            .O(N__34536),
            .I(\nx.n1608 ));
    CascadeMux I__6932 (
            .O(N__34533),
            .I(N__34530));
    InMux I__6931 (
            .O(N__34530),
            .I(N__34527));
    LocalMux I__6930 (
            .O(N__34527),
            .I(N__34524));
    Span4Mux_h I__6929 (
            .O(N__34524),
            .I(N__34521));
    Odrv4 I__6928 (
            .O(N__34521),
            .I(\nx.n1675 ));
    InMux I__6927 (
            .O(N__34518),
            .I(N__34512));
    CascadeMux I__6926 (
            .O(N__34517),
            .I(N__34508));
    InMux I__6925 (
            .O(N__34516),
            .I(N__34505));
    CascadeMux I__6924 (
            .O(N__34515),
            .I(N__34501));
    LocalMux I__6923 (
            .O(N__34512),
            .I(N__34496));
    InMux I__6922 (
            .O(N__34511),
            .I(N__34491));
    InMux I__6921 (
            .O(N__34508),
            .I(N__34491));
    LocalMux I__6920 (
            .O(N__34505),
            .I(N__34488));
    InMux I__6919 (
            .O(N__34504),
            .I(N__34483));
    InMux I__6918 (
            .O(N__34501),
            .I(N__34483));
    CascadeMux I__6917 (
            .O(N__34500),
            .I(N__34477));
    InMux I__6916 (
            .O(N__34499),
            .I(N__34473));
    Span4Mux_v I__6915 (
            .O(N__34496),
            .I(N__34468));
    LocalMux I__6914 (
            .O(N__34491),
            .I(N__34468));
    Span4Mux_h I__6913 (
            .O(N__34488),
            .I(N__34463));
    LocalMux I__6912 (
            .O(N__34483),
            .I(N__34463));
    InMux I__6911 (
            .O(N__34482),
            .I(N__34458));
    InMux I__6910 (
            .O(N__34481),
            .I(N__34458));
    InMux I__6909 (
            .O(N__34480),
            .I(N__34455));
    InMux I__6908 (
            .O(N__34477),
            .I(N__34450));
    InMux I__6907 (
            .O(N__34476),
            .I(N__34450));
    LocalMux I__6906 (
            .O(N__34473),
            .I(\nx.n1631 ));
    Odrv4 I__6905 (
            .O(N__34468),
            .I(\nx.n1631 ));
    Odrv4 I__6904 (
            .O(N__34463),
            .I(\nx.n1631 ));
    LocalMux I__6903 (
            .O(N__34458),
            .I(\nx.n1631 ));
    LocalMux I__6902 (
            .O(N__34455),
            .I(\nx.n1631 ));
    LocalMux I__6901 (
            .O(N__34450),
            .I(\nx.n1631 ));
    CascadeMux I__6900 (
            .O(N__34437),
            .I(\nx.n1707_cascade_ ));
    InMux I__6899 (
            .O(N__34434),
            .I(N__34429));
    InMux I__6898 (
            .O(N__34433),
            .I(N__34426));
    CascadeMux I__6897 (
            .O(N__34432),
            .I(N__34423));
    LocalMux I__6896 (
            .O(N__34429),
            .I(N__34420));
    LocalMux I__6895 (
            .O(N__34426),
            .I(N__34417));
    InMux I__6894 (
            .O(N__34423),
            .I(N__34414));
    Span4Mux_v I__6893 (
            .O(N__34420),
            .I(N__34411));
    Odrv4 I__6892 (
            .O(N__34417),
            .I(\nx.n1806 ));
    LocalMux I__6891 (
            .O(N__34414),
            .I(\nx.n1806 ));
    Odrv4 I__6890 (
            .O(N__34411),
            .I(\nx.n1806 ));
    InMux I__6889 (
            .O(N__34404),
            .I(N__34401));
    LocalMux I__6888 (
            .O(N__34401),
            .I(\nx.n2074 ));
    InMux I__6887 (
            .O(N__34398),
            .I(N__34395));
    LocalMux I__6886 (
            .O(N__34395),
            .I(\nx.n2064 ));
    CascadeMux I__6885 (
            .O(N__34392),
            .I(N__34389));
    InMux I__6884 (
            .O(N__34389),
            .I(N__34385));
    CascadeMux I__6883 (
            .O(N__34388),
            .I(N__34382));
    LocalMux I__6882 (
            .O(N__34385),
            .I(N__34379));
    InMux I__6881 (
            .O(N__34382),
            .I(N__34376));
    Span4Mux_v I__6880 (
            .O(N__34379),
            .I(N__34370));
    LocalMux I__6879 (
            .O(N__34376),
            .I(N__34370));
    InMux I__6878 (
            .O(N__34375),
            .I(N__34367));
    Span4Mux_h I__6877 (
            .O(N__34370),
            .I(N__34364));
    LocalMux I__6876 (
            .O(N__34367),
            .I(N__34361));
    Odrv4 I__6875 (
            .O(N__34364),
            .I(\nx.n1997 ));
    Odrv12 I__6874 (
            .O(N__34361),
            .I(\nx.n1997 ));
    InMux I__6873 (
            .O(N__34356),
            .I(N__34353));
    LocalMux I__6872 (
            .O(N__34353),
            .I(\nx.n2062 ));
    CascadeMux I__6871 (
            .O(N__34350),
            .I(N__34347));
    InMux I__6870 (
            .O(N__34347),
            .I(N__34343));
    CascadeMux I__6869 (
            .O(N__34346),
            .I(N__34340));
    LocalMux I__6868 (
            .O(N__34343),
            .I(N__34336));
    InMux I__6867 (
            .O(N__34340),
            .I(N__34333));
    CascadeMux I__6866 (
            .O(N__34339),
            .I(N__34330));
    Span4Mux_v I__6865 (
            .O(N__34336),
            .I(N__34325));
    LocalMux I__6864 (
            .O(N__34333),
            .I(N__34325));
    InMux I__6863 (
            .O(N__34330),
            .I(N__34322));
    Span4Mux_h I__6862 (
            .O(N__34325),
            .I(N__34319));
    LocalMux I__6861 (
            .O(N__34322),
            .I(N__34316));
    Odrv4 I__6860 (
            .O(N__34319),
            .I(\nx.n1995 ));
    Odrv12 I__6859 (
            .O(N__34316),
            .I(\nx.n1995 ));
    InMux I__6858 (
            .O(N__34311),
            .I(N__34308));
    LocalMux I__6857 (
            .O(N__34308),
            .I(N__34305));
    Odrv4 I__6856 (
            .O(N__34305),
            .I(\nx.n26_adj_667 ));
    CascadeMux I__6855 (
            .O(N__34302),
            .I(\nx.n30_adj_668_cascade_ ));
    InMux I__6854 (
            .O(N__34299),
            .I(N__34296));
    LocalMux I__6853 (
            .O(N__34296),
            .I(N__34293));
    Odrv4 I__6852 (
            .O(N__34293),
            .I(\nx.n28_adj_669 ));
    CascadeMux I__6851 (
            .O(N__34290),
            .I(N__34286));
    InMux I__6850 (
            .O(N__34289),
            .I(N__34283));
    InMux I__6849 (
            .O(N__34286),
            .I(N__34280));
    LocalMux I__6848 (
            .O(N__34283),
            .I(N__34277));
    LocalMux I__6847 (
            .O(N__34280),
            .I(N__34273));
    Span4Mux_v I__6846 (
            .O(N__34277),
            .I(N__34270));
    InMux I__6845 (
            .O(N__34276),
            .I(N__34267));
    Span4Mux_h I__6844 (
            .O(N__34273),
            .I(N__34264));
    Odrv4 I__6843 (
            .O(N__34270),
            .I(\nx.n2008 ));
    LocalMux I__6842 (
            .O(N__34267),
            .I(\nx.n2008 ));
    Odrv4 I__6841 (
            .O(N__34264),
            .I(\nx.n2008 ));
    CascadeMux I__6840 (
            .O(N__34257),
            .I(N__34254));
    InMux I__6839 (
            .O(N__34254),
            .I(N__34251));
    LocalMux I__6838 (
            .O(N__34251),
            .I(\nx.n2075 ));
    CascadeMux I__6837 (
            .O(N__34248),
            .I(\nx.n2107_cascade_ ));
    InMux I__6836 (
            .O(N__34245),
            .I(N__34242));
    LocalMux I__6835 (
            .O(N__34242),
            .I(\nx.n29_adj_670 ));
    InMux I__6834 (
            .O(N__34239),
            .I(N__34236));
    LocalMux I__6833 (
            .O(N__34236),
            .I(\nx.n2065 ));
    InMux I__6832 (
            .O(N__34233),
            .I(N__34228));
    CascadeMux I__6831 (
            .O(N__34232),
            .I(N__34225));
    CascadeMux I__6830 (
            .O(N__34231),
            .I(N__34222));
    LocalMux I__6829 (
            .O(N__34228),
            .I(N__34219));
    InMux I__6828 (
            .O(N__34225),
            .I(N__34216));
    InMux I__6827 (
            .O(N__34222),
            .I(N__34213));
    Span4Mux_h I__6826 (
            .O(N__34219),
            .I(N__34210));
    LocalMux I__6825 (
            .O(N__34216),
            .I(N__34205));
    LocalMux I__6824 (
            .O(N__34213),
            .I(N__34205));
    Span4Mux_v I__6823 (
            .O(N__34210),
            .I(N__34200));
    Span4Mux_v I__6822 (
            .O(N__34205),
            .I(N__34200));
    Odrv4 I__6821 (
            .O(N__34200),
            .I(\nx.n1998 ));
    CascadeMux I__6820 (
            .O(N__34197),
            .I(N__34186));
    CascadeMux I__6819 (
            .O(N__34196),
            .I(N__34180));
    CascadeMux I__6818 (
            .O(N__34195),
            .I(N__34177));
    InMux I__6817 (
            .O(N__34194),
            .I(N__34172));
    InMux I__6816 (
            .O(N__34193),
            .I(N__34172));
    InMux I__6815 (
            .O(N__34192),
            .I(N__34169));
    CascadeMux I__6814 (
            .O(N__34191),
            .I(N__34165));
    CascadeMux I__6813 (
            .O(N__34190),
            .I(N__34161));
    InMux I__6812 (
            .O(N__34189),
            .I(N__34156));
    InMux I__6811 (
            .O(N__34186),
            .I(N__34143));
    InMux I__6810 (
            .O(N__34185),
            .I(N__34143));
    InMux I__6809 (
            .O(N__34184),
            .I(N__34143));
    InMux I__6808 (
            .O(N__34183),
            .I(N__34143));
    InMux I__6807 (
            .O(N__34180),
            .I(N__34143));
    InMux I__6806 (
            .O(N__34177),
            .I(N__34143));
    LocalMux I__6805 (
            .O(N__34172),
            .I(N__34138));
    LocalMux I__6804 (
            .O(N__34169),
            .I(N__34138));
    InMux I__6803 (
            .O(N__34168),
            .I(N__34131));
    InMux I__6802 (
            .O(N__34165),
            .I(N__34131));
    InMux I__6801 (
            .O(N__34164),
            .I(N__34131));
    InMux I__6800 (
            .O(N__34161),
            .I(N__34124));
    InMux I__6799 (
            .O(N__34160),
            .I(N__34124));
    InMux I__6798 (
            .O(N__34159),
            .I(N__34124));
    LocalMux I__6797 (
            .O(N__34156),
            .I(\nx.n2027 ));
    LocalMux I__6796 (
            .O(N__34143),
            .I(\nx.n2027 ));
    Odrv4 I__6795 (
            .O(N__34138),
            .I(\nx.n2027 ));
    LocalMux I__6794 (
            .O(N__34131),
            .I(\nx.n2027 ));
    LocalMux I__6793 (
            .O(N__34124),
            .I(\nx.n2027 ));
    CascadeMux I__6792 (
            .O(N__34113),
            .I(\nx.n2394_cascade_ ));
    InMux I__6791 (
            .O(N__34110),
            .I(N__34107));
    LocalMux I__6790 (
            .O(N__34107),
            .I(\nx.n2077 ));
    InMux I__6789 (
            .O(N__34104),
            .I(N__34101));
    LocalMux I__6788 (
            .O(N__34101),
            .I(\nx.n2070 ));
    CascadeMux I__6787 (
            .O(N__34098),
            .I(N__34095));
    InMux I__6786 (
            .O(N__34095),
            .I(N__34092));
    LocalMux I__6785 (
            .O(N__34092),
            .I(\nx.n2069 ));
    InMux I__6784 (
            .O(N__34089),
            .I(N__34086));
    LocalMux I__6783 (
            .O(N__34086),
            .I(\nx.n2076 ));
    InMux I__6782 (
            .O(N__34083),
            .I(N__34080));
    LocalMux I__6781 (
            .O(N__34080),
            .I(N__34077));
    Span4Mux_v I__6780 (
            .O(N__34077),
            .I(N__34071));
    InMux I__6779 (
            .O(N__34076),
            .I(N__34068));
    InMux I__6778 (
            .O(N__34075),
            .I(N__34065));
    InMux I__6777 (
            .O(N__34074),
            .I(N__34061));
    Sp12to4 I__6776 (
            .O(N__34071),
            .I(N__34054));
    LocalMux I__6775 (
            .O(N__34068),
            .I(N__34054));
    LocalMux I__6774 (
            .O(N__34065),
            .I(N__34054));
    InMux I__6773 (
            .O(N__34064),
            .I(N__34051));
    LocalMux I__6772 (
            .O(N__34061),
            .I(N__34046));
    Span12Mux_h I__6771 (
            .O(N__34054),
            .I(N__34046));
    LocalMux I__6770 (
            .O(N__34051),
            .I(\nx.bit_ctr_15 ));
    Odrv12 I__6769 (
            .O(N__34046),
            .I(\nx.bit_ctr_15 ));
    CascadeMux I__6768 (
            .O(N__34041),
            .I(N__34036));
    InMux I__6767 (
            .O(N__34040),
            .I(N__34031));
    InMux I__6766 (
            .O(N__34039),
            .I(N__34031));
    InMux I__6765 (
            .O(N__34036),
            .I(N__34028));
    LocalMux I__6764 (
            .O(N__34031),
            .I(N__34023));
    LocalMux I__6763 (
            .O(N__34028),
            .I(N__34023));
    Span4Mux_h I__6762 (
            .O(N__34023),
            .I(N__34020));
    Odrv4 I__6761 (
            .O(N__34020),
            .I(\nx.n2003 ));
    CascadeMux I__6760 (
            .O(N__34017),
            .I(N__34012));
    CascadeMux I__6759 (
            .O(N__34016),
            .I(N__34009));
    InMux I__6758 (
            .O(N__34015),
            .I(N__34004));
    InMux I__6757 (
            .O(N__34012),
            .I(N__34004));
    InMux I__6756 (
            .O(N__34009),
            .I(N__34001));
    LocalMux I__6755 (
            .O(N__34004),
            .I(N__33996));
    LocalMux I__6754 (
            .O(N__34001),
            .I(N__33996));
    Span4Mux_h I__6753 (
            .O(N__33996),
            .I(N__33993));
    Odrv4 I__6752 (
            .O(N__33993),
            .I(\nx.n2009 ));
    InMux I__6751 (
            .O(N__33990),
            .I(N__33987));
    LocalMux I__6750 (
            .O(N__33987),
            .I(\nx.n27_adj_665 ));
    InMux I__6749 (
            .O(N__33984),
            .I(N__33981));
    LocalMux I__6748 (
            .O(N__33981),
            .I(\nx.n36 ));
    InMux I__6747 (
            .O(N__33978),
            .I(N__33975));
    LocalMux I__6746 (
            .O(N__33975),
            .I(N__33972));
    Span4Mux_h I__6745 (
            .O(N__33972),
            .I(N__33969));
    Odrv4 I__6744 (
            .O(N__33969),
            .I(\nx.n41 ));
    InMux I__6743 (
            .O(N__33966),
            .I(N__33963));
    LocalMux I__6742 (
            .O(N__33963),
            .I(\nx.n2656 ));
    CascadeMux I__6741 (
            .O(N__33960),
            .I(\nx.n31_adj_655_cascade_ ));
    InMux I__6740 (
            .O(N__33957),
            .I(N__33954));
    LocalMux I__6739 (
            .O(N__33954),
            .I(N__33951));
    Span4Mux_h I__6738 (
            .O(N__33951),
            .I(N__33948));
    Span4Mux_v I__6737 (
            .O(N__33948),
            .I(N__33945));
    Odrv4 I__6736 (
            .O(N__33945),
            .I(\nx.n24_adj_654 ));
    CascadeMux I__6735 (
            .O(N__33942),
            .I(\nx.n36_adj_656_cascade_ ));
    InMux I__6734 (
            .O(N__33939),
            .I(N__33936));
    LocalMux I__6733 (
            .O(N__33936),
            .I(N__33933));
    Span4Mux_h I__6732 (
            .O(N__33933),
            .I(N__33930));
    Odrv4 I__6731 (
            .O(N__33930),
            .I(\nx.n33_adj_659 ));
    CascadeMux I__6730 (
            .O(N__33927),
            .I(\nx.n2423_cascade_ ));
    CascadeMux I__6729 (
            .O(N__33924),
            .I(\nx.n2491_cascade_ ));
    InMux I__6728 (
            .O(N__33921),
            .I(\nx.n10788 ));
    InMux I__6727 (
            .O(N__33918),
            .I(\nx.n10789 ));
    CascadeMux I__6726 (
            .O(N__33915),
            .I(N__33912));
    InMux I__6725 (
            .O(N__33912),
            .I(N__33909));
    LocalMux I__6724 (
            .O(N__33909),
            .I(\nx.n2660 ));
    CascadeMux I__6723 (
            .O(N__33906),
            .I(N__33903));
    InMux I__6722 (
            .O(N__33903),
            .I(N__33899));
    CascadeMux I__6721 (
            .O(N__33902),
            .I(N__33896));
    LocalMux I__6720 (
            .O(N__33899),
            .I(N__33893));
    InMux I__6719 (
            .O(N__33896),
            .I(N__33890));
    Span4Mux_v I__6718 (
            .O(N__33893),
            .I(N__33885));
    LocalMux I__6717 (
            .O(N__33890),
            .I(N__33885));
    Span4Mux_h I__6716 (
            .O(N__33885),
            .I(N__33881));
    InMux I__6715 (
            .O(N__33884),
            .I(N__33878));
    Odrv4 I__6714 (
            .O(N__33881),
            .I(\nx.n2692 ));
    LocalMux I__6713 (
            .O(N__33878),
            .I(\nx.n2692 ));
    CascadeMux I__6712 (
            .O(N__33873),
            .I(\nx.n34_adj_603_cascade_ ));
    CascadeMux I__6711 (
            .O(N__33870),
            .I(\nx.n39_cascade_ ));
    CascadeMux I__6710 (
            .O(N__33867),
            .I(\nx.n2621_cascade_ ));
    InMux I__6709 (
            .O(N__33864),
            .I(N__33861));
    LocalMux I__6708 (
            .O(N__33861),
            .I(\nx.n2661 ));
    CascadeMux I__6707 (
            .O(N__33858),
            .I(N__33854));
    InMux I__6706 (
            .O(N__33857),
            .I(N__33850));
    InMux I__6705 (
            .O(N__33854),
            .I(N__33847));
    InMux I__6704 (
            .O(N__33853),
            .I(N__33844));
    LocalMux I__6703 (
            .O(N__33850),
            .I(N__33841));
    LocalMux I__6702 (
            .O(N__33847),
            .I(N__33838));
    LocalMux I__6701 (
            .O(N__33844),
            .I(N__33835));
    Span4Mux_v I__6700 (
            .O(N__33841),
            .I(N__33830));
    Span4Mux_v I__6699 (
            .O(N__33838),
            .I(N__33830));
    Span4Mux_h I__6698 (
            .O(N__33835),
            .I(N__33827));
    Odrv4 I__6697 (
            .O(N__33830),
            .I(\nx.n2693 ));
    Odrv4 I__6696 (
            .O(N__33827),
            .I(\nx.n2693 ));
    InMux I__6695 (
            .O(N__33822),
            .I(N__33819));
    LocalMux I__6694 (
            .O(N__33819),
            .I(N__33816));
    Odrv4 I__6693 (
            .O(N__33816),
            .I(\nx.n2667 ));
    CascadeMux I__6692 (
            .O(N__33813),
            .I(N__33810));
    InMux I__6691 (
            .O(N__33810),
            .I(N__33806));
    CascadeMux I__6690 (
            .O(N__33809),
            .I(N__33803));
    LocalMux I__6689 (
            .O(N__33806),
            .I(N__33800));
    InMux I__6688 (
            .O(N__33803),
            .I(N__33797));
    Span4Mux_h I__6687 (
            .O(N__33800),
            .I(N__33792));
    LocalMux I__6686 (
            .O(N__33797),
            .I(N__33792));
    Odrv4 I__6685 (
            .O(N__33792),
            .I(\nx.n2699 ));
    CascadeMux I__6684 (
            .O(N__33789),
            .I(N__33786));
    InMux I__6683 (
            .O(N__33786),
            .I(N__33783));
    LocalMux I__6682 (
            .O(N__33783),
            .I(N__33780));
    Span4Mux_h I__6681 (
            .O(N__33780),
            .I(N__33776));
    InMux I__6680 (
            .O(N__33779),
            .I(N__33773));
    Odrv4 I__6679 (
            .O(N__33776),
            .I(\nx.n2687 ));
    LocalMux I__6678 (
            .O(N__33773),
            .I(\nx.n2687 ));
    CascadeMux I__6677 (
            .O(N__33768),
            .I(\nx.n2699_cascade_ ));
    CascadeMux I__6676 (
            .O(N__33765),
            .I(N__33762));
    InMux I__6675 (
            .O(N__33762),
            .I(N__33759));
    LocalMux I__6674 (
            .O(N__33759),
            .I(\nx.n2665 ));
    InMux I__6673 (
            .O(N__33756),
            .I(\nx.n10779 ));
    InMux I__6672 (
            .O(N__33753),
            .I(N__33750));
    LocalMux I__6671 (
            .O(N__33750),
            .I(N__33747));
    Span4Mux_v I__6670 (
            .O(N__33747),
            .I(N__33744));
    Span4Mux_h I__6669 (
            .O(N__33744),
            .I(N__33741));
    Odrv4 I__6668 (
            .O(N__33741),
            .I(\nx.n2664 ));
    InMux I__6667 (
            .O(N__33738),
            .I(\nx.n10780 ));
    CascadeMux I__6666 (
            .O(N__33735),
            .I(N__33732));
    InMux I__6665 (
            .O(N__33732),
            .I(N__33729));
    LocalMux I__6664 (
            .O(N__33729),
            .I(\nx.n2663 ));
    InMux I__6663 (
            .O(N__33726),
            .I(\nx.n10781 ));
    CascadeMux I__6662 (
            .O(N__33723),
            .I(N__33720));
    InMux I__6661 (
            .O(N__33720),
            .I(N__33716));
    InMux I__6660 (
            .O(N__33719),
            .I(N__33713));
    LocalMux I__6659 (
            .O(N__33716),
            .I(N__33710));
    LocalMux I__6658 (
            .O(N__33713),
            .I(N__33707));
    Span4Mux_h I__6657 (
            .O(N__33710),
            .I(N__33704));
    Odrv4 I__6656 (
            .O(N__33707),
            .I(\nx.n2595 ));
    Odrv4 I__6655 (
            .O(N__33704),
            .I(\nx.n2595 ));
    InMux I__6654 (
            .O(N__33699),
            .I(N__33696));
    LocalMux I__6653 (
            .O(N__33696),
            .I(\nx.n2662 ));
    InMux I__6652 (
            .O(N__33693),
            .I(\nx.n10782 ));
    InMux I__6651 (
            .O(N__33690),
            .I(bfn_10_19_0_));
    InMux I__6650 (
            .O(N__33687),
            .I(\nx.n10784 ));
    CascadeMux I__6649 (
            .O(N__33684),
            .I(N__33681));
    InMux I__6648 (
            .O(N__33681),
            .I(N__33677));
    InMux I__6647 (
            .O(N__33680),
            .I(N__33674));
    LocalMux I__6646 (
            .O(N__33677),
            .I(\nx.n2592 ));
    LocalMux I__6645 (
            .O(N__33674),
            .I(\nx.n2592 ));
    InMux I__6644 (
            .O(N__33669),
            .I(N__33666));
    LocalMux I__6643 (
            .O(N__33666),
            .I(\nx.n2659 ));
    InMux I__6642 (
            .O(N__33663),
            .I(\nx.n10785 ));
    InMux I__6641 (
            .O(N__33660),
            .I(N__33657));
    LocalMux I__6640 (
            .O(N__33657),
            .I(\nx.n2658 ));
    InMux I__6639 (
            .O(N__33654),
            .I(\nx.n10786 ));
    InMux I__6638 (
            .O(N__33651),
            .I(N__33648));
    LocalMux I__6637 (
            .O(N__33648),
            .I(\nx.n2657 ));
    InMux I__6636 (
            .O(N__33645),
            .I(\nx.n10787 ));
    InMux I__6635 (
            .O(N__33642),
            .I(\nx.n10771 ));
    InMux I__6634 (
            .O(N__33639),
            .I(N__33636));
    LocalMux I__6633 (
            .O(N__33636),
            .I(N__33633));
    Odrv4 I__6632 (
            .O(N__33633),
            .I(\nx.n2672 ));
    InMux I__6631 (
            .O(N__33630),
            .I(\nx.n10772 ));
    InMux I__6630 (
            .O(N__33627),
            .I(N__33624));
    LocalMux I__6629 (
            .O(N__33624),
            .I(N__33621));
    Odrv4 I__6628 (
            .O(N__33621),
            .I(\nx.n2671 ));
    InMux I__6627 (
            .O(N__33618),
            .I(\nx.n10773 ));
    CascadeMux I__6626 (
            .O(N__33615),
            .I(N__33612));
    InMux I__6625 (
            .O(N__33612),
            .I(N__33609));
    LocalMux I__6624 (
            .O(N__33609),
            .I(N__33606));
    Odrv4 I__6623 (
            .O(N__33606),
            .I(\nx.n2670 ));
    InMux I__6622 (
            .O(N__33603),
            .I(\nx.n10774 ));
    InMux I__6621 (
            .O(N__33600),
            .I(N__33597));
    LocalMux I__6620 (
            .O(N__33597),
            .I(N__33594));
    Odrv4 I__6619 (
            .O(N__33594),
            .I(\nx.n2669 ));
    InMux I__6618 (
            .O(N__33591),
            .I(bfn_10_18_0_));
    CascadeMux I__6617 (
            .O(N__33588),
            .I(N__33585));
    InMux I__6616 (
            .O(N__33585),
            .I(N__33582));
    LocalMux I__6615 (
            .O(N__33582),
            .I(N__33579));
    Odrv12 I__6614 (
            .O(N__33579),
            .I(\nx.n2668 ));
    InMux I__6613 (
            .O(N__33576),
            .I(\nx.n10776 ));
    InMux I__6612 (
            .O(N__33573),
            .I(\nx.n10777 ));
    InMux I__6611 (
            .O(N__33570),
            .I(N__33567));
    LocalMux I__6610 (
            .O(N__33567),
            .I(\nx.n2666 ));
    InMux I__6609 (
            .O(N__33564),
            .I(\nx.n10778 ));
    IoInMux I__6608 (
            .O(N__33561),
            .I(N__33558));
    LocalMux I__6607 (
            .O(N__33558),
            .I(N__33555));
    Span4Mux_s2_h I__6606 (
            .O(N__33555),
            .I(N__33552));
    Span4Mux_v I__6605 (
            .O(N__33552),
            .I(N__33549));
    Sp12to4 I__6604 (
            .O(N__33549),
            .I(N__33545));
    CascadeMux I__6603 (
            .O(N__33548),
            .I(N__33542));
    Span12Mux_s9_h I__6602 (
            .O(N__33545),
            .I(N__33538));
    InMux I__6601 (
            .O(N__33542),
            .I(N__33535));
    InMux I__6600 (
            .O(N__33541),
            .I(N__33532));
    Odrv12 I__6599 (
            .O(N__33538),
            .I(pin_out_6));
    LocalMux I__6598 (
            .O(N__33535),
            .I(pin_out_6));
    LocalMux I__6597 (
            .O(N__33532),
            .I(pin_out_6));
    InMux I__6596 (
            .O(N__33525),
            .I(N__33522));
    LocalMux I__6595 (
            .O(N__33522),
            .I(N__33519));
    Odrv4 I__6594 (
            .O(N__33519),
            .I(n7262));
    IoInMux I__6593 (
            .O(N__33516),
            .I(N__33513));
    LocalMux I__6592 (
            .O(N__33513),
            .I(N__33510));
    Span12Mux_s1_h I__6591 (
            .O(N__33510),
            .I(N__33506));
    CascadeMux I__6590 (
            .O(N__33509),
            .I(N__33503));
    Span12Mux_v I__6589 (
            .O(N__33506),
            .I(N__33499));
    InMux I__6588 (
            .O(N__33503),
            .I(N__33496));
    InMux I__6587 (
            .O(N__33502),
            .I(N__33493));
    Odrv12 I__6586 (
            .O(N__33499),
            .I(pin_out_7));
    LocalMux I__6585 (
            .O(N__33496),
            .I(pin_out_7));
    LocalMux I__6584 (
            .O(N__33493),
            .I(pin_out_7));
    InMux I__6583 (
            .O(N__33486),
            .I(N__33483));
    LocalMux I__6582 (
            .O(N__33483),
            .I(n8_adj_780));
    CascadeMux I__6581 (
            .O(N__33480),
            .I(n8_adj_780_cascade_));
    InMux I__6580 (
            .O(N__33477),
            .I(N__33474));
    LocalMux I__6579 (
            .O(N__33474),
            .I(n7274));
    InMux I__6578 (
            .O(N__33471),
            .I(N__33468));
    LocalMux I__6577 (
            .O(N__33468),
            .I(N__33465));
    Odrv4 I__6576 (
            .O(N__33465),
            .I(\nx.n2677 ));
    InMux I__6575 (
            .O(N__33462),
            .I(bfn_10_17_0_));
    CascadeMux I__6574 (
            .O(N__33459),
            .I(N__33456));
    InMux I__6573 (
            .O(N__33456),
            .I(N__33453));
    LocalMux I__6572 (
            .O(N__33453),
            .I(N__33450));
    Span4Mux_h I__6571 (
            .O(N__33450),
            .I(N__33447));
    Odrv4 I__6570 (
            .O(N__33447),
            .I(\nx.n2676 ));
    InMux I__6569 (
            .O(N__33444),
            .I(\nx.n10768 ));
    InMux I__6568 (
            .O(N__33441),
            .I(N__33438));
    LocalMux I__6567 (
            .O(N__33438),
            .I(N__33435));
    Span4Mux_v I__6566 (
            .O(N__33435),
            .I(N__33432));
    Odrv4 I__6565 (
            .O(N__33432),
            .I(\nx.n2675 ));
    InMux I__6564 (
            .O(N__33429),
            .I(\nx.n10769 ));
    InMux I__6563 (
            .O(N__33426),
            .I(N__33423));
    LocalMux I__6562 (
            .O(N__33423),
            .I(N__33420));
    Span4Mux_h I__6561 (
            .O(N__33420),
            .I(N__33417));
    Odrv4 I__6560 (
            .O(N__33417),
            .I(\nx.n2674 ));
    InMux I__6559 (
            .O(N__33414),
            .I(\nx.n10770 ));
    InMux I__6558 (
            .O(N__33411),
            .I(N__33408));
    LocalMux I__6557 (
            .O(N__33408),
            .I(N__33405));
    Span4Mux_h I__6556 (
            .O(N__33405),
            .I(N__33402));
    Odrv4 I__6555 (
            .O(N__33402),
            .I(\nx.n1668 ));
    CascadeMux I__6554 (
            .O(N__33399),
            .I(N__33396));
    InMux I__6553 (
            .O(N__33396),
            .I(N__33393));
    LocalMux I__6552 (
            .O(N__33393),
            .I(N__33389));
    CascadeMux I__6551 (
            .O(N__33392),
            .I(N__33386));
    Span4Mux_h I__6550 (
            .O(N__33389),
            .I(N__33382));
    InMux I__6549 (
            .O(N__33386),
            .I(N__33379));
    InMux I__6548 (
            .O(N__33385),
            .I(N__33376));
    Odrv4 I__6547 (
            .O(N__33382),
            .I(\nx.n1601 ));
    LocalMux I__6546 (
            .O(N__33379),
            .I(\nx.n1601 ));
    LocalMux I__6545 (
            .O(N__33376),
            .I(\nx.n1601 ));
    InMux I__6544 (
            .O(N__33369),
            .I(N__33366));
    LocalMux I__6543 (
            .O(N__33366),
            .I(N__33363));
    Span4Mux_h I__6542 (
            .O(N__33363),
            .I(N__33359));
    CascadeMux I__6541 (
            .O(N__33362),
            .I(N__33356));
    IoSpan4Mux I__6540 (
            .O(N__33359),
            .I(N__33353));
    InMux I__6539 (
            .O(N__33356),
            .I(N__33350));
    Span4Mux_s1_v I__6538 (
            .O(N__33353),
            .I(N__33345));
    LocalMux I__6537 (
            .O(N__33350),
            .I(N__33345));
    Span4Mux_h I__6536 (
            .O(N__33345),
            .I(N__33342));
    Odrv4 I__6535 (
            .O(N__33342),
            .I(\nx.n1509 ));
    CascadeMux I__6534 (
            .O(N__33339),
            .I(N__33336));
    InMux I__6533 (
            .O(N__33336),
            .I(N__33333));
    LocalMux I__6532 (
            .O(N__33333),
            .I(N__33330));
    Span4Mux_h I__6531 (
            .O(N__33330),
            .I(N__33327));
    Odrv4 I__6530 (
            .O(N__33327),
            .I(\nx.n1576 ));
    CascadeMux I__6529 (
            .O(N__33324),
            .I(\nx.n1608_cascade_ ));
    InMux I__6528 (
            .O(N__33321),
            .I(N__33318));
    LocalMux I__6527 (
            .O(N__33318),
            .I(N__33315));
    Odrv4 I__6526 (
            .O(N__33315),
            .I(\nx.n18 ));
    InMux I__6525 (
            .O(N__33312),
            .I(N__33309));
    LocalMux I__6524 (
            .O(N__33309),
            .I(N__33305));
    CascadeMux I__6523 (
            .O(N__33308),
            .I(N__33302));
    Span4Mux_v I__6522 (
            .O(N__33305),
            .I(N__33299));
    InMux I__6521 (
            .O(N__33302),
            .I(N__33296));
    Odrv4 I__6520 (
            .O(N__33299),
            .I(\nx.n1506 ));
    LocalMux I__6519 (
            .O(N__33296),
            .I(\nx.n1506 ));
    CascadeMux I__6518 (
            .O(N__33291),
            .I(N__33288));
    InMux I__6517 (
            .O(N__33288),
            .I(N__33285));
    LocalMux I__6516 (
            .O(N__33285),
            .I(N__33282));
    Span4Mux_h I__6515 (
            .O(N__33282),
            .I(N__33279));
    Odrv4 I__6514 (
            .O(N__33279),
            .I(\nx.n1573 ));
    CascadeMux I__6513 (
            .O(N__33276),
            .I(N__33267));
    CascadeMux I__6512 (
            .O(N__33275),
            .I(N__33264));
    CascadeMux I__6511 (
            .O(N__33274),
            .I(N__33259));
    CascadeMux I__6510 (
            .O(N__33273),
            .I(N__33256));
    CascadeMux I__6509 (
            .O(N__33272),
            .I(N__33252));
    InMux I__6508 (
            .O(N__33271),
            .I(N__33246));
    InMux I__6507 (
            .O(N__33270),
            .I(N__33246));
    InMux I__6506 (
            .O(N__33267),
            .I(N__33243));
    InMux I__6505 (
            .O(N__33264),
            .I(N__33236));
    InMux I__6504 (
            .O(N__33263),
            .I(N__33236));
    InMux I__6503 (
            .O(N__33262),
            .I(N__33236));
    InMux I__6502 (
            .O(N__33259),
            .I(N__33231));
    InMux I__6501 (
            .O(N__33256),
            .I(N__33231));
    InMux I__6500 (
            .O(N__33255),
            .I(N__33224));
    InMux I__6499 (
            .O(N__33252),
            .I(N__33224));
    InMux I__6498 (
            .O(N__33251),
            .I(N__33224));
    LocalMux I__6497 (
            .O(N__33246),
            .I(N__33221));
    LocalMux I__6496 (
            .O(N__33243),
            .I(N__33218));
    LocalMux I__6495 (
            .O(N__33236),
            .I(\nx.n1532 ));
    LocalMux I__6494 (
            .O(N__33231),
            .I(\nx.n1532 ));
    LocalMux I__6493 (
            .O(N__33224),
            .I(\nx.n1532 ));
    Odrv4 I__6492 (
            .O(N__33221),
            .I(\nx.n1532 ));
    Odrv12 I__6491 (
            .O(N__33218),
            .I(\nx.n1532 ));
    CascadeMux I__6490 (
            .O(N__33207),
            .I(N__33204));
    InMux I__6489 (
            .O(N__33204),
            .I(N__33200));
    InMux I__6488 (
            .O(N__33203),
            .I(N__33197));
    LocalMux I__6487 (
            .O(N__33200),
            .I(N__33193));
    LocalMux I__6486 (
            .O(N__33197),
            .I(N__33190));
    InMux I__6485 (
            .O(N__33196),
            .I(N__33187));
    Span4Mux_s3_v I__6484 (
            .O(N__33193),
            .I(N__33184));
    Odrv4 I__6483 (
            .O(N__33190),
            .I(\nx.n1605 ));
    LocalMux I__6482 (
            .O(N__33187),
            .I(\nx.n1605 ));
    Odrv4 I__6481 (
            .O(N__33184),
            .I(\nx.n1605 ));
    InMux I__6480 (
            .O(N__33177),
            .I(N__33173));
    CascadeMux I__6479 (
            .O(N__33176),
            .I(N__33169));
    LocalMux I__6478 (
            .O(N__33173),
            .I(N__33166));
    InMux I__6477 (
            .O(N__33172),
            .I(N__33163));
    InMux I__6476 (
            .O(N__33169),
            .I(N__33160));
    Odrv12 I__6475 (
            .O(N__33166),
            .I(\nx.n1604 ));
    LocalMux I__6474 (
            .O(N__33163),
            .I(\nx.n1604 ));
    LocalMux I__6473 (
            .O(N__33160),
            .I(\nx.n1604 ));
    CascadeMux I__6472 (
            .O(N__33153),
            .I(N__33150));
    InMux I__6471 (
            .O(N__33150),
            .I(N__33147));
    LocalMux I__6470 (
            .O(N__33147),
            .I(N__33144));
    Span4Mux_h I__6469 (
            .O(N__33144),
            .I(N__33141));
    Odrv4 I__6468 (
            .O(N__33141),
            .I(\nx.n1671 ));
    InMux I__6467 (
            .O(N__33138),
            .I(N__33134));
    CascadeMux I__6466 (
            .O(N__33137),
            .I(N__33131));
    LocalMux I__6465 (
            .O(N__33134),
            .I(N__33128));
    InMux I__6464 (
            .O(N__33131),
            .I(N__33125));
    Odrv4 I__6463 (
            .O(N__33128),
            .I(\nx.n1606 ));
    LocalMux I__6462 (
            .O(N__33125),
            .I(\nx.n1606 ));
    InMux I__6461 (
            .O(N__33120),
            .I(N__33117));
    LocalMux I__6460 (
            .O(N__33117),
            .I(N__33114));
    Span4Mux_h I__6459 (
            .O(N__33114),
            .I(N__33111));
    Odrv4 I__6458 (
            .O(N__33111),
            .I(\nx.n1673 ));
    CascadeMux I__6457 (
            .O(N__33108),
            .I(n21_cascade_));
    InMux I__6456 (
            .O(N__33105),
            .I(N__33102));
    LocalMux I__6455 (
            .O(N__33102),
            .I(N__33099));
    Span4Mux_h I__6454 (
            .O(N__33099),
            .I(N__33095));
    InMux I__6453 (
            .O(N__33098),
            .I(N__33092));
    Odrv4 I__6452 (
            .O(N__33095),
            .I(n6150));
    LocalMux I__6451 (
            .O(N__33092),
            .I(n6150));
    InMux I__6450 (
            .O(N__33087),
            .I(N__33084));
    LocalMux I__6449 (
            .O(N__33084),
            .I(N__33081));
    Odrv4 I__6448 (
            .O(N__33081),
            .I(\nx.n1870 ));
    InMux I__6447 (
            .O(N__33078),
            .I(\nx.n10634 ));
    InMux I__6446 (
            .O(N__33075),
            .I(N__33072));
    LocalMux I__6445 (
            .O(N__33072),
            .I(N__33069));
    Odrv4 I__6444 (
            .O(N__33069),
            .I(\nx.n1869 ));
    InMux I__6443 (
            .O(N__33066),
            .I(bfn_9_28_0_));
    InMux I__6442 (
            .O(N__33063),
            .I(N__33059));
    CascadeMux I__6441 (
            .O(N__33062),
            .I(N__33056));
    LocalMux I__6440 (
            .O(N__33059),
            .I(N__33053));
    InMux I__6439 (
            .O(N__33056),
            .I(N__33050));
    Span4Mux_h I__6438 (
            .O(N__33053),
            .I(N__33047));
    LocalMux I__6437 (
            .O(N__33050),
            .I(N__33044));
    Odrv4 I__6436 (
            .O(N__33047),
            .I(\nx.n1801 ));
    Odrv4 I__6435 (
            .O(N__33044),
            .I(\nx.n1801 ));
    CascadeMux I__6434 (
            .O(N__33039),
            .I(N__33036));
    InMux I__6433 (
            .O(N__33036),
            .I(N__33033));
    LocalMux I__6432 (
            .O(N__33033),
            .I(N__33030));
    Odrv4 I__6431 (
            .O(N__33030),
            .I(\nx.n1868 ));
    InMux I__6430 (
            .O(N__33027),
            .I(\nx.n10636 ));
    CascadeMux I__6429 (
            .O(N__33024),
            .I(N__33021));
    InMux I__6428 (
            .O(N__33021),
            .I(N__33017));
    InMux I__6427 (
            .O(N__33020),
            .I(N__33013));
    LocalMux I__6426 (
            .O(N__33017),
            .I(N__33010));
    InMux I__6425 (
            .O(N__33016),
            .I(N__33007));
    LocalMux I__6424 (
            .O(N__33013),
            .I(\nx.n1800 ));
    Odrv4 I__6423 (
            .O(N__33010),
            .I(\nx.n1800 ));
    LocalMux I__6422 (
            .O(N__33007),
            .I(\nx.n1800 ));
    CascadeMux I__6421 (
            .O(N__33000),
            .I(N__32997));
    InMux I__6420 (
            .O(N__32997),
            .I(N__32994));
    LocalMux I__6419 (
            .O(N__32994),
            .I(N__32991));
    Span4Mux_h I__6418 (
            .O(N__32991),
            .I(N__32988));
    Odrv4 I__6417 (
            .O(N__32988),
            .I(\nx.n1867 ));
    InMux I__6416 (
            .O(N__32985),
            .I(\nx.n10637 ));
    InMux I__6415 (
            .O(N__32982),
            .I(N__32979));
    LocalMux I__6414 (
            .O(N__32979),
            .I(N__32975));
    InMux I__6413 (
            .O(N__32978),
            .I(N__32972));
    Odrv4 I__6412 (
            .O(N__32975),
            .I(\nx.n1799 ));
    LocalMux I__6411 (
            .O(N__32972),
            .I(\nx.n1799 ));
    InMux I__6410 (
            .O(N__32967),
            .I(N__32964));
    LocalMux I__6409 (
            .O(N__32964),
            .I(N__32961));
    Odrv4 I__6408 (
            .O(N__32961),
            .I(\nx.n1866 ));
    InMux I__6407 (
            .O(N__32958),
            .I(\nx.n10638 ));
    InMux I__6406 (
            .O(N__32955),
            .I(N__32952));
    LocalMux I__6405 (
            .O(N__32952),
            .I(N__32949));
    Span4Mux_h I__6404 (
            .O(N__32949),
            .I(N__32946));
    Odrv4 I__6403 (
            .O(N__32946),
            .I(\nx.n1865 ));
    InMux I__6402 (
            .O(N__32943),
            .I(\nx.n10639 ));
    CascadeMux I__6401 (
            .O(N__32940),
            .I(N__32937));
    InMux I__6400 (
            .O(N__32937),
            .I(N__32934));
    LocalMux I__6399 (
            .O(N__32934),
            .I(N__32930));
    InMux I__6398 (
            .O(N__32933),
            .I(N__32927));
    Odrv4 I__6397 (
            .O(N__32930),
            .I(\nx.n1797 ));
    LocalMux I__6396 (
            .O(N__32927),
            .I(\nx.n1797 ));
    InMux I__6395 (
            .O(N__32922),
            .I(N__32919));
    LocalMux I__6394 (
            .O(N__32919),
            .I(N__32916));
    Odrv4 I__6393 (
            .O(N__32916),
            .I(\nx.n1864 ));
    InMux I__6392 (
            .O(N__32913),
            .I(\nx.n10640 ));
    CascadeMux I__6391 (
            .O(N__32910),
            .I(N__32907));
    InMux I__6390 (
            .O(N__32907),
            .I(N__32904));
    LocalMux I__6389 (
            .O(N__32904),
            .I(N__32893));
    InMux I__6388 (
            .O(N__32903),
            .I(N__32888));
    InMux I__6387 (
            .O(N__32902),
            .I(N__32888));
    CascadeMux I__6386 (
            .O(N__32901),
            .I(N__32884));
    CascadeMux I__6385 (
            .O(N__32900),
            .I(N__32879));
    CascadeMux I__6384 (
            .O(N__32899),
            .I(N__32875));
    InMux I__6383 (
            .O(N__32898),
            .I(N__32867));
    InMux I__6382 (
            .O(N__32897),
            .I(N__32867));
    InMux I__6381 (
            .O(N__32896),
            .I(N__32867));
    Span4Mux_v I__6380 (
            .O(N__32893),
            .I(N__32862));
    LocalMux I__6379 (
            .O(N__32888),
            .I(N__32862));
    InMux I__6378 (
            .O(N__32887),
            .I(N__32859));
    InMux I__6377 (
            .O(N__32884),
            .I(N__32854));
    InMux I__6376 (
            .O(N__32883),
            .I(N__32854));
    InMux I__6375 (
            .O(N__32882),
            .I(N__32851));
    InMux I__6374 (
            .O(N__32879),
            .I(N__32842));
    InMux I__6373 (
            .O(N__32878),
            .I(N__32842));
    InMux I__6372 (
            .O(N__32875),
            .I(N__32842));
    InMux I__6371 (
            .O(N__32874),
            .I(N__32842));
    LocalMux I__6370 (
            .O(N__32867),
            .I(N__32839));
    Span4Mux_h I__6369 (
            .O(N__32862),
            .I(N__32836));
    LocalMux I__6368 (
            .O(N__32859),
            .I(\nx.n1829 ));
    LocalMux I__6367 (
            .O(N__32854),
            .I(\nx.n1829 ));
    LocalMux I__6366 (
            .O(N__32851),
            .I(\nx.n1829 ));
    LocalMux I__6365 (
            .O(N__32842),
            .I(\nx.n1829 ));
    Odrv4 I__6364 (
            .O(N__32839),
            .I(\nx.n1829 ));
    Odrv4 I__6363 (
            .O(N__32836),
            .I(\nx.n1829 ));
    InMux I__6362 (
            .O(N__32823),
            .I(\nx.n10641 ));
    InMux I__6361 (
            .O(N__32820),
            .I(N__32816));
    InMux I__6360 (
            .O(N__32819),
            .I(N__32813));
    LocalMux I__6359 (
            .O(N__32816),
            .I(N__32807));
    LocalMux I__6358 (
            .O(N__32813),
            .I(N__32807));
    InMux I__6357 (
            .O(N__32812),
            .I(N__32804));
    Span4Mux_h I__6356 (
            .O(N__32807),
            .I(N__32801));
    LocalMux I__6355 (
            .O(N__32804),
            .I(N__32798));
    Odrv4 I__6354 (
            .O(N__32801),
            .I(\nx.n1895 ));
    Odrv12 I__6353 (
            .O(N__32798),
            .I(\nx.n1895 ));
    InMux I__6352 (
            .O(N__32793),
            .I(N__32788));
    InMux I__6351 (
            .O(N__32792),
            .I(N__32785));
    CascadeMux I__6350 (
            .O(N__32791),
            .I(N__32782));
    LocalMux I__6349 (
            .O(N__32788),
            .I(N__32777));
    LocalMux I__6348 (
            .O(N__32785),
            .I(N__32777));
    InMux I__6347 (
            .O(N__32782),
            .I(N__32774));
    Odrv4 I__6346 (
            .O(N__32777),
            .I(\nx.n1896 ));
    LocalMux I__6345 (
            .O(N__32774),
            .I(\nx.n1896 ));
    InMux I__6344 (
            .O(N__32769),
            .I(N__32766));
    LocalMux I__6343 (
            .O(N__32766),
            .I(N__32760));
    InMux I__6342 (
            .O(N__32765),
            .I(N__32757));
    InMux I__6341 (
            .O(N__32764),
            .I(N__32754));
    InMux I__6340 (
            .O(N__32763),
            .I(N__32751));
    Span4Mux_h I__6339 (
            .O(N__32760),
            .I(N__32746));
    LocalMux I__6338 (
            .O(N__32757),
            .I(N__32746));
    LocalMux I__6337 (
            .O(N__32754),
            .I(N__32740));
    LocalMux I__6336 (
            .O(N__32751),
            .I(N__32740));
    Span4Mux_h I__6335 (
            .O(N__32746),
            .I(N__32737));
    InMux I__6334 (
            .O(N__32745),
            .I(N__32734));
    Span4Mux_h I__6333 (
            .O(N__32740),
            .I(N__32731));
    Span4Mux_h I__6332 (
            .O(N__32737),
            .I(N__32728));
    LocalMux I__6331 (
            .O(N__32734),
            .I(\nx.bit_ctr_17 ));
    Odrv4 I__6330 (
            .O(N__32731),
            .I(\nx.bit_ctr_17 ));
    Odrv4 I__6329 (
            .O(N__32728),
            .I(\nx.bit_ctr_17 ));
    InMux I__6328 (
            .O(N__32721),
            .I(N__32718));
    LocalMux I__6327 (
            .O(N__32718),
            .I(N__32714));
    InMux I__6326 (
            .O(N__32717),
            .I(N__32711));
    Span4Mux_h I__6325 (
            .O(N__32714),
            .I(N__32705));
    LocalMux I__6324 (
            .O(N__32711),
            .I(N__32702));
    InMux I__6323 (
            .O(N__32710),
            .I(N__32699));
    InMux I__6322 (
            .O(N__32709),
            .I(N__32694));
    InMux I__6321 (
            .O(N__32708),
            .I(N__32694));
    Span4Mux_h I__6320 (
            .O(N__32705),
            .I(N__32689));
    Span4Mux_s3_h I__6319 (
            .O(N__32702),
            .I(N__32689));
    LocalMux I__6318 (
            .O(N__32699),
            .I(\nx.bit_ctr_22 ));
    LocalMux I__6317 (
            .O(N__32694),
            .I(\nx.bit_ctr_22 ));
    Odrv4 I__6316 (
            .O(N__32689),
            .I(\nx.bit_ctr_22 ));
    InMux I__6315 (
            .O(N__32682),
            .I(N__32679));
    LocalMux I__6314 (
            .O(N__32679),
            .I(N__32676));
    Span4Mux_h I__6313 (
            .O(N__32676),
            .I(N__32673));
    Span4Mux_h I__6312 (
            .O(N__32673),
            .I(N__32670));
    Odrv4 I__6311 (
            .O(N__32670),
            .I(\nx.n30_adj_703 ));
    CascadeMux I__6310 (
            .O(N__32667),
            .I(N__32663));
    InMux I__6309 (
            .O(N__32666),
            .I(N__32659));
    InMux I__6308 (
            .O(N__32663),
            .I(N__32656));
    InMux I__6307 (
            .O(N__32662),
            .I(N__32653));
    LocalMux I__6306 (
            .O(N__32659),
            .I(N__32648));
    LocalMux I__6305 (
            .O(N__32656),
            .I(N__32648));
    LocalMux I__6304 (
            .O(N__32653),
            .I(\nx.n1809 ));
    Odrv4 I__6303 (
            .O(N__32648),
            .I(\nx.n1809 ));
    InMux I__6302 (
            .O(N__32643),
            .I(N__32640));
    LocalMux I__6301 (
            .O(N__32640),
            .I(N__32637));
    Span4Mux_v I__6300 (
            .O(N__32637),
            .I(N__32634));
    Odrv4 I__6299 (
            .O(N__32634),
            .I(\nx.n1876 ));
    InMux I__6298 (
            .O(N__32631),
            .I(\nx.n10628 ));
    CascadeMux I__6297 (
            .O(N__32628),
            .I(N__32625));
    InMux I__6296 (
            .O(N__32625),
            .I(N__32620));
    InMux I__6295 (
            .O(N__32624),
            .I(N__32615));
    InMux I__6294 (
            .O(N__32623),
            .I(N__32615));
    LocalMux I__6293 (
            .O(N__32620),
            .I(N__32612));
    LocalMux I__6292 (
            .O(N__32615),
            .I(\nx.n1808 ));
    Odrv12 I__6291 (
            .O(N__32612),
            .I(\nx.n1808 ));
    InMux I__6290 (
            .O(N__32607),
            .I(N__32604));
    LocalMux I__6289 (
            .O(N__32604),
            .I(N__32601));
    Span4Mux_h I__6288 (
            .O(N__32601),
            .I(N__32598));
    Odrv4 I__6287 (
            .O(N__32598),
            .I(\nx.n1875 ));
    InMux I__6286 (
            .O(N__32595),
            .I(\nx.n10629 ));
    CascadeMux I__6285 (
            .O(N__32592),
            .I(N__32589));
    InMux I__6284 (
            .O(N__32589),
            .I(N__32582));
    InMux I__6283 (
            .O(N__32588),
            .I(N__32582));
    CascadeMux I__6282 (
            .O(N__32587),
            .I(N__32579));
    LocalMux I__6281 (
            .O(N__32582),
            .I(N__32576));
    InMux I__6280 (
            .O(N__32579),
            .I(N__32573));
    Odrv4 I__6279 (
            .O(N__32576),
            .I(\nx.n1807 ));
    LocalMux I__6278 (
            .O(N__32573),
            .I(\nx.n1807 ));
    InMux I__6277 (
            .O(N__32568),
            .I(N__32565));
    LocalMux I__6276 (
            .O(N__32565),
            .I(N__32562));
    Span4Mux_h I__6275 (
            .O(N__32562),
            .I(N__32559));
    Odrv4 I__6274 (
            .O(N__32559),
            .I(\nx.n1874 ));
    InMux I__6273 (
            .O(N__32556),
            .I(\nx.n10630 ));
    CascadeMux I__6272 (
            .O(N__32553),
            .I(N__32550));
    InMux I__6271 (
            .O(N__32550),
            .I(N__32547));
    LocalMux I__6270 (
            .O(N__32547),
            .I(N__32544));
    Odrv4 I__6269 (
            .O(N__32544),
            .I(\nx.n1873 ));
    InMux I__6268 (
            .O(N__32541),
            .I(\nx.n10631 ));
    InMux I__6267 (
            .O(N__32538),
            .I(N__32534));
    CascadeMux I__6266 (
            .O(N__32537),
            .I(N__32531));
    LocalMux I__6265 (
            .O(N__32534),
            .I(N__32527));
    InMux I__6264 (
            .O(N__32531),
            .I(N__32524));
    InMux I__6263 (
            .O(N__32530),
            .I(N__32521));
    Span4Mux_v I__6262 (
            .O(N__32527),
            .I(N__32516));
    LocalMux I__6261 (
            .O(N__32524),
            .I(N__32516));
    LocalMux I__6260 (
            .O(N__32521),
            .I(\nx.n1805 ));
    Odrv4 I__6259 (
            .O(N__32516),
            .I(\nx.n1805 ));
    CascadeMux I__6258 (
            .O(N__32511),
            .I(N__32508));
    InMux I__6257 (
            .O(N__32508),
            .I(N__32505));
    LocalMux I__6256 (
            .O(N__32505),
            .I(N__32502));
    Span4Mux_v I__6255 (
            .O(N__32502),
            .I(N__32499));
    Span4Mux_h I__6254 (
            .O(N__32499),
            .I(N__32496));
    Odrv4 I__6253 (
            .O(N__32496),
            .I(\nx.n1872 ));
    InMux I__6252 (
            .O(N__32493),
            .I(\nx.n10632 ));
    CascadeMux I__6251 (
            .O(N__32490),
            .I(N__32487));
    InMux I__6250 (
            .O(N__32487),
            .I(N__32483));
    InMux I__6249 (
            .O(N__32486),
            .I(N__32480));
    LocalMux I__6248 (
            .O(N__32483),
            .I(N__32477));
    LocalMux I__6247 (
            .O(N__32480),
            .I(\nx.n1804 ));
    Odrv4 I__6246 (
            .O(N__32477),
            .I(\nx.n1804 ));
    InMux I__6245 (
            .O(N__32472),
            .I(N__32469));
    LocalMux I__6244 (
            .O(N__32469),
            .I(N__32466));
    Span4Mux_h I__6243 (
            .O(N__32466),
            .I(N__32463));
    Odrv4 I__6242 (
            .O(N__32463),
            .I(\nx.n1871 ));
    InMux I__6241 (
            .O(N__32460),
            .I(\nx.n10633 ));
    InMux I__6240 (
            .O(N__32457),
            .I(N__32453));
    InMux I__6239 (
            .O(N__32456),
            .I(N__32450));
    LocalMux I__6238 (
            .O(N__32453),
            .I(N__32444));
    LocalMux I__6237 (
            .O(N__32450),
            .I(N__32444));
    InMux I__6236 (
            .O(N__32449),
            .I(N__32441));
    Span4Mux_h I__6235 (
            .O(N__32444),
            .I(N__32438));
    LocalMux I__6234 (
            .O(N__32441),
            .I(N__32435));
    Odrv4 I__6233 (
            .O(N__32438),
            .I(\nx.n1901 ));
    Odrv4 I__6232 (
            .O(N__32435),
            .I(\nx.n1901 ));
    InMux I__6231 (
            .O(N__32430),
            .I(N__32426));
    InMux I__6230 (
            .O(N__32429),
            .I(N__32423));
    LocalMux I__6229 (
            .O(N__32426),
            .I(N__32417));
    LocalMux I__6228 (
            .O(N__32423),
            .I(N__32417));
    InMux I__6227 (
            .O(N__32422),
            .I(N__32414));
    Odrv4 I__6226 (
            .O(N__32417),
            .I(\nx.n1905 ));
    LocalMux I__6225 (
            .O(N__32414),
            .I(\nx.n1905 ));
    InMux I__6224 (
            .O(N__32409),
            .I(N__32406));
    LocalMux I__6223 (
            .O(N__32406),
            .I(N__32403));
    Odrv4 I__6222 (
            .O(N__32403),
            .I(\nx.n25_adj_606 ));
    CascadeMux I__6221 (
            .O(N__32400),
            .I(N__32397));
    InMux I__6220 (
            .O(N__32397),
            .I(N__32394));
    LocalMux I__6219 (
            .O(N__32394),
            .I(N__32391));
    Odrv12 I__6218 (
            .O(N__32391),
            .I(\nx.n22 ));
    InMux I__6217 (
            .O(N__32388),
            .I(N__32384));
    InMux I__6216 (
            .O(N__32387),
            .I(N__32381));
    LocalMux I__6215 (
            .O(N__32384),
            .I(N__32375));
    LocalMux I__6214 (
            .O(N__32381),
            .I(N__32375));
    InMux I__6213 (
            .O(N__32380),
            .I(N__32372));
    Odrv4 I__6212 (
            .O(N__32375),
            .I(\nx.n1900 ));
    LocalMux I__6211 (
            .O(N__32372),
            .I(\nx.n1900 ));
    CascadeMux I__6210 (
            .O(N__32367),
            .I(\nx.n1799_cascade_ ));
    InMux I__6209 (
            .O(N__32364),
            .I(N__32360));
    InMux I__6208 (
            .O(N__32363),
            .I(N__32357));
    LocalMux I__6207 (
            .O(N__32360),
            .I(N__32351));
    LocalMux I__6206 (
            .O(N__32357),
            .I(N__32351));
    InMux I__6205 (
            .O(N__32356),
            .I(N__32348));
    Span4Mux_h I__6204 (
            .O(N__32351),
            .I(N__32345));
    LocalMux I__6203 (
            .O(N__32348),
            .I(N__32342));
    Odrv4 I__6202 (
            .O(N__32345),
            .I(\nx.n1898 ));
    Odrv12 I__6201 (
            .O(N__32342),
            .I(\nx.n1898 ));
    CascadeMux I__6200 (
            .O(N__32337),
            .I(\nx.n1797_cascade_ ));
    CascadeMux I__6199 (
            .O(N__32334),
            .I(N__32329));
    InMux I__6198 (
            .O(N__32333),
            .I(N__32324));
    InMux I__6197 (
            .O(N__32332),
            .I(N__32324));
    InMux I__6196 (
            .O(N__32329),
            .I(N__32321));
    LocalMux I__6195 (
            .O(N__32324),
            .I(N__32318));
    LocalMux I__6194 (
            .O(N__32321),
            .I(N__32315));
    Span4Mux_h I__6193 (
            .O(N__32318),
            .I(N__32312));
    Span4Mux_h I__6192 (
            .O(N__32315),
            .I(N__32309));
    Odrv4 I__6191 (
            .O(N__32312),
            .I(\nx.n2001 ));
    Odrv4 I__6190 (
            .O(N__32309),
            .I(\nx.n2001 ));
    InMux I__6189 (
            .O(N__32304),
            .I(N__32301));
    LocalMux I__6188 (
            .O(N__32301),
            .I(N__32298));
    Odrv4 I__6187 (
            .O(N__32298),
            .I(\nx.n2068 ));
    InMux I__6186 (
            .O(N__32295),
            .I(\nx.n10665 ));
    CascadeMux I__6185 (
            .O(N__32292),
            .I(N__32288));
    CascadeMux I__6184 (
            .O(N__32291),
            .I(N__32284));
    InMux I__6183 (
            .O(N__32288),
            .I(N__32279));
    InMux I__6182 (
            .O(N__32287),
            .I(N__32279));
    InMux I__6181 (
            .O(N__32284),
            .I(N__32276));
    LocalMux I__6180 (
            .O(N__32279),
            .I(N__32273));
    LocalMux I__6179 (
            .O(N__32276),
            .I(N__32270));
    Span4Mux_h I__6178 (
            .O(N__32273),
            .I(N__32267));
    Span4Mux_h I__6177 (
            .O(N__32270),
            .I(N__32264));
    Odrv4 I__6176 (
            .O(N__32267),
            .I(\nx.n2000 ));
    Odrv4 I__6175 (
            .O(N__32264),
            .I(\nx.n2000 ));
    InMux I__6174 (
            .O(N__32259),
            .I(N__32256));
    LocalMux I__6173 (
            .O(N__32256),
            .I(N__32253));
    Odrv4 I__6172 (
            .O(N__32253),
            .I(\nx.n2067 ));
    InMux I__6171 (
            .O(N__32250),
            .I(\nx.n10666 ));
    CascadeMux I__6170 (
            .O(N__32247),
            .I(N__32242));
    CascadeMux I__6169 (
            .O(N__32246),
            .I(N__32239));
    InMux I__6168 (
            .O(N__32245),
            .I(N__32234));
    InMux I__6167 (
            .O(N__32242),
            .I(N__32234));
    InMux I__6166 (
            .O(N__32239),
            .I(N__32231));
    LocalMux I__6165 (
            .O(N__32234),
            .I(N__32228));
    LocalMux I__6164 (
            .O(N__32231),
            .I(N__32225));
    Span4Mux_h I__6163 (
            .O(N__32228),
            .I(N__32222));
    Span4Mux_v I__6162 (
            .O(N__32225),
            .I(N__32219));
    Odrv4 I__6161 (
            .O(N__32222),
            .I(\nx.n1999 ));
    Odrv4 I__6160 (
            .O(N__32219),
            .I(\nx.n1999 ));
    InMux I__6159 (
            .O(N__32214),
            .I(N__32211));
    LocalMux I__6158 (
            .O(N__32211),
            .I(N__32208));
    Odrv4 I__6157 (
            .O(N__32208),
            .I(\nx.n2066 ));
    InMux I__6156 (
            .O(N__32205),
            .I(\nx.n10667 ));
    InMux I__6155 (
            .O(N__32202),
            .I(\nx.n10668 ));
    InMux I__6154 (
            .O(N__32199),
            .I(\nx.n10669 ));
    InMux I__6153 (
            .O(N__32196),
            .I(N__32192));
    CascadeMux I__6152 (
            .O(N__32195),
            .I(N__32189));
    LocalMux I__6151 (
            .O(N__32192),
            .I(N__32186));
    InMux I__6150 (
            .O(N__32189),
            .I(N__32183));
    Span4Mux_h I__6149 (
            .O(N__32186),
            .I(N__32179));
    LocalMux I__6148 (
            .O(N__32183),
            .I(N__32176));
    InMux I__6147 (
            .O(N__32182),
            .I(N__32173));
    Span4Mux_v I__6146 (
            .O(N__32179),
            .I(N__32170));
    Span4Mux_h I__6145 (
            .O(N__32176),
            .I(N__32167));
    LocalMux I__6144 (
            .O(N__32173),
            .I(N__32164));
    Odrv4 I__6143 (
            .O(N__32170),
            .I(\nx.n1996 ));
    Odrv4 I__6142 (
            .O(N__32167),
            .I(\nx.n1996 ));
    Odrv12 I__6141 (
            .O(N__32164),
            .I(\nx.n1996 ));
    CascadeMux I__6140 (
            .O(N__32157),
            .I(N__32154));
    InMux I__6139 (
            .O(N__32154),
            .I(N__32151));
    LocalMux I__6138 (
            .O(N__32151),
            .I(N__32148));
    Span4Mux_h I__6137 (
            .O(N__32148),
            .I(N__32145));
    Odrv4 I__6136 (
            .O(N__32145),
            .I(\nx.n2063 ));
    InMux I__6135 (
            .O(N__32142),
            .I(\nx.n10670 ));
    InMux I__6134 (
            .O(N__32139),
            .I(\nx.n10671 ));
    CascadeMux I__6133 (
            .O(N__32136),
            .I(N__32133));
    InMux I__6132 (
            .O(N__32133),
            .I(N__32130));
    LocalMux I__6131 (
            .O(N__32130),
            .I(N__32126));
    InMux I__6130 (
            .O(N__32129),
            .I(N__32123));
    Span4Mux_h I__6129 (
            .O(N__32126),
            .I(N__32120));
    LocalMux I__6128 (
            .O(N__32123),
            .I(N__32117));
    Odrv4 I__6127 (
            .O(N__32120),
            .I(\nx.n1994 ));
    Odrv12 I__6126 (
            .O(N__32117),
            .I(\nx.n1994 ));
    InMux I__6125 (
            .O(N__32112),
            .I(bfn_9_25_0_));
    InMux I__6124 (
            .O(N__32109),
            .I(bfn_9_23_0_));
    InMux I__6123 (
            .O(N__32106),
            .I(\nx.n10657 ));
    InMux I__6122 (
            .O(N__32103),
            .I(\nx.n10658 ));
    InMux I__6121 (
            .O(N__32100),
            .I(\nx.n10659 ));
    InMux I__6120 (
            .O(N__32097),
            .I(N__32093));
    CascadeMux I__6119 (
            .O(N__32096),
            .I(N__32090));
    LocalMux I__6118 (
            .O(N__32093),
            .I(N__32086));
    InMux I__6117 (
            .O(N__32090),
            .I(N__32083));
    CascadeMux I__6116 (
            .O(N__32089),
            .I(N__32080));
    Span4Mux_h I__6115 (
            .O(N__32086),
            .I(N__32077));
    LocalMux I__6114 (
            .O(N__32083),
            .I(N__32074));
    InMux I__6113 (
            .O(N__32080),
            .I(N__32071));
    Span4Mux_v I__6112 (
            .O(N__32077),
            .I(N__32066));
    Span4Mux_v I__6111 (
            .O(N__32074),
            .I(N__32066));
    LocalMux I__6110 (
            .O(N__32071),
            .I(\nx.n2006 ));
    Odrv4 I__6109 (
            .O(N__32066),
            .I(\nx.n2006 ));
    InMux I__6108 (
            .O(N__32061),
            .I(N__32058));
    LocalMux I__6107 (
            .O(N__32058),
            .I(N__32055));
    Odrv12 I__6106 (
            .O(N__32055),
            .I(\nx.n2073 ));
    InMux I__6105 (
            .O(N__32052),
            .I(\nx.n10660 ));
    CascadeMux I__6104 (
            .O(N__32049),
            .I(N__32045));
    CascadeMux I__6103 (
            .O(N__32048),
            .I(N__32042));
    InMux I__6102 (
            .O(N__32045),
            .I(N__32039));
    InMux I__6101 (
            .O(N__32042),
            .I(N__32036));
    LocalMux I__6100 (
            .O(N__32039),
            .I(N__32033));
    LocalMux I__6099 (
            .O(N__32036),
            .I(N__32029));
    Span4Mux_h I__6098 (
            .O(N__32033),
            .I(N__32026));
    InMux I__6097 (
            .O(N__32032),
            .I(N__32023));
    Span4Mux_h I__6096 (
            .O(N__32029),
            .I(N__32020));
    Odrv4 I__6095 (
            .O(N__32026),
            .I(\nx.n2005 ));
    LocalMux I__6094 (
            .O(N__32023),
            .I(\nx.n2005 ));
    Odrv4 I__6093 (
            .O(N__32020),
            .I(\nx.n2005 ));
    InMux I__6092 (
            .O(N__32013),
            .I(N__32010));
    LocalMux I__6091 (
            .O(N__32010),
            .I(N__32007));
    Odrv4 I__6090 (
            .O(N__32007),
            .I(\nx.n2072 ));
    InMux I__6089 (
            .O(N__32004),
            .I(\nx.n10661 ));
    CascadeMux I__6088 (
            .O(N__32001),
            .I(N__31997));
    CascadeMux I__6087 (
            .O(N__32000),
            .I(N__31994));
    InMux I__6086 (
            .O(N__31997),
            .I(N__31991));
    InMux I__6085 (
            .O(N__31994),
            .I(N__31988));
    LocalMux I__6084 (
            .O(N__31991),
            .I(N__31985));
    LocalMux I__6083 (
            .O(N__31988),
            .I(N__31981));
    Span4Mux_v I__6082 (
            .O(N__31985),
            .I(N__31978));
    InMux I__6081 (
            .O(N__31984),
            .I(N__31975));
    Span4Mux_h I__6080 (
            .O(N__31981),
            .I(N__31972));
    Odrv4 I__6079 (
            .O(N__31978),
            .I(\nx.n2004 ));
    LocalMux I__6078 (
            .O(N__31975),
            .I(\nx.n2004 ));
    Odrv4 I__6077 (
            .O(N__31972),
            .I(\nx.n2004 ));
    InMux I__6076 (
            .O(N__31965),
            .I(N__31962));
    LocalMux I__6075 (
            .O(N__31962),
            .I(\nx.n2071 ));
    InMux I__6074 (
            .O(N__31959),
            .I(\nx.n10662 ));
    InMux I__6073 (
            .O(N__31956),
            .I(\nx.n10663 ));
    InMux I__6072 (
            .O(N__31953),
            .I(bfn_9_24_0_));
    CascadeMux I__6071 (
            .O(N__31950),
            .I(\nx.n2595_cascade_ ));
    InMux I__6070 (
            .O(N__31947),
            .I(N__31944));
    LocalMux I__6069 (
            .O(N__31944),
            .I(N__31941));
    Span4Mux_h I__6068 (
            .O(N__31941),
            .I(N__31938));
    Odrv4 I__6067 (
            .O(N__31938),
            .I(\nx.n28_adj_663 ));
    CascadeMux I__6066 (
            .O(N__31935),
            .I(\nx.n26_adj_664_cascade_ ));
    InMux I__6065 (
            .O(N__31932),
            .I(N__31929));
    LocalMux I__6064 (
            .O(N__31929),
            .I(N__31926));
    Odrv4 I__6063 (
            .O(N__31926),
            .I(\nx.n25_adj_666 ));
    CascadeMux I__6062 (
            .O(N__31923),
            .I(\nx.n2027_cascade_ ));
    CascadeMux I__6061 (
            .O(N__31920),
            .I(\nx.n2099_cascade_ ));
    InMux I__6060 (
            .O(N__31917),
            .I(N__31914));
    LocalMux I__6059 (
            .O(N__31914),
            .I(N__31910));
    CascadeMux I__6058 (
            .O(N__31913),
            .I(N__31907));
    Span4Mux_h I__6057 (
            .O(N__31910),
            .I(N__31903));
    InMux I__6056 (
            .O(N__31907),
            .I(N__31900));
    InMux I__6055 (
            .O(N__31906),
            .I(N__31897));
    Odrv4 I__6054 (
            .O(N__31903),
            .I(\nx.n2904 ));
    LocalMux I__6053 (
            .O(N__31900),
            .I(\nx.n2904 ));
    LocalMux I__6052 (
            .O(N__31897),
            .I(\nx.n2904 ));
    CascadeMux I__6051 (
            .O(N__31890),
            .I(N__31887));
    InMux I__6050 (
            .O(N__31887),
            .I(N__31884));
    LocalMux I__6049 (
            .O(N__31884),
            .I(N__31881));
    Odrv12 I__6048 (
            .O(N__31881),
            .I(\nx.n2971 ));
    InMux I__6047 (
            .O(N__31878),
            .I(N__31871));
    CascadeMux I__6046 (
            .O(N__31877),
            .I(N__31868));
    CascadeMux I__6045 (
            .O(N__31876),
            .I(N__31860));
    CascadeMux I__6044 (
            .O(N__31875),
            .I(N__31855));
    InMux I__6043 (
            .O(N__31874),
            .I(N__31848));
    LocalMux I__6042 (
            .O(N__31871),
            .I(N__31845));
    InMux I__6041 (
            .O(N__31868),
            .I(N__31840));
    InMux I__6040 (
            .O(N__31867),
            .I(N__31840));
    CascadeMux I__6039 (
            .O(N__31866),
            .I(N__31830));
    CascadeMux I__6038 (
            .O(N__31865),
            .I(N__31827));
    CascadeMux I__6037 (
            .O(N__31864),
            .I(N__31823));
    CascadeMux I__6036 (
            .O(N__31863),
            .I(N__31819));
    InMux I__6035 (
            .O(N__31860),
            .I(N__31814));
    InMux I__6034 (
            .O(N__31859),
            .I(N__31814));
    InMux I__6033 (
            .O(N__31858),
            .I(N__31807));
    InMux I__6032 (
            .O(N__31855),
            .I(N__31807));
    InMux I__6031 (
            .O(N__31854),
            .I(N__31807));
    InMux I__6030 (
            .O(N__31853),
            .I(N__31800));
    InMux I__6029 (
            .O(N__31852),
            .I(N__31800));
    InMux I__6028 (
            .O(N__31851),
            .I(N__31800));
    LocalMux I__6027 (
            .O(N__31848),
            .I(N__31797));
    Span4Mux_v I__6026 (
            .O(N__31845),
            .I(N__31794));
    LocalMux I__6025 (
            .O(N__31840),
            .I(N__31791));
    InMux I__6024 (
            .O(N__31839),
            .I(N__31784));
    InMux I__6023 (
            .O(N__31838),
            .I(N__31784));
    InMux I__6022 (
            .O(N__31837),
            .I(N__31784));
    InMux I__6021 (
            .O(N__31836),
            .I(N__31775));
    InMux I__6020 (
            .O(N__31835),
            .I(N__31775));
    InMux I__6019 (
            .O(N__31834),
            .I(N__31775));
    InMux I__6018 (
            .O(N__31833),
            .I(N__31775));
    InMux I__6017 (
            .O(N__31830),
            .I(N__31762));
    InMux I__6016 (
            .O(N__31827),
            .I(N__31762));
    InMux I__6015 (
            .O(N__31826),
            .I(N__31762));
    InMux I__6014 (
            .O(N__31823),
            .I(N__31762));
    InMux I__6013 (
            .O(N__31822),
            .I(N__31762));
    InMux I__6012 (
            .O(N__31819),
            .I(N__31762));
    LocalMux I__6011 (
            .O(N__31814),
            .I(N__31759));
    LocalMux I__6010 (
            .O(N__31807),
            .I(N__31756));
    LocalMux I__6009 (
            .O(N__31800),
            .I(N__31749));
    Span4Mux_s1_h I__6008 (
            .O(N__31797),
            .I(N__31749));
    Span4Mux_h I__6007 (
            .O(N__31794),
            .I(N__31749));
    Odrv4 I__6006 (
            .O(N__31791),
            .I(\nx.n2918 ));
    LocalMux I__6005 (
            .O(N__31784),
            .I(\nx.n2918 ));
    LocalMux I__6004 (
            .O(N__31775),
            .I(\nx.n2918 ));
    LocalMux I__6003 (
            .O(N__31762),
            .I(\nx.n2918 ));
    Odrv4 I__6002 (
            .O(N__31759),
            .I(\nx.n2918 ));
    Odrv4 I__6001 (
            .O(N__31756),
            .I(\nx.n2918 ));
    Odrv4 I__6000 (
            .O(N__31749),
            .I(\nx.n2918 ));
    CascadeMux I__5999 (
            .O(N__31734),
            .I(N__31729));
    InMux I__5998 (
            .O(N__31733),
            .I(N__31726));
    InMux I__5997 (
            .O(N__31732),
            .I(N__31723));
    InMux I__5996 (
            .O(N__31729),
            .I(N__31720));
    LocalMux I__5995 (
            .O(N__31726),
            .I(N__31717));
    LocalMux I__5994 (
            .O(N__31723),
            .I(N__31714));
    LocalMux I__5993 (
            .O(N__31720),
            .I(N__31711));
    Span4Mux_h I__5992 (
            .O(N__31717),
            .I(N__31708));
    Span4Mux_v I__5991 (
            .O(N__31714),
            .I(N__31703));
    Span4Mux_v I__5990 (
            .O(N__31711),
            .I(N__31703));
    Span4Mux_h I__5989 (
            .O(N__31708),
            .I(N__31700));
    Span4Mux_h I__5988 (
            .O(N__31703),
            .I(N__31697));
    Odrv4 I__5987 (
            .O(N__31700),
            .I(\nx.n3003 ));
    Odrv4 I__5986 (
            .O(N__31697),
            .I(\nx.n3003 ));
    CascadeMux I__5985 (
            .O(N__31692),
            .I(N__31689));
    InMux I__5984 (
            .O(N__31689),
            .I(N__31685));
    InMux I__5983 (
            .O(N__31688),
            .I(N__31682));
    LocalMux I__5982 (
            .O(N__31685),
            .I(N__31679));
    LocalMux I__5981 (
            .O(N__31682),
            .I(N__31676));
    Span4Mux_v I__5980 (
            .O(N__31679),
            .I(N__31673));
    Odrv4 I__5979 (
            .O(N__31676),
            .I(\nx.n2689 ));
    Odrv4 I__5978 (
            .O(N__31673),
            .I(\nx.n2689 ));
    CascadeMux I__5977 (
            .O(N__31668),
            .I(N__31664));
    CascadeMux I__5976 (
            .O(N__31667),
            .I(N__31661));
    InMux I__5975 (
            .O(N__31664),
            .I(N__31658));
    InMux I__5974 (
            .O(N__31661),
            .I(N__31655));
    LocalMux I__5973 (
            .O(N__31658),
            .I(N__31652));
    LocalMux I__5972 (
            .O(N__31655),
            .I(N__31649));
    Span4Mux_v I__5971 (
            .O(N__31652),
            .I(N__31645));
    Span4Mux_h I__5970 (
            .O(N__31649),
            .I(N__31642));
    InMux I__5969 (
            .O(N__31648),
            .I(N__31639));
    Odrv4 I__5968 (
            .O(N__31645),
            .I(\nx.n2690 ));
    Odrv4 I__5967 (
            .O(N__31642),
            .I(\nx.n2690 ));
    LocalMux I__5966 (
            .O(N__31639),
            .I(\nx.n2690 ));
    CascadeMux I__5965 (
            .O(N__31632),
            .I(\nx.n2689_cascade_ ));
    CascadeMux I__5964 (
            .O(N__31629),
            .I(N__31625));
    CascadeMux I__5963 (
            .O(N__31628),
            .I(N__31622));
    InMux I__5962 (
            .O(N__31625),
            .I(N__31619));
    InMux I__5961 (
            .O(N__31622),
            .I(N__31616));
    LocalMux I__5960 (
            .O(N__31619),
            .I(N__31611));
    LocalMux I__5959 (
            .O(N__31616),
            .I(N__31611));
    Span4Mux_v I__5958 (
            .O(N__31611),
            .I(N__31607));
    InMux I__5957 (
            .O(N__31610),
            .I(N__31604));
    Odrv4 I__5956 (
            .O(N__31607),
            .I(\nx.n2691 ));
    LocalMux I__5955 (
            .O(N__31604),
            .I(\nx.n2691 ));
    InMux I__5954 (
            .O(N__31599),
            .I(N__31595));
    CascadeMux I__5953 (
            .O(N__31598),
            .I(N__31592));
    LocalMux I__5952 (
            .O(N__31595),
            .I(N__31589));
    InMux I__5951 (
            .O(N__31592),
            .I(N__31586));
    Span4Mux_h I__5950 (
            .O(N__31589),
            .I(N__31580));
    LocalMux I__5949 (
            .O(N__31586),
            .I(N__31580));
    InMux I__5948 (
            .O(N__31585),
            .I(N__31577));
    Odrv4 I__5947 (
            .O(N__31580),
            .I(\nx.n2701 ));
    LocalMux I__5946 (
            .O(N__31577),
            .I(\nx.n2701 ));
    CascadeMux I__5945 (
            .O(N__31572),
            .I(\nx.n2105_cascade_ ));
    InMux I__5944 (
            .O(N__31569),
            .I(N__31565));
    CascadeMux I__5943 (
            .O(N__31568),
            .I(N__31561));
    LocalMux I__5942 (
            .O(N__31565),
            .I(N__31558));
    InMux I__5941 (
            .O(N__31564),
            .I(N__31555));
    InMux I__5940 (
            .O(N__31561),
            .I(N__31552));
    Span4Mux_v I__5939 (
            .O(N__31558),
            .I(N__31545));
    LocalMux I__5938 (
            .O(N__31555),
            .I(N__31545));
    LocalMux I__5937 (
            .O(N__31552),
            .I(N__31545));
    Odrv4 I__5936 (
            .O(N__31545),
            .I(\nx.n2704 ));
    CascadeMux I__5935 (
            .O(N__31542),
            .I(N__31539));
    InMux I__5934 (
            .O(N__31539),
            .I(N__31534));
    InMux I__5933 (
            .O(N__31538),
            .I(N__31529));
    InMux I__5932 (
            .O(N__31537),
            .I(N__31529));
    LocalMux I__5931 (
            .O(N__31534),
            .I(N__31526));
    LocalMux I__5930 (
            .O(N__31529),
            .I(N__31523));
    Span4Mux_v I__5929 (
            .O(N__31526),
            .I(N__31518));
    Span4Mux_h I__5928 (
            .O(N__31523),
            .I(N__31518));
    Odrv4 I__5927 (
            .O(N__31518),
            .I(\nx.n2695 ));
    CascadeMux I__5926 (
            .O(N__31515),
            .I(N__31512));
    InMux I__5925 (
            .O(N__31512),
            .I(N__31508));
    InMux I__5924 (
            .O(N__31511),
            .I(N__31505));
    LocalMux I__5923 (
            .O(N__31508),
            .I(N__31500));
    LocalMux I__5922 (
            .O(N__31505),
            .I(N__31500));
    Span4Mux_v I__5921 (
            .O(N__31500),
            .I(N__31497));
    Odrv4 I__5920 (
            .O(N__31497),
            .I(\nx.n2698 ));
    CascadeMux I__5919 (
            .O(N__31494),
            .I(\nx.n2698_cascade_ ));
    InMux I__5918 (
            .O(N__31491),
            .I(N__31488));
    LocalMux I__5917 (
            .O(N__31488),
            .I(N__31485));
    Odrv4 I__5916 (
            .O(N__31485),
            .I(\nx.n39_adj_610 ));
    InMux I__5915 (
            .O(N__31482),
            .I(N__31478));
    CascadeMux I__5914 (
            .O(N__31481),
            .I(N__31475));
    LocalMux I__5913 (
            .O(N__31478),
            .I(N__31471));
    InMux I__5912 (
            .O(N__31475),
            .I(N__31468));
    InMux I__5911 (
            .O(N__31474),
            .I(N__31465));
    Span4Mux_h I__5910 (
            .O(N__31471),
            .I(N__31460));
    LocalMux I__5909 (
            .O(N__31468),
            .I(N__31460));
    LocalMux I__5908 (
            .O(N__31465),
            .I(\nx.n2703 ));
    Odrv4 I__5907 (
            .O(N__31460),
            .I(\nx.n2703 ));
    InMux I__5906 (
            .O(N__31455),
            .I(N__31450));
    InMux I__5905 (
            .O(N__31454),
            .I(N__31447));
    CascadeMux I__5904 (
            .O(N__31453),
            .I(N__31444));
    LocalMux I__5903 (
            .O(N__31450),
            .I(N__31441));
    LocalMux I__5902 (
            .O(N__31447),
            .I(N__31438));
    InMux I__5901 (
            .O(N__31444),
            .I(N__31435));
    Span4Mux_v I__5900 (
            .O(N__31441),
            .I(N__31428));
    Span4Mux_h I__5899 (
            .O(N__31438),
            .I(N__31428));
    LocalMux I__5898 (
            .O(N__31435),
            .I(N__31428));
    Odrv4 I__5897 (
            .O(N__31428),
            .I(\nx.n2709 ));
    CascadeMux I__5896 (
            .O(N__31425),
            .I(\nx.n2592_cascade_ ));
    InMux I__5895 (
            .O(N__31422),
            .I(N__31419));
    LocalMux I__5894 (
            .O(N__31419),
            .I(N__31416));
    Span4Mux_h I__5893 (
            .O(N__31416),
            .I(N__31413));
    Odrv4 I__5892 (
            .O(N__31413),
            .I(n13146));
    CascadeMux I__5891 (
            .O(N__31410),
            .I(n13462_cascade_));
    InMux I__5890 (
            .O(N__31407),
            .I(N__31404));
    LocalMux I__5889 (
            .O(N__31404),
            .I(n13153));
    IoInMux I__5888 (
            .O(N__31401),
            .I(N__31398));
    LocalMux I__5887 (
            .O(N__31398),
            .I(N__31395));
    IoSpan4Mux I__5886 (
            .O(N__31395),
            .I(N__31392));
    Span4Mux_s3_h I__5885 (
            .O(N__31392),
            .I(N__31389));
    Span4Mux_h I__5884 (
            .O(N__31389),
            .I(N__31384));
    InMux I__5883 (
            .O(N__31388),
            .I(N__31379));
    InMux I__5882 (
            .O(N__31387),
            .I(N__31379));
    Odrv4 I__5881 (
            .O(N__31384),
            .I(pin_out_3));
    LocalMux I__5880 (
            .O(N__31379),
            .I(pin_out_3));
    IoInMux I__5879 (
            .O(N__31374),
            .I(N__31371));
    LocalMux I__5878 (
            .O(N__31371),
            .I(N__31368));
    IoSpan4Mux I__5877 (
            .O(N__31368),
            .I(N__31365));
    Span4Mux_s0_h I__5876 (
            .O(N__31365),
            .I(N__31362));
    Span4Mux_h I__5875 (
            .O(N__31362),
            .I(N__31357));
    InMux I__5874 (
            .O(N__31361),
            .I(N__31354));
    InMux I__5873 (
            .O(N__31360),
            .I(N__31351));
    Span4Mux_h I__5872 (
            .O(N__31357),
            .I(N__31346));
    LocalMux I__5871 (
            .O(N__31354),
            .I(N__31346));
    LocalMux I__5870 (
            .O(N__31351),
            .I(pin_out_2));
    Odrv4 I__5869 (
            .O(N__31346),
            .I(pin_out_2));
    InMux I__5868 (
            .O(N__31341),
            .I(N__31338));
    LocalMux I__5867 (
            .O(N__31338),
            .I(n13147));
    InMux I__5866 (
            .O(N__31335),
            .I(N__31332));
    LocalMux I__5865 (
            .O(N__31332),
            .I(n13168));
    CascadeMux I__5864 (
            .O(N__31329),
            .I(n13167_cascade_));
    InMux I__5863 (
            .O(N__31326),
            .I(N__31323));
    LocalMux I__5862 (
            .O(N__31323),
            .I(N__31320));
    Odrv12 I__5861 (
            .O(N__31320),
            .I(n13450));
    InMux I__5860 (
            .O(N__31317),
            .I(N__31313));
    InMux I__5859 (
            .O(N__31316),
            .I(N__31309));
    LocalMux I__5858 (
            .O(N__31313),
            .I(N__31306));
    InMux I__5857 (
            .O(N__31312),
            .I(N__31303));
    LocalMux I__5856 (
            .O(N__31309),
            .I(N__31300));
    Span4Mux_v I__5855 (
            .O(N__31306),
            .I(N__31295));
    LocalMux I__5854 (
            .O(N__31303),
            .I(N__31295));
    Span4Mux_v I__5853 (
            .O(N__31300),
            .I(N__31290));
    Span4Mux_h I__5852 (
            .O(N__31295),
            .I(N__31290));
    Odrv4 I__5851 (
            .O(N__31290),
            .I(\nx.n2694 ));
    CascadeMux I__5850 (
            .O(N__31287),
            .I(N__31283));
    CascadeMux I__5849 (
            .O(N__31286),
            .I(N__31279));
    InMux I__5848 (
            .O(N__31283),
            .I(N__31276));
    InMux I__5847 (
            .O(N__31282),
            .I(N__31271));
    InMux I__5846 (
            .O(N__31279),
            .I(N__31271));
    LocalMux I__5845 (
            .O(N__31276),
            .I(N__31268));
    LocalMux I__5844 (
            .O(N__31271),
            .I(N__31265));
    Span4Mux_h I__5843 (
            .O(N__31268),
            .I(N__31262));
    Odrv12 I__5842 (
            .O(N__31265),
            .I(\nx.n2697 ));
    Odrv4 I__5841 (
            .O(N__31262),
            .I(\nx.n2697 ));
    CascadeMux I__5840 (
            .O(N__31257),
            .I(n7258_cascade_));
    InMux I__5839 (
            .O(N__31254),
            .I(N__31251));
    LocalMux I__5838 (
            .O(N__31251),
            .I(N__31248));
    Odrv4 I__5837 (
            .O(N__31248),
            .I(n7236));
    CascadeMux I__5836 (
            .O(N__31245),
            .I(n7270_cascade_));
    InMux I__5835 (
            .O(N__31242),
            .I(N__31239));
    LocalMux I__5834 (
            .O(N__31239),
            .I(N__31236));
    Span4Mux_h I__5833 (
            .O(N__31236),
            .I(N__31233));
    Odrv4 I__5832 (
            .O(N__31233),
            .I(n7254));
    IoInMux I__5831 (
            .O(N__31230),
            .I(N__31227));
    LocalMux I__5830 (
            .O(N__31227),
            .I(N__31224));
    IoSpan4Mux I__5829 (
            .O(N__31224),
            .I(N__31221));
    Sp12to4 I__5828 (
            .O(N__31221),
            .I(N__31218));
    Span12Mux_s6_h I__5827 (
            .O(N__31218),
            .I(N__31215));
    Span12Mux_v I__5826 (
            .O(N__31215),
            .I(N__31210));
    InMux I__5825 (
            .O(N__31214),
            .I(N__31207));
    InMux I__5824 (
            .O(N__31213),
            .I(N__31204));
    Odrv12 I__5823 (
            .O(N__31210),
            .I(pin_out_5));
    LocalMux I__5822 (
            .O(N__31207),
            .I(pin_out_5));
    LocalMux I__5821 (
            .O(N__31204),
            .I(pin_out_5));
    CascadeMux I__5820 (
            .O(N__31197),
            .I(n13152_cascade_));
    InMux I__5819 (
            .O(N__31194),
            .I(\nx.n10608 ));
    CascadeMux I__5818 (
            .O(N__31191),
            .I(N__31188));
    InMux I__5817 (
            .O(N__31188),
            .I(N__31183));
    InMux I__5816 (
            .O(N__31187),
            .I(N__31178));
    InMux I__5815 (
            .O(N__31186),
            .I(N__31178));
    LocalMux I__5814 (
            .O(N__31183),
            .I(\nx.n1603 ));
    LocalMux I__5813 (
            .O(N__31178),
            .I(\nx.n1603 ));
    CascadeMux I__5812 (
            .O(N__31173),
            .I(N__31170));
    InMux I__5811 (
            .O(N__31170),
            .I(N__31167));
    LocalMux I__5810 (
            .O(N__31167),
            .I(\nx.n1670 ));
    InMux I__5809 (
            .O(N__31164),
            .I(\nx.n10609 ));
    CascadeMux I__5808 (
            .O(N__31161),
            .I(N__31157));
    CascadeMux I__5807 (
            .O(N__31160),
            .I(N__31153));
    InMux I__5806 (
            .O(N__31157),
            .I(N__31150));
    InMux I__5805 (
            .O(N__31156),
            .I(N__31147));
    InMux I__5804 (
            .O(N__31153),
            .I(N__31144));
    LocalMux I__5803 (
            .O(N__31150),
            .I(N__31141));
    LocalMux I__5802 (
            .O(N__31147),
            .I(N__31138));
    LocalMux I__5801 (
            .O(N__31144),
            .I(\nx.n1602 ));
    Odrv4 I__5800 (
            .O(N__31141),
            .I(\nx.n1602 ));
    Odrv4 I__5799 (
            .O(N__31138),
            .I(\nx.n1602 ));
    InMux I__5798 (
            .O(N__31131),
            .I(N__31128));
    LocalMux I__5797 (
            .O(N__31128),
            .I(N__31125));
    Odrv4 I__5796 (
            .O(N__31125),
            .I(\nx.n1669 ));
    InMux I__5795 (
            .O(N__31122),
            .I(bfn_7_31_0_));
    InMux I__5794 (
            .O(N__31119),
            .I(\nx.n10611 ));
    InMux I__5793 (
            .O(N__31116),
            .I(\nx.n10612 ));
    CascadeMux I__5792 (
            .O(N__31113),
            .I(N__31110));
    InMux I__5791 (
            .O(N__31110),
            .I(N__31106));
    InMux I__5790 (
            .O(N__31109),
            .I(N__31103));
    LocalMux I__5789 (
            .O(N__31106),
            .I(\nx.n1599 ));
    LocalMux I__5788 (
            .O(N__31103),
            .I(\nx.n1599 ));
    InMux I__5787 (
            .O(N__31098),
            .I(N__31095));
    LocalMux I__5786 (
            .O(N__31095),
            .I(\nx.n1666 ));
    InMux I__5785 (
            .O(N__31092),
            .I(\nx.n10613 ));
    InMux I__5784 (
            .O(N__31089),
            .I(N__31085));
    InMux I__5783 (
            .O(N__31088),
            .I(N__31082));
    LocalMux I__5782 (
            .O(N__31085),
            .I(N__31079));
    LocalMux I__5781 (
            .O(N__31082),
            .I(\nx.n1598 ));
    Odrv4 I__5780 (
            .O(N__31079),
            .I(\nx.n1598 ));
    InMux I__5779 (
            .O(N__31074),
            .I(\nx.n10614 ));
    CascadeMux I__5778 (
            .O(N__31071),
            .I(N__31066));
    CascadeMux I__5777 (
            .O(N__31070),
            .I(N__31063));
    InMux I__5776 (
            .O(N__31069),
            .I(N__31058));
    InMux I__5775 (
            .O(N__31066),
            .I(N__31058));
    InMux I__5774 (
            .O(N__31063),
            .I(N__31055));
    LocalMux I__5773 (
            .O(N__31058),
            .I(\nx.n1600 ));
    LocalMux I__5772 (
            .O(N__31055),
            .I(\nx.n1600 ));
    CascadeMux I__5771 (
            .O(N__31050),
            .I(N__31047));
    InMux I__5770 (
            .O(N__31047),
            .I(N__31044));
    LocalMux I__5769 (
            .O(N__31044),
            .I(\nx.n1667 ));
    InMux I__5768 (
            .O(N__31041),
            .I(N__31038));
    LocalMux I__5767 (
            .O(N__31038),
            .I(N__31035));
    Odrv4 I__5766 (
            .O(N__31035),
            .I(\nx.n1570 ));
    CascadeMux I__5765 (
            .O(N__31032),
            .I(N__31028));
    InMux I__5764 (
            .O(N__31031),
            .I(N__31025));
    InMux I__5763 (
            .O(N__31028),
            .I(N__31022));
    LocalMux I__5762 (
            .O(N__31025),
            .I(N__31017));
    LocalMux I__5761 (
            .O(N__31022),
            .I(N__31017));
    Span4Mux_v I__5760 (
            .O(N__31017),
            .I(N__31013));
    InMux I__5759 (
            .O(N__31016),
            .I(N__31010));
    Odrv4 I__5758 (
            .O(N__31013),
            .I(\nx.n1503 ));
    LocalMux I__5757 (
            .O(N__31010),
            .I(\nx.n1503 ));
    InMux I__5756 (
            .O(N__31005),
            .I(N__31000));
    InMux I__5755 (
            .O(N__31004),
            .I(N__30996));
    InMux I__5754 (
            .O(N__31003),
            .I(N__30992));
    LocalMux I__5753 (
            .O(N__31000),
            .I(N__30989));
    InMux I__5752 (
            .O(N__30999),
            .I(N__30986));
    LocalMux I__5751 (
            .O(N__30996),
            .I(N__30983));
    InMux I__5750 (
            .O(N__30995),
            .I(N__30980));
    LocalMux I__5749 (
            .O(N__30992),
            .I(N__30977));
    Span4Mux_h I__5748 (
            .O(N__30989),
            .I(N__30974));
    LocalMux I__5747 (
            .O(N__30986),
            .I(N__30971));
    Span4Mux_h I__5746 (
            .O(N__30983),
            .I(N__30968));
    LocalMux I__5745 (
            .O(N__30980),
            .I(\nx.bit_ctr_19 ));
    Odrv4 I__5744 (
            .O(N__30977),
            .I(\nx.bit_ctr_19 ));
    Odrv4 I__5743 (
            .O(N__30974),
            .I(\nx.bit_ctr_19 ));
    Odrv4 I__5742 (
            .O(N__30971),
            .I(\nx.bit_ctr_19 ));
    Odrv4 I__5741 (
            .O(N__30968),
            .I(\nx.bit_ctr_19 ));
    InMux I__5740 (
            .O(N__30957),
            .I(N__30954));
    LocalMux I__5739 (
            .O(N__30954),
            .I(N__30951));
    Span4Mux_h I__5738 (
            .O(N__30951),
            .I(N__30948));
    Odrv4 I__5737 (
            .O(N__30948),
            .I(\nx.n1677 ));
    InMux I__5736 (
            .O(N__30945),
            .I(bfn_7_30_0_));
    CascadeMux I__5735 (
            .O(N__30942),
            .I(N__30938));
    InMux I__5734 (
            .O(N__30941),
            .I(N__30935));
    InMux I__5733 (
            .O(N__30938),
            .I(N__30932));
    LocalMux I__5732 (
            .O(N__30935),
            .I(\nx.n1609 ));
    LocalMux I__5731 (
            .O(N__30932),
            .I(\nx.n1609 ));
    InMux I__5730 (
            .O(N__30927),
            .I(N__30924));
    LocalMux I__5729 (
            .O(N__30924),
            .I(\nx.n1676 ));
    InMux I__5728 (
            .O(N__30921),
            .I(\nx.n10603 ));
    InMux I__5727 (
            .O(N__30918),
            .I(\nx.n10604 ));
    CascadeMux I__5726 (
            .O(N__30915),
            .I(N__30911));
    CascadeMux I__5725 (
            .O(N__30914),
            .I(N__30907));
    InMux I__5724 (
            .O(N__30911),
            .I(N__30904));
    InMux I__5723 (
            .O(N__30910),
            .I(N__30901));
    InMux I__5722 (
            .O(N__30907),
            .I(N__30898));
    LocalMux I__5721 (
            .O(N__30904),
            .I(\nx.n1607 ));
    LocalMux I__5720 (
            .O(N__30901),
            .I(\nx.n1607 ));
    LocalMux I__5719 (
            .O(N__30898),
            .I(\nx.n1607 ));
    InMux I__5718 (
            .O(N__30891),
            .I(N__30888));
    LocalMux I__5717 (
            .O(N__30888),
            .I(N__30885));
    Odrv4 I__5716 (
            .O(N__30885),
            .I(\nx.n1674 ));
    InMux I__5715 (
            .O(N__30882),
            .I(\nx.n10605 ));
    InMux I__5714 (
            .O(N__30879),
            .I(\nx.n10606 ));
    InMux I__5713 (
            .O(N__30876),
            .I(N__30873));
    LocalMux I__5712 (
            .O(N__30873),
            .I(\nx.n1672 ));
    InMux I__5711 (
            .O(N__30870),
            .I(\nx.n10607 ));
    CascadeMux I__5710 (
            .O(N__30867),
            .I(\nx.n1701_cascade_ ));
    CascadeMux I__5709 (
            .O(N__30864),
            .I(\nx.n1801_cascade_ ));
    InMux I__5708 (
            .O(N__30861),
            .I(N__30858));
    LocalMux I__5707 (
            .O(N__30858),
            .I(\nx.n23 ));
    InMux I__5706 (
            .O(N__30855),
            .I(N__30852));
    LocalMux I__5705 (
            .O(N__30852),
            .I(N__30849));
    Odrv4 I__5704 (
            .O(N__30849),
            .I(\nx.n1577 ));
    InMux I__5703 (
            .O(N__30846),
            .I(N__30841));
    InMux I__5702 (
            .O(N__30845),
            .I(N__30838));
    InMux I__5701 (
            .O(N__30844),
            .I(N__30833));
    LocalMux I__5700 (
            .O(N__30841),
            .I(N__30828));
    LocalMux I__5699 (
            .O(N__30838),
            .I(N__30828));
    InMux I__5698 (
            .O(N__30837),
            .I(N__30825));
    InMux I__5697 (
            .O(N__30836),
            .I(N__30822));
    LocalMux I__5696 (
            .O(N__30833),
            .I(N__30819));
    Span4Mux_h I__5695 (
            .O(N__30828),
            .I(N__30816));
    LocalMux I__5694 (
            .O(N__30825),
            .I(N__30813));
    LocalMux I__5693 (
            .O(N__30822),
            .I(\nx.bit_ctr_20 ));
    Odrv4 I__5692 (
            .O(N__30819),
            .I(\nx.bit_ctr_20 ));
    Odrv4 I__5691 (
            .O(N__30816),
            .I(\nx.bit_ctr_20 ));
    Odrv12 I__5690 (
            .O(N__30813),
            .I(\nx.bit_ctr_20 ));
    CascadeMux I__5689 (
            .O(N__30804),
            .I(\nx.n1609_cascade_ ));
    InMux I__5688 (
            .O(N__30801),
            .I(N__30798));
    LocalMux I__5687 (
            .O(N__30798),
            .I(\nx.n16_adj_646 ));
    InMux I__5686 (
            .O(N__30795),
            .I(\nx.n10653 ));
    InMux I__5685 (
            .O(N__30792),
            .I(\nx.n10654 ));
    InMux I__5684 (
            .O(N__30789),
            .I(\nx.n10655 ));
    CascadeMux I__5683 (
            .O(N__30786),
            .I(N__30770));
    CascadeMux I__5682 (
            .O(N__30785),
            .I(N__30767));
    CascadeMux I__5681 (
            .O(N__30784),
            .I(N__30764));
    CascadeMux I__5680 (
            .O(N__30783),
            .I(N__30761));
    CascadeMux I__5679 (
            .O(N__30782),
            .I(N__30758));
    CascadeMux I__5678 (
            .O(N__30781),
            .I(N__30755));
    CascadeMux I__5677 (
            .O(N__30780),
            .I(N__30752));
    CascadeMux I__5676 (
            .O(N__30779),
            .I(N__30749));
    CascadeMux I__5675 (
            .O(N__30778),
            .I(N__30746));
    CascadeMux I__5674 (
            .O(N__30777),
            .I(N__30743));
    CascadeMux I__5673 (
            .O(N__30776),
            .I(N__30740));
    CascadeMux I__5672 (
            .O(N__30775),
            .I(N__30737));
    CascadeMux I__5671 (
            .O(N__30774),
            .I(N__30734));
    CascadeMux I__5670 (
            .O(N__30773),
            .I(N__30731));
    InMux I__5669 (
            .O(N__30770),
            .I(N__30722));
    InMux I__5668 (
            .O(N__30767),
            .I(N__30722));
    InMux I__5667 (
            .O(N__30764),
            .I(N__30722));
    InMux I__5666 (
            .O(N__30761),
            .I(N__30722));
    InMux I__5665 (
            .O(N__30758),
            .I(N__30713));
    InMux I__5664 (
            .O(N__30755),
            .I(N__30713));
    InMux I__5663 (
            .O(N__30752),
            .I(N__30713));
    InMux I__5662 (
            .O(N__30749),
            .I(N__30713));
    InMux I__5661 (
            .O(N__30746),
            .I(N__30706));
    InMux I__5660 (
            .O(N__30743),
            .I(N__30706));
    InMux I__5659 (
            .O(N__30740),
            .I(N__30706));
    InMux I__5658 (
            .O(N__30737),
            .I(N__30699));
    InMux I__5657 (
            .O(N__30734),
            .I(N__30699));
    InMux I__5656 (
            .O(N__30731),
            .I(N__30699));
    LocalMux I__5655 (
            .O(N__30722),
            .I(\nx.n1928 ));
    LocalMux I__5654 (
            .O(N__30713),
            .I(\nx.n1928 ));
    LocalMux I__5653 (
            .O(N__30706),
            .I(\nx.n1928 ));
    LocalMux I__5652 (
            .O(N__30699),
            .I(\nx.n1928 ));
    InMux I__5651 (
            .O(N__30690),
            .I(\nx.n10656 ));
    InMux I__5650 (
            .O(N__30687),
            .I(N__30682));
    InMux I__5649 (
            .O(N__30686),
            .I(N__30679));
    InMux I__5648 (
            .O(N__30685),
            .I(N__30676));
    LocalMux I__5647 (
            .O(N__30682),
            .I(N__30673));
    LocalMux I__5646 (
            .O(N__30679),
            .I(\nx.n1897 ));
    LocalMux I__5645 (
            .O(N__30676),
            .I(\nx.n1897 ));
    Odrv4 I__5644 (
            .O(N__30673),
            .I(\nx.n1897 ));
    InMux I__5643 (
            .O(N__30666),
            .I(N__30662));
    InMux I__5642 (
            .O(N__30665),
            .I(N__30659));
    LocalMux I__5641 (
            .O(N__30662),
            .I(N__30653));
    LocalMux I__5640 (
            .O(N__30659),
            .I(N__30653));
    InMux I__5639 (
            .O(N__30658),
            .I(N__30650));
    Odrv4 I__5638 (
            .O(N__30653),
            .I(\nx.n1902 ));
    LocalMux I__5637 (
            .O(N__30650),
            .I(\nx.n1902 ));
    CascadeMux I__5636 (
            .O(N__30645),
            .I(N__30640));
    InMux I__5635 (
            .O(N__30644),
            .I(N__30636));
    InMux I__5634 (
            .O(N__30643),
            .I(N__30633));
    InMux I__5633 (
            .O(N__30640),
            .I(N__30628));
    InMux I__5632 (
            .O(N__30639),
            .I(N__30628));
    LocalMux I__5631 (
            .O(N__30636),
            .I(N__30622));
    LocalMux I__5630 (
            .O(N__30633),
            .I(N__30619));
    LocalMux I__5629 (
            .O(N__30628),
            .I(N__30616));
    InMux I__5628 (
            .O(N__30627),
            .I(N__30609));
    InMux I__5627 (
            .O(N__30626),
            .I(N__30609));
    InMux I__5626 (
            .O(N__30625),
            .I(N__30609));
    Span4Mux_h I__5625 (
            .O(N__30622),
            .I(N__30606));
    Odrv4 I__5624 (
            .O(N__30619),
            .I(\nx.n10994 ));
    Odrv4 I__5623 (
            .O(N__30616),
            .I(\nx.n10994 ));
    LocalMux I__5622 (
            .O(N__30609),
            .I(\nx.n10994 ));
    Odrv4 I__5621 (
            .O(N__30606),
            .I(\nx.n10994 ));
    InMux I__5620 (
            .O(N__30597),
            .I(N__30594));
    LocalMux I__5619 (
            .O(N__30594),
            .I(\nx.n13425 ));
    InMux I__5618 (
            .O(N__30591),
            .I(N__30587));
    InMux I__5617 (
            .O(N__30590),
            .I(N__30584));
    LocalMux I__5616 (
            .O(N__30587),
            .I(\nx.n1906 ));
    LocalMux I__5615 (
            .O(N__30584),
            .I(\nx.n1906 ));
    InMux I__5614 (
            .O(N__30579),
            .I(\nx.n10645 ));
    InMux I__5613 (
            .O(N__30576),
            .I(\nx.n10646 ));
    CascadeMux I__5612 (
            .O(N__30573),
            .I(N__30568));
    InMux I__5611 (
            .O(N__30572),
            .I(N__30565));
    InMux I__5610 (
            .O(N__30571),
            .I(N__30562));
    InMux I__5609 (
            .O(N__30568),
            .I(N__30559));
    LocalMux I__5608 (
            .O(N__30565),
            .I(\nx.n1904 ));
    LocalMux I__5607 (
            .O(N__30562),
            .I(\nx.n1904 ));
    LocalMux I__5606 (
            .O(N__30559),
            .I(\nx.n1904 ));
    InMux I__5605 (
            .O(N__30552),
            .I(\nx.n10647 ));
    InMux I__5604 (
            .O(N__30549),
            .I(N__30544));
    InMux I__5603 (
            .O(N__30548),
            .I(N__30541));
    InMux I__5602 (
            .O(N__30547),
            .I(N__30538));
    LocalMux I__5601 (
            .O(N__30544),
            .I(\nx.n1903 ));
    LocalMux I__5600 (
            .O(N__30541),
            .I(\nx.n1903 ));
    LocalMux I__5599 (
            .O(N__30538),
            .I(\nx.n1903 ));
    InMux I__5598 (
            .O(N__30531),
            .I(\nx.n10648 ));
    InMux I__5597 (
            .O(N__30528),
            .I(bfn_7_26_0_));
    InMux I__5596 (
            .O(N__30525),
            .I(\nx.n10650 ));
    InMux I__5595 (
            .O(N__30522),
            .I(\nx.n10651 ));
    InMux I__5594 (
            .O(N__30519),
            .I(N__30514));
    InMux I__5593 (
            .O(N__30518),
            .I(N__30511));
    InMux I__5592 (
            .O(N__30517),
            .I(N__30508));
    LocalMux I__5591 (
            .O(N__30514),
            .I(N__30505));
    LocalMux I__5590 (
            .O(N__30511),
            .I(\nx.n1899 ));
    LocalMux I__5589 (
            .O(N__30508),
            .I(\nx.n1899 ));
    Odrv4 I__5588 (
            .O(N__30505),
            .I(\nx.n1899 ));
    InMux I__5587 (
            .O(N__30498),
            .I(\nx.n10652 ));
    CascadeMux I__5586 (
            .O(N__30495),
            .I(N__30492));
    InMux I__5585 (
            .O(N__30492),
            .I(N__30489));
    LocalMux I__5584 (
            .O(N__30489),
            .I(N__30485));
    CascadeMux I__5583 (
            .O(N__30488),
            .I(N__30482));
    Span4Mux_v I__5582 (
            .O(N__30485),
            .I(N__30478));
    InMux I__5581 (
            .O(N__30482),
            .I(N__30475));
    InMux I__5580 (
            .O(N__30481),
            .I(N__30472));
    Odrv4 I__5579 (
            .O(N__30478),
            .I(\nx.n2888 ));
    LocalMux I__5578 (
            .O(N__30475),
            .I(\nx.n2888 ));
    LocalMux I__5577 (
            .O(N__30472),
            .I(\nx.n2888 ));
    CascadeMux I__5576 (
            .O(N__30465),
            .I(\nx.n2887_cascade_ ));
    InMux I__5575 (
            .O(N__30462),
            .I(N__30459));
    LocalMux I__5574 (
            .O(N__30459),
            .I(N__30456));
    Span4Mux_h I__5573 (
            .O(N__30456),
            .I(N__30453));
    Odrv4 I__5572 (
            .O(N__30453),
            .I(\nx.n39_adj_679 ));
    InMux I__5571 (
            .O(N__30450),
            .I(N__30447));
    LocalMux I__5570 (
            .O(N__30447),
            .I(N__30443));
    CascadeMux I__5569 (
            .O(N__30446),
            .I(N__30439));
    Span4Mux_v I__5568 (
            .O(N__30443),
            .I(N__30436));
    InMux I__5567 (
            .O(N__30442),
            .I(N__30433));
    InMux I__5566 (
            .O(N__30439),
            .I(N__30430));
    Odrv4 I__5565 (
            .O(N__30436),
            .I(\nx.n2803 ));
    LocalMux I__5564 (
            .O(N__30433),
            .I(\nx.n2803 ));
    LocalMux I__5563 (
            .O(N__30430),
            .I(\nx.n2803 ));
    InMux I__5562 (
            .O(N__30423),
            .I(N__30420));
    LocalMux I__5561 (
            .O(N__30420),
            .I(N__30417));
    Span4Mux_h I__5560 (
            .O(N__30417),
            .I(N__30414));
    Odrv4 I__5559 (
            .O(N__30414),
            .I(\nx.n2870 ));
    InMux I__5558 (
            .O(N__30411),
            .I(N__30406));
    CascadeMux I__5557 (
            .O(N__30410),
            .I(N__30403));
    CascadeMux I__5556 (
            .O(N__30409),
            .I(N__30400));
    LocalMux I__5555 (
            .O(N__30406),
            .I(N__30397));
    InMux I__5554 (
            .O(N__30403),
            .I(N__30394));
    InMux I__5553 (
            .O(N__30400),
            .I(N__30391));
    Span4Mux_s2_h I__5552 (
            .O(N__30397),
            .I(N__30384));
    LocalMux I__5551 (
            .O(N__30394),
            .I(N__30384));
    LocalMux I__5550 (
            .O(N__30391),
            .I(N__30384));
    Span4Mux_h I__5549 (
            .O(N__30384),
            .I(N__30381));
    Odrv4 I__5548 (
            .O(N__30381),
            .I(\nx.n2902 ));
    InMux I__5547 (
            .O(N__30378),
            .I(N__30375));
    LocalMux I__5546 (
            .O(N__30375),
            .I(N__30372));
    Odrv4 I__5545 (
            .O(N__30372),
            .I(\nx.n2871 ));
    CascadeMux I__5544 (
            .O(N__30369),
            .I(N__30365));
    CascadeMux I__5543 (
            .O(N__30368),
            .I(N__30362));
    InMux I__5542 (
            .O(N__30365),
            .I(N__30358));
    InMux I__5541 (
            .O(N__30362),
            .I(N__30355));
    InMux I__5540 (
            .O(N__30361),
            .I(N__30352));
    LocalMux I__5539 (
            .O(N__30358),
            .I(N__30349));
    LocalMux I__5538 (
            .O(N__30355),
            .I(N__30346));
    LocalMux I__5537 (
            .O(N__30352),
            .I(N__30343));
    Span4Mux_h I__5536 (
            .O(N__30349),
            .I(N__30340));
    Span4Mux_h I__5535 (
            .O(N__30346),
            .I(N__30337));
    Odrv4 I__5534 (
            .O(N__30343),
            .I(\nx.n2903 ));
    Odrv4 I__5533 (
            .O(N__30340),
            .I(\nx.n2903 ));
    Odrv4 I__5532 (
            .O(N__30337),
            .I(\nx.n2903 ));
    InMux I__5531 (
            .O(N__30330),
            .I(N__30326));
    CascadeMux I__5530 (
            .O(N__30329),
            .I(N__30323));
    LocalMux I__5529 (
            .O(N__30326),
            .I(N__30319));
    InMux I__5528 (
            .O(N__30323),
            .I(N__30316));
    InMux I__5527 (
            .O(N__30322),
            .I(N__30313));
    Odrv4 I__5526 (
            .O(N__30319),
            .I(\nx.n2790 ));
    LocalMux I__5525 (
            .O(N__30316),
            .I(\nx.n2790 ));
    LocalMux I__5524 (
            .O(N__30313),
            .I(\nx.n2790 ));
    CascadeMux I__5523 (
            .O(N__30306),
            .I(N__30298));
    CascadeMux I__5522 (
            .O(N__30305),
            .I(N__30295));
    CascadeMux I__5521 (
            .O(N__30304),
            .I(N__30290));
    CascadeMux I__5520 (
            .O(N__30303),
            .I(N__30287));
    InMux I__5519 (
            .O(N__30302),
            .I(N__30278));
    InMux I__5518 (
            .O(N__30301),
            .I(N__30278));
    InMux I__5517 (
            .O(N__30298),
            .I(N__30263));
    InMux I__5516 (
            .O(N__30295),
            .I(N__30263));
    InMux I__5515 (
            .O(N__30294),
            .I(N__30263));
    InMux I__5514 (
            .O(N__30293),
            .I(N__30263));
    InMux I__5513 (
            .O(N__30290),
            .I(N__30263));
    InMux I__5512 (
            .O(N__30287),
            .I(N__30258));
    InMux I__5511 (
            .O(N__30286),
            .I(N__30258));
    CascadeMux I__5510 (
            .O(N__30285),
            .I(N__30252));
    CascadeMux I__5509 (
            .O(N__30284),
            .I(N__30247));
    CascadeMux I__5508 (
            .O(N__30283),
            .I(N__30243));
    LocalMux I__5507 (
            .O(N__30278),
            .I(N__30240));
    CascadeMux I__5506 (
            .O(N__30277),
            .I(N__30237));
    CascadeMux I__5505 (
            .O(N__30276),
            .I(N__30234));
    CascadeMux I__5504 (
            .O(N__30275),
            .I(N__30231));
    CascadeMux I__5503 (
            .O(N__30274),
            .I(N__30228));
    LocalMux I__5502 (
            .O(N__30263),
            .I(N__30224));
    LocalMux I__5501 (
            .O(N__30258),
            .I(N__30221));
    InMux I__5500 (
            .O(N__30257),
            .I(N__30218));
    CascadeMux I__5499 (
            .O(N__30256),
            .I(N__30215));
    CascadeMux I__5498 (
            .O(N__30255),
            .I(N__30212));
    InMux I__5497 (
            .O(N__30252),
            .I(N__30206));
    InMux I__5496 (
            .O(N__30251),
            .I(N__30206));
    InMux I__5495 (
            .O(N__30250),
            .I(N__30197));
    InMux I__5494 (
            .O(N__30247),
            .I(N__30197));
    InMux I__5493 (
            .O(N__30246),
            .I(N__30197));
    InMux I__5492 (
            .O(N__30243),
            .I(N__30197));
    Span4Mux_h I__5491 (
            .O(N__30240),
            .I(N__30194));
    InMux I__5490 (
            .O(N__30237),
            .I(N__30183));
    InMux I__5489 (
            .O(N__30234),
            .I(N__30183));
    InMux I__5488 (
            .O(N__30231),
            .I(N__30183));
    InMux I__5487 (
            .O(N__30228),
            .I(N__30183));
    InMux I__5486 (
            .O(N__30227),
            .I(N__30183));
    Span4Mux_v I__5485 (
            .O(N__30224),
            .I(N__30180));
    Span4Mux_h I__5484 (
            .O(N__30221),
            .I(N__30177));
    LocalMux I__5483 (
            .O(N__30218),
            .I(N__30174));
    InMux I__5482 (
            .O(N__30215),
            .I(N__30167));
    InMux I__5481 (
            .O(N__30212),
            .I(N__30167));
    InMux I__5480 (
            .O(N__30211),
            .I(N__30167));
    LocalMux I__5479 (
            .O(N__30206),
            .I(\nx.n2819 ));
    LocalMux I__5478 (
            .O(N__30197),
            .I(\nx.n2819 ));
    Odrv4 I__5477 (
            .O(N__30194),
            .I(\nx.n2819 ));
    LocalMux I__5476 (
            .O(N__30183),
            .I(\nx.n2819 ));
    Odrv4 I__5475 (
            .O(N__30180),
            .I(\nx.n2819 ));
    Odrv4 I__5474 (
            .O(N__30177),
            .I(\nx.n2819 ));
    Odrv12 I__5473 (
            .O(N__30174),
            .I(\nx.n2819 ));
    LocalMux I__5472 (
            .O(N__30167),
            .I(\nx.n2819 ));
    InMux I__5471 (
            .O(N__30150),
            .I(N__30147));
    LocalMux I__5470 (
            .O(N__30147),
            .I(\nx.n2857 ));
    InMux I__5469 (
            .O(N__30144),
            .I(N__30140));
    CascadeMux I__5468 (
            .O(N__30143),
            .I(N__30137));
    LocalMux I__5467 (
            .O(N__30140),
            .I(N__30134));
    InMux I__5466 (
            .O(N__30137),
            .I(N__30131));
    Span4Mux_v I__5465 (
            .O(N__30134),
            .I(N__30125));
    LocalMux I__5464 (
            .O(N__30131),
            .I(N__30125));
    InMux I__5463 (
            .O(N__30130),
            .I(N__30122));
    Odrv4 I__5462 (
            .O(N__30125),
            .I(\nx.n2889 ));
    LocalMux I__5461 (
            .O(N__30122),
            .I(\nx.n2889 ));
    InMux I__5460 (
            .O(N__30117),
            .I(N__30112));
    InMux I__5459 (
            .O(N__30116),
            .I(N__30109));
    CascadeMux I__5458 (
            .O(N__30115),
            .I(N__30105));
    LocalMux I__5457 (
            .O(N__30112),
            .I(N__30100));
    LocalMux I__5456 (
            .O(N__30109),
            .I(N__30100));
    InMux I__5455 (
            .O(N__30108),
            .I(N__30097));
    InMux I__5454 (
            .O(N__30105),
            .I(N__30093));
    Span4Mux_h I__5453 (
            .O(N__30100),
            .I(N__30090));
    LocalMux I__5452 (
            .O(N__30097),
            .I(N__30087));
    InMux I__5451 (
            .O(N__30096),
            .I(N__30084));
    LocalMux I__5450 (
            .O(N__30093),
            .I(N__30081));
    Span4Mux_s3_h I__5449 (
            .O(N__30090),
            .I(N__30078));
    Span4Mux_v I__5448 (
            .O(N__30087),
            .I(N__30075));
    LocalMux I__5447 (
            .O(N__30084),
            .I(\nx.bit_ctr_16 ));
    Odrv4 I__5446 (
            .O(N__30081),
            .I(\nx.bit_ctr_16 ));
    Odrv4 I__5445 (
            .O(N__30078),
            .I(\nx.bit_ctr_16 ));
    Odrv4 I__5444 (
            .O(N__30075),
            .I(\nx.bit_ctr_16 ));
    InMux I__5443 (
            .O(N__30066),
            .I(bfn_7_25_0_));
    InMux I__5442 (
            .O(N__30063),
            .I(N__30058));
    InMux I__5441 (
            .O(N__30062),
            .I(N__30055));
    InMux I__5440 (
            .O(N__30061),
            .I(N__30052));
    LocalMux I__5439 (
            .O(N__30058),
            .I(\nx.n1909 ));
    LocalMux I__5438 (
            .O(N__30055),
            .I(\nx.n1909 ));
    LocalMux I__5437 (
            .O(N__30052),
            .I(\nx.n1909 ));
    CascadeMux I__5436 (
            .O(N__30045),
            .I(N__30041));
    CascadeMux I__5435 (
            .O(N__30044),
            .I(N__30038));
    InMux I__5434 (
            .O(N__30041),
            .I(N__30035));
    InMux I__5433 (
            .O(N__30038),
            .I(N__30032));
    LocalMux I__5432 (
            .O(N__30035),
            .I(\nx.n13435 ));
    LocalMux I__5431 (
            .O(N__30032),
            .I(\nx.n13435 ));
    InMux I__5430 (
            .O(N__30027),
            .I(\nx.n10642 ));
    InMux I__5429 (
            .O(N__30024),
            .I(N__30020));
    InMux I__5428 (
            .O(N__30023),
            .I(N__30017));
    LocalMux I__5427 (
            .O(N__30020),
            .I(\nx.n1908 ));
    LocalMux I__5426 (
            .O(N__30017),
            .I(\nx.n1908 ));
    InMux I__5425 (
            .O(N__30012),
            .I(\nx.n10643 ));
    InMux I__5424 (
            .O(N__30009),
            .I(N__30004));
    InMux I__5423 (
            .O(N__30008),
            .I(N__30001));
    InMux I__5422 (
            .O(N__30007),
            .I(N__29998));
    LocalMux I__5421 (
            .O(N__30004),
            .I(\nx.n1907 ));
    LocalMux I__5420 (
            .O(N__30001),
            .I(\nx.n1907 ));
    LocalMux I__5419 (
            .O(N__29998),
            .I(\nx.n1907 ));
    InMux I__5418 (
            .O(N__29991),
            .I(\nx.n10644 ));
    InMux I__5417 (
            .O(N__29988),
            .I(N__29985));
    LocalMux I__5416 (
            .O(N__29985),
            .I(N__29982));
    Span4Mux_h I__5415 (
            .O(N__29982),
            .I(N__29979));
    Odrv4 I__5414 (
            .O(N__29979),
            .I(\nx.n44 ));
    InMux I__5413 (
            .O(N__29976),
            .I(N__29973));
    LocalMux I__5412 (
            .O(N__29973),
            .I(\nx.n2854 ));
    CascadeMux I__5411 (
            .O(N__29970),
            .I(\nx.n2819_cascade_ ));
    CascadeMux I__5410 (
            .O(N__29967),
            .I(N__29963));
    InMux I__5409 (
            .O(N__29966),
            .I(N__29960));
    InMux I__5408 (
            .O(N__29963),
            .I(N__29957));
    LocalMux I__5407 (
            .O(N__29960),
            .I(N__29953));
    LocalMux I__5406 (
            .O(N__29957),
            .I(N__29950));
    InMux I__5405 (
            .O(N__29956),
            .I(N__29947));
    Span4Mux_v I__5404 (
            .O(N__29953),
            .I(N__29944));
    Span4Mux_v I__5403 (
            .O(N__29950),
            .I(N__29939));
    LocalMux I__5402 (
            .O(N__29947),
            .I(N__29939));
    Odrv4 I__5401 (
            .O(N__29944),
            .I(\nx.n2886 ));
    Odrv4 I__5400 (
            .O(N__29939),
            .I(\nx.n2886 ));
    CascadeMux I__5399 (
            .O(N__29934),
            .I(N__29930));
    CascadeMux I__5398 (
            .O(N__29933),
            .I(N__29927));
    InMux I__5397 (
            .O(N__29930),
            .I(N__29924));
    InMux I__5396 (
            .O(N__29927),
            .I(N__29921));
    LocalMux I__5395 (
            .O(N__29924),
            .I(\nx.n2789 ));
    LocalMux I__5394 (
            .O(N__29921),
            .I(\nx.n2789 ));
    InMux I__5393 (
            .O(N__29916),
            .I(N__29913));
    LocalMux I__5392 (
            .O(N__29913),
            .I(\nx.n26_adj_615 ));
    InMux I__5391 (
            .O(N__29910),
            .I(N__29907));
    LocalMux I__5390 (
            .O(N__29907),
            .I(\nx.n2863 ));
    InMux I__5389 (
            .O(N__29904),
            .I(N__29900));
    CascadeMux I__5388 (
            .O(N__29903),
            .I(N__29897));
    LocalMux I__5387 (
            .O(N__29900),
            .I(N__29894));
    InMux I__5386 (
            .O(N__29897),
            .I(N__29891));
    Span4Mux_v I__5385 (
            .O(N__29894),
            .I(N__29887));
    LocalMux I__5384 (
            .O(N__29891),
            .I(N__29884));
    InMux I__5383 (
            .O(N__29890),
            .I(N__29881));
    Odrv4 I__5382 (
            .O(N__29887),
            .I(\nx.n2796 ));
    Odrv12 I__5381 (
            .O(N__29884),
            .I(\nx.n2796 ));
    LocalMux I__5380 (
            .O(N__29881),
            .I(\nx.n2796 ));
    InMux I__5379 (
            .O(N__29874),
            .I(N__29869));
    CascadeMux I__5378 (
            .O(N__29873),
            .I(N__29866));
    InMux I__5377 (
            .O(N__29872),
            .I(N__29863));
    LocalMux I__5376 (
            .O(N__29869),
            .I(N__29860));
    InMux I__5375 (
            .O(N__29866),
            .I(N__29857));
    LocalMux I__5374 (
            .O(N__29863),
            .I(N__29854));
    Span4Mux_v I__5373 (
            .O(N__29860),
            .I(N__29849));
    LocalMux I__5372 (
            .O(N__29857),
            .I(N__29849));
    Span4Mux_h I__5371 (
            .O(N__29854),
            .I(N__29846));
    Odrv4 I__5370 (
            .O(N__29849),
            .I(\nx.n2895 ));
    Odrv4 I__5369 (
            .O(N__29846),
            .I(\nx.n2895 ));
    InMux I__5368 (
            .O(N__29841),
            .I(N__29838));
    LocalMux I__5367 (
            .O(N__29838),
            .I(N__29835));
    Span4Mux_v I__5366 (
            .O(N__29835),
            .I(N__29832));
    Odrv4 I__5365 (
            .O(N__29832),
            .I(\nx.n2877 ));
    InMux I__5364 (
            .O(N__29829),
            .I(N__29823));
    InMux I__5363 (
            .O(N__29828),
            .I(N__29820));
    InMux I__5362 (
            .O(N__29827),
            .I(N__29817));
    InMux I__5361 (
            .O(N__29826),
            .I(N__29814));
    LocalMux I__5360 (
            .O(N__29823),
            .I(N__29809));
    LocalMux I__5359 (
            .O(N__29820),
            .I(N__29809));
    LocalMux I__5358 (
            .O(N__29817),
            .I(N__29805));
    LocalMux I__5357 (
            .O(N__29814),
            .I(N__29802));
    Span4Mux_v I__5356 (
            .O(N__29809),
            .I(N__29799));
    InMux I__5355 (
            .O(N__29808),
            .I(N__29796));
    Span12Mux_s5_v I__5354 (
            .O(N__29805),
            .I(N__29791));
    Span12Mux_v I__5353 (
            .O(N__29802),
            .I(N__29791));
    Span4Mux_v I__5352 (
            .O(N__29799),
            .I(N__29788));
    LocalMux I__5351 (
            .O(N__29796),
            .I(\nx.bit_ctr_7 ));
    Odrv12 I__5350 (
            .O(N__29791),
            .I(\nx.bit_ctr_7 ));
    Odrv4 I__5349 (
            .O(N__29788),
            .I(\nx.bit_ctr_7 ));
    CascadeMux I__5348 (
            .O(N__29781),
            .I(N__29778));
    InMux I__5347 (
            .O(N__29778),
            .I(N__29773));
    InMux I__5346 (
            .O(N__29777),
            .I(N__29770));
    InMux I__5345 (
            .O(N__29776),
            .I(N__29767));
    LocalMux I__5344 (
            .O(N__29773),
            .I(N__29764));
    LocalMux I__5343 (
            .O(N__29770),
            .I(N__29761));
    LocalMux I__5342 (
            .O(N__29767),
            .I(N__29758));
    Span4Mux_h I__5341 (
            .O(N__29764),
            .I(N__29755));
    Span4Mux_h I__5340 (
            .O(N__29761),
            .I(N__29752));
    Odrv12 I__5339 (
            .O(N__29758),
            .I(\nx.n2909 ));
    Odrv4 I__5338 (
            .O(N__29755),
            .I(\nx.n2909 ));
    Odrv4 I__5337 (
            .O(N__29752),
            .I(\nx.n2909 ));
    InMux I__5336 (
            .O(N__29745),
            .I(N__29742));
    LocalMux I__5335 (
            .O(N__29742),
            .I(\nx.n2868 ));
    InMux I__5334 (
            .O(N__29739),
            .I(N__29735));
    CascadeMux I__5333 (
            .O(N__29738),
            .I(N__29732));
    LocalMux I__5332 (
            .O(N__29735),
            .I(N__29729));
    InMux I__5331 (
            .O(N__29732),
            .I(N__29726));
    Span4Mux_v I__5330 (
            .O(N__29729),
            .I(N__29723));
    LocalMux I__5329 (
            .O(N__29726),
            .I(N__29720));
    Odrv4 I__5328 (
            .O(N__29723),
            .I(\nx.n2801 ));
    Odrv12 I__5327 (
            .O(N__29720),
            .I(\nx.n2801 ));
    InMux I__5326 (
            .O(N__29715),
            .I(N__29711));
    CascadeMux I__5325 (
            .O(N__29714),
            .I(N__29708));
    LocalMux I__5324 (
            .O(N__29711),
            .I(N__29704));
    InMux I__5323 (
            .O(N__29708),
            .I(N__29701));
    InMux I__5322 (
            .O(N__29707),
            .I(N__29698));
    Span4Mux_s3_h I__5321 (
            .O(N__29704),
            .I(N__29691));
    LocalMux I__5320 (
            .O(N__29701),
            .I(N__29691));
    LocalMux I__5319 (
            .O(N__29698),
            .I(N__29691));
    Odrv4 I__5318 (
            .O(N__29691),
            .I(\nx.n2900 ));
    InMux I__5317 (
            .O(N__29688),
            .I(N__29685));
    LocalMux I__5316 (
            .O(N__29685),
            .I(\nx.n2861 ));
    InMux I__5315 (
            .O(N__29682),
            .I(N__29678));
    CascadeMux I__5314 (
            .O(N__29681),
            .I(N__29675));
    LocalMux I__5313 (
            .O(N__29678),
            .I(N__29672));
    InMux I__5312 (
            .O(N__29675),
            .I(N__29669));
    Span4Mux_v I__5311 (
            .O(N__29672),
            .I(N__29665));
    LocalMux I__5310 (
            .O(N__29669),
            .I(N__29662));
    InMux I__5309 (
            .O(N__29668),
            .I(N__29659));
    Odrv4 I__5308 (
            .O(N__29665),
            .I(\nx.n2794 ));
    Odrv12 I__5307 (
            .O(N__29662),
            .I(\nx.n2794 ));
    LocalMux I__5306 (
            .O(N__29659),
            .I(\nx.n2794 ));
    InMux I__5305 (
            .O(N__29652),
            .I(N__29647));
    CascadeMux I__5304 (
            .O(N__29651),
            .I(N__29644));
    InMux I__5303 (
            .O(N__29650),
            .I(N__29641));
    LocalMux I__5302 (
            .O(N__29647),
            .I(N__29638));
    InMux I__5301 (
            .O(N__29644),
            .I(N__29635));
    LocalMux I__5300 (
            .O(N__29641),
            .I(N__29632));
    Span4Mux_v I__5299 (
            .O(N__29638),
            .I(N__29627));
    LocalMux I__5298 (
            .O(N__29635),
            .I(N__29627));
    Span4Mux_h I__5297 (
            .O(N__29632),
            .I(N__29624));
    Odrv4 I__5296 (
            .O(N__29627),
            .I(\nx.n2893 ));
    Odrv4 I__5295 (
            .O(N__29624),
            .I(\nx.n2893 ));
    InMux I__5294 (
            .O(N__29619),
            .I(N__29614));
    InMux I__5293 (
            .O(N__29618),
            .I(N__29611));
    InMux I__5292 (
            .O(N__29617),
            .I(N__29608));
    LocalMux I__5291 (
            .O(N__29614),
            .I(N__29601));
    LocalMux I__5290 (
            .O(N__29611),
            .I(N__29601));
    LocalMux I__5289 (
            .O(N__29608),
            .I(N__29601));
    Span4Mux_v I__5288 (
            .O(N__29601),
            .I(N__29598));
    Odrv4 I__5287 (
            .O(N__29598),
            .I(\nx.n2788 ));
    InMux I__5286 (
            .O(N__29595),
            .I(N__29592));
    LocalMux I__5285 (
            .O(N__29592),
            .I(\nx.n2855 ));
    InMux I__5284 (
            .O(N__29589),
            .I(N__29586));
    LocalMux I__5283 (
            .O(N__29586),
            .I(N__29582));
    InMux I__5282 (
            .O(N__29585),
            .I(N__29579));
    Span4Mux_v I__5281 (
            .O(N__29582),
            .I(N__29574));
    LocalMux I__5280 (
            .O(N__29579),
            .I(N__29574));
    Odrv4 I__5279 (
            .O(N__29574),
            .I(\nx.n2887 ));
    InMux I__5278 (
            .O(N__29571),
            .I(N__29567));
    CascadeMux I__5277 (
            .O(N__29570),
            .I(N__29564));
    LocalMux I__5276 (
            .O(N__29567),
            .I(N__29560));
    InMux I__5275 (
            .O(N__29564),
            .I(N__29557));
    InMux I__5274 (
            .O(N__29563),
            .I(N__29554));
    Odrv4 I__5273 (
            .O(N__29560),
            .I(\nx.n2890 ));
    LocalMux I__5272 (
            .O(N__29557),
            .I(\nx.n2890 ));
    LocalMux I__5271 (
            .O(N__29554),
            .I(\nx.n2890 ));
    CascadeMux I__5270 (
            .O(N__29547),
            .I(N__29544));
    InMux I__5269 (
            .O(N__29544),
            .I(N__29541));
    LocalMux I__5268 (
            .O(N__29541),
            .I(\nx.n2761 ));
    InMux I__5267 (
            .O(N__29538),
            .I(N__29535));
    LocalMux I__5266 (
            .O(N__29535),
            .I(\nx.n2860 ));
    CascadeMux I__5265 (
            .O(N__29532),
            .I(\nx.n2793_cascade_ ));
    CascadeMux I__5264 (
            .O(N__29529),
            .I(N__29525));
    InMux I__5263 (
            .O(N__29528),
            .I(N__29522));
    InMux I__5262 (
            .O(N__29525),
            .I(N__29519));
    LocalMux I__5261 (
            .O(N__29522),
            .I(N__29515));
    LocalMux I__5260 (
            .O(N__29519),
            .I(N__29512));
    InMux I__5259 (
            .O(N__29518),
            .I(N__29509));
    Span4Mux_h I__5258 (
            .O(N__29515),
            .I(N__29506));
    Span4Mux_v I__5257 (
            .O(N__29512),
            .I(N__29503));
    LocalMux I__5256 (
            .O(N__29509),
            .I(N__29500));
    Odrv4 I__5255 (
            .O(N__29506),
            .I(\nx.n2892 ));
    Odrv4 I__5254 (
            .O(N__29503),
            .I(\nx.n2892 ));
    Odrv4 I__5253 (
            .O(N__29500),
            .I(\nx.n2892 ));
    InMux I__5252 (
            .O(N__29493),
            .I(N__29490));
    LocalMux I__5251 (
            .O(N__29490),
            .I(\nx.n2758 ));
    InMux I__5250 (
            .O(N__29487),
            .I(N__29484));
    LocalMux I__5249 (
            .O(N__29484),
            .I(\nx.n2760 ));
    InMux I__5248 (
            .O(N__29481),
            .I(N__29478));
    LocalMux I__5247 (
            .O(N__29478),
            .I(\nx.n2873 ));
    InMux I__5246 (
            .O(N__29475),
            .I(N__29471));
    CascadeMux I__5245 (
            .O(N__29474),
            .I(N__29467));
    LocalMux I__5244 (
            .O(N__29471),
            .I(N__29464));
    InMux I__5243 (
            .O(N__29470),
            .I(N__29461));
    InMux I__5242 (
            .O(N__29467),
            .I(N__29458));
    Odrv4 I__5241 (
            .O(N__29464),
            .I(\nx.n2806 ));
    LocalMux I__5240 (
            .O(N__29461),
            .I(\nx.n2806 ));
    LocalMux I__5239 (
            .O(N__29458),
            .I(\nx.n2806 ));
    InMux I__5238 (
            .O(N__29451),
            .I(N__29447));
    InMux I__5237 (
            .O(N__29450),
            .I(N__29444));
    LocalMux I__5236 (
            .O(N__29447),
            .I(N__29438));
    LocalMux I__5235 (
            .O(N__29444),
            .I(N__29438));
    InMux I__5234 (
            .O(N__29443),
            .I(N__29435));
    Span4Mux_v I__5233 (
            .O(N__29438),
            .I(N__29430));
    LocalMux I__5232 (
            .O(N__29435),
            .I(N__29430));
    Odrv4 I__5231 (
            .O(N__29430),
            .I(\nx.n2905 ));
    CascadeMux I__5230 (
            .O(N__29427),
            .I(N__29424));
    InMux I__5229 (
            .O(N__29424),
            .I(N__29420));
    InMux I__5228 (
            .O(N__29423),
            .I(N__29417));
    LocalMux I__5227 (
            .O(N__29420),
            .I(\nx.n2793 ));
    LocalMux I__5226 (
            .O(N__29417),
            .I(\nx.n2793 ));
    CascadeMux I__5225 (
            .O(N__29412),
            .I(N__29409));
    InMux I__5224 (
            .O(N__29409),
            .I(N__29405));
    InMux I__5223 (
            .O(N__29408),
            .I(N__29402));
    LocalMux I__5222 (
            .O(N__29405),
            .I(\nx.n2791 ));
    LocalMux I__5221 (
            .O(N__29402),
            .I(\nx.n2791 ));
    InMux I__5220 (
            .O(N__29397),
            .I(N__29392));
    CascadeMux I__5219 (
            .O(N__29396),
            .I(N__29389));
    CascadeMux I__5218 (
            .O(N__29395),
            .I(N__29386));
    LocalMux I__5217 (
            .O(N__29392),
            .I(N__29383));
    InMux I__5216 (
            .O(N__29389),
            .I(N__29380));
    InMux I__5215 (
            .O(N__29386),
            .I(N__29377));
    Odrv4 I__5214 (
            .O(N__29383),
            .I(\nx.n2792 ));
    LocalMux I__5213 (
            .O(N__29380),
            .I(\nx.n2792 ));
    LocalMux I__5212 (
            .O(N__29377),
            .I(\nx.n2792 ));
    InMux I__5211 (
            .O(N__29370),
            .I(N__29366));
    InMux I__5210 (
            .O(N__29369),
            .I(N__29363));
    LocalMux I__5209 (
            .O(N__29366),
            .I(N__29358));
    LocalMux I__5208 (
            .O(N__29363),
            .I(N__29358));
    Odrv4 I__5207 (
            .O(N__29358),
            .I(\nx.n2786 ));
    CascadeMux I__5206 (
            .O(N__29355),
            .I(\nx.n38_adj_625_cascade_ ));
    InMux I__5205 (
            .O(N__29352),
            .I(N__29349));
    LocalMux I__5204 (
            .O(N__29349),
            .I(N__29346));
    Span4Mux_v I__5203 (
            .O(N__29346),
            .I(N__29343));
    Odrv4 I__5202 (
            .O(N__29343),
            .I(\nx.n42_adj_635 ));
    InMux I__5201 (
            .O(N__29340),
            .I(N__29337));
    LocalMux I__5200 (
            .O(N__29337),
            .I(N__29334));
    Odrv4 I__5199 (
            .O(N__29334),
            .I(\nx.n41_adj_643 ));
    CascadeMux I__5198 (
            .O(N__29331),
            .I(\nx.n43_cascade_ ));
    InMux I__5197 (
            .O(N__29328),
            .I(\nx.n10806 ));
    InMux I__5196 (
            .O(N__29325),
            .I(N__29322));
    LocalMux I__5195 (
            .O(N__29322),
            .I(N__29319));
    Odrv4 I__5194 (
            .O(N__29319),
            .I(\nx.n2759 ));
    InMux I__5193 (
            .O(N__29316),
            .I(\nx.n10807 ));
    InMux I__5192 (
            .O(N__29313),
            .I(\nx.n10808 ));
    InMux I__5191 (
            .O(N__29310),
            .I(N__29307));
    LocalMux I__5190 (
            .O(N__29307),
            .I(N__29304));
    Odrv4 I__5189 (
            .O(N__29304),
            .I(\nx.n2757 ));
    InMux I__5188 (
            .O(N__29301),
            .I(\nx.n10809 ));
    InMux I__5187 (
            .O(N__29298),
            .I(N__29295));
    LocalMux I__5186 (
            .O(N__29295),
            .I(\nx.n2756 ));
    InMux I__5185 (
            .O(N__29292),
            .I(\nx.n10810 ));
    InMux I__5184 (
            .O(N__29289),
            .I(\nx.n10811 ));
    InMux I__5183 (
            .O(N__29286),
            .I(\nx.n10812 ));
    InMux I__5182 (
            .O(N__29283),
            .I(N__29280));
    LocalMux I__5181 (
            .O(N__29280),
            .I(N__29277));
    Span4Mux_v I__5180 (
            .O(N__29277),
            .I(N__29273));
    InMux I__5179 (
            .O(N__29276),
            .I(N__29270));
    Span4Mux_v I__5178 (
            .O(N__29273),
            .I(N__29267));
    LocalMux I__5177 (
            .O(N__29270),
            .I(neo_pixel_transmitter_t0_22));
    Odrv4 I__5176 (
            .O(N__29267),
            .I(neo_pixel_transmitter_t0_22));
    CascadeMux I__5175 (
            .O(N__29262),
            .I(N__29259));
    InMux I__5174 (
            .O(N__29259),
            .I(N__29256));
    LocalMux I__5173 (
            .O(N__29256),
            .I(N__29253));
    Span4Mux_v I__5172 (
            .O(N__29253),
            .I(N__29250));
    Span4Mux_h I__5171 (
            .O(N__29250),
            .I(N__29247));
    Odrv4 I__5170 (
            .O(N__29247),
            .I(\nx.n11 ));
    InMux I__5169 (
            .O(N__29244),
            .I(N__29241));
    LocalMux I__5168 (
            .O(N__29241),
            .I(N__29238));
    Odrv4 I__5167 (
            .O(N__29238),
            .I(\nx.n2768 ));
    InMux I__5166 (
            .O(N__29235),
            .I(\nx.n10798 ));
    CascadeMux I__5165 (
            .O(N__29232),
            .I(N__29228));
    CascadeMux I__5164 (
            .O(N__29231),
            .I(N__29225));
    InMux I__5163 (
            .O(N__29228),
            .I(N__29222));
    InMux I__5162 (
            .O(N__29225),
            .I(N__29219));
    LocalMux I__5161 (
            .O(N__29222),
            .I(N__29214));
    LocalMux I__5160 (
            .O(N__29219),
            .I(N__29214));
    Odrv4 I__5159 (
            .O(N__29214),
            .I(\nx.n2700 ));
    InMux I__5158 (
            .O(N__29211),
            .I(N__29208));
    LocalMux I__5157 (
            .O(N__29208),
            .I(\nx.n2767 ));
    InMux I__5156 (
            .O(N__29205),
            .I(\nx.n10799 ));
    InMux I__5155 (
            .O(N__29202),
            .I(N__29199));
    LocalMux I__5154 (
            .O(N__29199),
            .I(\nx.n2766 ));
    InMux I__5153 (
            .O(N__29196),
            .I(\nx.n10800 ));
    InMux I__5152 (
            .O(N__29193),
            .I(N__29190));
    LocalMux I__5151 (
            .O(N__29190),
            .I(\nx.n2765 ));
    InMux I__5150 (
            .O(N__29187),
            .I(\nx.n10801 ));
    CascadeMux I__5149 (
            .O(N__29184),
            .I(N__29181));
    InMux I__5148 (
            .O(N__29181),
            .I(N__29178));
    LocalMux I__5147 (
            .O(N__29178),
            .I(\nx.n2764 ));
    InMux I__5146 (
            .O(N__29175),
            .I(\nx.n10802 ));
    CascadeMux I__5145 (
            .O(N__29172),
            .I(N__29168));
    InMux I__5144 (
            .O(N__29171),
            .I(N__29164));
    InMux I__5143 (
            .O(N__29168),
            .I(N__29161));
    InMux I__5142 (
            .O(N__29167),
            .I(N__29158));
    LocalMux I__5141 (
            .O(N__29164),
            .I(N__29153));
    LocalMux I__5140 (
            .O(N__29161),
            .I(N__29153));
    LocalMux I__5139 (
            .O(N__29158),
            .I(N__29150));
    Span4Mux_h I__5138 (
            .O(N__29153),
            .I(N__29147));
    Odrv12 I__5137 (
            .O(N__29150),
            .I(\nx.n2696 ));
    Odrv4 I__5136 (
            .O(N__29147),
            .I(\nx.n2696 ));
    CascadeMux I__5135 (
            .O(N__29142),
            .I(N__29139));
    InMux I__5134 (
            .O(N__29139),
            .I(N__29136));
    LocalMux I__5133 (
            .O(N__29136),
            .I(\nx.n2763 ));
    InMux I__5132 (
            .O(N__29133),
            .I(\nx.n10803 ));
    InMux I__5131 (
            .O(N__29130),
            .I(N__29127));
    LocalMux I__5130 (
            .O(N__29127),
            .I(\nx.n2762 ));
    InMux I__5129 (
            .O(N__29124),
            .I(\nx.n10804 ));
    InMux I__5128 (
            .O(N__29121),
            .I(bfn_7_21_0_));
    CascadeMux I__5127 (
            .O(N__29118),
            .I(N__29115));
    InMux I__5126 (
            .O(N__29115),
            .I(N__29112));
    LocalMux I__5125 (
            .O(N__29112),
            .I(\nx.n2776 ));
    InMux I__5124 (
            .O(N__29109),
            .I(\nx.n10790 ));
    CascadeMux I__5123 (
            .O(N__29106),
            .I(N__29102));
    CascadeMux I__5122 (
            .O(N__29105),
            .I(N__29098));
    InMux I__5121 (
            .O(N__29102),
            .I(N__29095));
    InMux I__5120 (
            .O(N__29101),
            .I(N__29092));
    InMux I__5119 (
            .O(N__29098),
            .I(N__29089));
    LocalMux I__5118 (
            .O(N__29095),
            .I(\nx.n2708 ));
    LocalMux I__5117 (
            .O(N__29092),
            .I(\nx.n2708 ));
    LocalMux I__5116 (
            .O(N__29089),
            .I(\nx.n2708 ));
    InMux I__5115 (
            .O(N__29082),
            .I(N__29079));
    LocalMux I__5114 (
            .O(N__29079),
            .I(\nx.n2775 ));
    InMux I__5113 (
            .O(N__29076),
            .I(\nx.n10791 ));
    CascadeMux I__5112 (
            .O(N__29073),
            .I(N__29070));
    InMux I__5111 (
            .O(N__29070),
            .I(N__29065));
    CascadeMux I__5110 (
            .O(N__29069),
            .I(N__29062));
    CascadeMux I__5109 (
            .O(N__29068),
            .I(N__29059));
    LocalMux I__5108 (
            .O(N__29065),
            .I(N__29056));
    InMux I__5107 (
            .O(N__29062),
            .I(N__29053));
    InMux I__5106 (
            .O(N__29059),
            .I(N__29050));
    Odrv4 I__5105 (
            .O(N__29056),
            .I(\nx.n2707 ));
    LocalMux I__5104 (
            .O(N__29053),
            .I(\nx.n2707 ));
    LocalMux I__5103 (
            .O(N__29050),
            .I(\nx.n2707 ));
    InMux I__5102 (
            .O(N__29043),
            .I(N__29040));
    LocalMux I__5101 (
            .O(N__29040),
            .I(\nx.n2774 ));
    InMux I__5100 (
            .O(N__29037),
            .I(\nx.n10792 ));
    CascadeMux I__5099 (
            .O(N__29034),
            .I(N__29029));
    InMux I__5098 (
            .O(N__29033),
            .I(N__29026));
    InMux I__5097 (
            .O(N__29032),
            .I(N__29023));
    InMux I__5096 (
            .O(N__29029),
            .I(N__29020));
    LocalMux I__5095 (
            .O(N__29026),
            .I(\nx.n2706 ));
    LocalMux I__5094 (
            .O(N__29023),
            .I(\nx.n2706 ));
    LocalMux I__5093 (
            .O(N__29020),
            .I(\nx.n2706 ));
    CascadeMux I__5092 (
            .O(N__29013),
            .I(N__29010));
    InMux I__5091 (
            .O(N__29010),
            .I(N__29007));
    LocalMux I__5090 (
            .O(N__29007),
            .I(N__29004));
    Odrv4 I__5089 (
            .O(N__29004),
            .I(\nx.n2773 ));
    InMux I__5088 (
            .O(N__29001),
            .I(\nx.n10793 ));
    InMux I__5087 (
            .O(N__28998),
            .I(\nx.n10794 ));
    InMux I__5086 (
            .O(N__28995),
            .I(N__28992));
    LocalMux I__5085 (
            .O(N__28992),
            .I(\nx.n2771 ));
    InMux I__5084 (
            .O(N__28989),
            .I(\nx.n10795 ));
    InMux I__5083 (
            .O(N__28986),
            .I(N__28983));
    LocalMux I__5082 (
            .O(N__28983),
            .I(\nx.n2770 ));
    InMux I__5081 (
            .O(N__28980),
            .I(\nx.n10796 ));
    CascadeMux I__5080 (
            .O(N__28977),
            .I(N__28973));
    CascadeMux I__5079 (
            .O(N__28976),
            .I(N__28970));
    InMux I__5078 (
            .O(N__28973),
            .I(N__28966));
    InMux I__5077 (
            .O(N__28970),
            .I(N__28961));
    InMux I__5076 (
            .O(N__28969),
            .I(N__28961));
    LocalMux I__5075 (
            .O(N__28966),
            .I(N__28958));
    LocalMux I__5074 (
            .O(N__28961),
            .I(\nx.n2702 ));
    Odrv12 I__5073 (
            .O(N__28958),
            .I(\nx.n2702 ));
    InMux I__5072 (
            .O(N__28953),
            .I(N__28950));
    LocalMux I__5071 (
            .O(N__28950),
            .I(N__28947));
    Odrv4 I__5070 (
            .O(N__28947),
            .I(\nx.n2769 ));
    InMux I__5069 (
            .O(N__28944),
            .I(bfn_7_20_0_));
    InMux I__5068 (
            .O(N__28941),
            .I(N__28938));
    LocalMux I__5067 (
            .O(N__28938),
            .I(N__28934));
    InMux I__5066 (
            .O(N__28937),
            .I(N__28931));
    Span4Mux_s1_v I__5065 (
            .O(N__28934),
            .I(N__28926));
    LocalMux I__5064 (
            .O(N__28931),
            .I(N__28926));
    Span4Mux_h I__5063 (
            .O(N__28926),
            .I(N__28923));
    Odrv4 I__5062 (
            .O(N__28923),
            .I(\nx.n1499 ));
    InMux I__5061 (
            .O(N__28920),
            .I(\nx.n10602 ));
    InMux I__5060 (
            .O(N__28917),
            .I(N__28912));
    InMux I__5059 (
            .O(N__28916),
            .I(N__28909));
    InMux I__5058 (
            .O(N__28915),
            .I(N__28906));
    LocalMux I__5057 (
            .O(N__28912),
            .I(N__28901));
    LocalMux I__5056 (
            .O(N__28909),
            .I(N__28901));
    LocalMux I__5055 (
            .O(N__28906),
            .I(N__28898));
    Span4Mux_v I__5054 (
            .O(N__28901),
            .I(N__28894));
    Span4Mux_h I__5053 (
            .O(N__28898),
            .I(N__28891));
    InMux I__5052 (
            .O(N__28897),
            .I(N__28888));
    Span4Mux_h I__5051 (
            .O(N__28894),
            .I(N__28885));
    Odrv4 I__5050 (
            .O(N__28891),
            .I(neopxl_color_13));
    LocalMux I__5049 (
            .O(N__28888),
            .I(neopxl_color_13));
    Odrv4 I__5048 (
            .O(N__28885),
            .I(neopxl_color_13));
    InMux I__5047 (
            .O(N__28878),
            .I(N__28870));
    InMux I__5046 (
            .O(N__28877),
            .I(N__28867));
    InMux I__5045 (
            .O(N__28876),
            .I(N__28859));
    CascadeMux I__5044 (
            .O(N__28875),
            .I(N__28852));
    InMux I__5043 (
            .O(N__28874),
            .I(N__28847));
    CascadeMux I__5042 (
            .O(N__28873),
            .I(N__28844));
    LocalMux I__5041 (
            .O(N__28870),
            .I(N__28828));
    LocalMux I__5040 (
            .O(N__28867),
            .I(N__28828));
    InMux I__5039 (
            .O(N__28866),
            .I(N__28825));
    InMux I__5038 (
            .O(N__28865),
            .I(N__28822));
    InMux I__5037 (
            .O(N__28864),
            .I(N__28815));
    InMux I__5036 (
            .O(N__28863),
            .I(N__28815));
    InMux I__5035 (
            .O(N__28862),
            .I(N__28815));
    LocalMux I__5034 (
            .O(N__28859),
            .I(N__28812));
    InMux I__5033 (
            .O(N__28858),
            .I(N__28807));
    InMux I__5032 (
            .O(N__28857),
            .I(N__28807));
    InMux I__5031 (
            .O(N__28856),
            .I(N__28802));
    InMux I__5030 (
            .O(N__28855),
            .I(N__28802));
    InMux I__5029 (
            .O(N__28852),
            .I(N__28797));
    InMux I__5028 (
            .O(N__28851),
            .I(N__28797));
    InMux I__5027 (
            .O(N__28850),
            .I(N__28794));
    LocalMux I__5026 (
            .O(N__28847),
            .I(N__28791));
    InMux I__5025 (
            .O(N__28844),
            .I(N__28786));
    InMux I__5024 (
            .O(N__28843),
            .I(N__28786));
    InMux I__5023 (
            .O(N__28842),
            .I(N__28783));
    InMux I__5022 (
            .O(N__28841),
            .I(N__28778));
    InMux I__5021 (
            .O(N__28840),
            .I(N__28778));
    InMux I__5020 (
            .O(N__28839),
            .I(N__28769));
    InMux I__5019 (
            .O(N__28838),
            .I(N__28769));
    InMux I__5018 (
            .O(N__28837),
            .I(N__28764));
    InMux I__5017 (
            .O(N__28836),
            .I(N__28764));
    InMux I__5016 (
            .O(N__28835),
            .I(N__28757));
    InMux I__5015 (
            .O(N__28834),
            .I(N__28757));
    InMux I__5014 (
            .O(N__28833),
            .I(N__28757));
    Span4Mux_v I__5013 (
            .O(N__28828),
            .I(N__28750));
    LocalMux I__5012 (
            .O(N__28825),
            .I(N__28750));
    LocalMux I__5011 (
            .O(N__28822),
            .I(N__28750));
    LocalMux I__5010 (
            .O(N__28815),
            .I(N__28745));
    Span4Mux_h I__5009 (
            .O(N__28812),
            .I(N__28745));
    LocalMux I__5008 (
            .O(N__28807),
            .I(N__28742));
    LocalMux I__5007 (
            .O(N__28802),
            .I(N__28735));
    LocalMux I__5006 (
            .O(N__28797),
            .I(N__28735));
    LocalMux I__5005 (
            .O(N__28794),
            .I(N__28735));
    Span4Mux_v I__5004 (
            .O(N__28791),
            .I(N__28732));
    LocalMux I__5003 (
            .O(N__28786),
            .I(N__28725));
    LocalMux I__5002 (
            .O(N__28783),
            .I(N__28725));
    LocalMux I__5001 (
            .O(N__28778),
            .I(N__28725));
    InMux I__5000 (
            .O(N__28777),
            .I(N__28722));
    InMux I__4999 (
            .O(N__28776),
            .I(N__28717));
    InMux I__4998 (
            .O(N__28775),
            .I(N__28717));
    InMux I__4997 (
            .O(N__28774),
            .I(N__28714));
    LocalMux I__4996 (
            .O(N__28769),
            .I(N__28709));
    LocalMux I__4995 (
            .O(N__28764),
            .I(N__28709));
    LocalMux I__4994 (
            .O(N__28757),
            .I(N__28704));
    Span4Mux_v I__4993 (
            .O(N__28750),
            .I(N__28704));
    Span4Mux_v I__4992 (
            .O(N__28745),
            .I(N__28701));
    Span4Mux_v I__4991 (
            .O(N__28742),
            .I(N__28692));
    Span4Mux_v I__4990 (
            .O(N__28735),
            .I(N__28692));
    Span4Mux_h I__4989 (
            .O(N__28732),
            .I(N__28692));
    Span4Mux_v I__4988 (
            .O(N__28725),
            .I(N__28692));
    LocalMux I__4987 (
            .O(N__28722),
            .I(n11683));
    LocalMux I__4986 (
            .O(N__28717),
            .I(n11683));
    LocalMux I__4985 (
            .O(N__28714),
            .I(n11683));
    Odrv4 I__4984 (
            .O(N__28709),
            .I(n11683));
    Odrv4 I__4983 (
            .O(N__28704),
            .I(n11683));
    Odrv4 I__4982 (
            .O(N__28701),
            .I(n11683));
    Odrv4 I__4981 (
            .O(N__28692),
            .I(n11683));
    CascadeMux I__4980 (
            .O(N__28677),
            .I(N__28674));
    InMux I__4979 (
            .O(N__28674),
            .I(N__28670));
    InMux I__4978 (
            .O(N__28673),
            .I(N__28667));
    LocalMux I__4977 (
            .O(N__28670),
            .I(N__28663));
    LocalMux I__4976 (
            .O(N__28667),
            .I(N__28660));
    InMux I__4975 (
            .O(N__28666),
            .I(N__28657));
    Span4Mux_v I__4974 (
            .O(N__28663),
            .I(N__28654));
    Odrv12 I__4973 (
            .O(N__28660),
            .I(timer_0));
    LocalMux I__4972 (
            .O(N__28657),
            .I(timer_0));
    Odrv4 I__4971 (
            .O(N__28654),
            .I(timer_0));
    InMux I__4970 (
            .O(N__28647),
            .I(N__28643));
    InMux I__4969 (
            .O(N__28646),
            .I(N__28640));
    LocalMux I__4968 (
            .O(N__28643),
            .I(neo_pixel_transmitter_t0_0));
    LocalMux I__4967 (
            .O(N__28640),
            .I(neo_pixel_transmitter_t0_0));
    InMux I__4966 (
            .O(N__28635),
            .I(N__28632));
    LocalMux I__4965 (
            .O(N__28632),
            .I(N__28629));
    Span12Mux_v I__4964 (
            .O(N__28629),
            .I(N__28626));
    Odrv12 I__4963 (
            .O(N__28626),
            .I(\nx.n33_adj_652 ));
    IoInMux I__4962 (
            .O(N__28623),
            .I(N__28620));
    LocalMux I__4961 (
            .O(N__28620),
            .I(N__28617));
    Span12Mux_s4_v I__4960 (
            .O(N__28617),
            .I(N__28614));
    Span12Mux_h I__4959 (
            .O(N__28614),
            .I(N__28609));
    CascadeMux I__4958 (
            .O(N__28613),
            .I(N__28606));
    InMux I__4957 (
            .O(N__28612),
            .I(N__28603));
    Span12Mux_v I__4956 (
            .O(N__28609),
            .I(N__28600));
    InMux I__4955 (
            .O(N__28606),
            .I(N__28597));
    LocalMux I__4954 (
            .O(N__28603),
            .I(N__28594));
    Odrv12 I__4953 (
            .O(N__28600),
            .I(pin_out_0));
    LocalMux I__4952 (
            .O(N__28597),
            .I(pin_out_0));
    Odrv4 I__4951 (
            .O(N__28594),
            .I(pin_out_0));
    IoInMux I__4950 (
            .O(N__28587),
            .I(N__28584));
    LocalMux I__4949 (
            .O(N__28584),
            .I(N__28581));
    IoSpan4Mux I__4948 (
            .O(N__28581),
            .I(N__28578));
    Span4Mux_s3_v I__4947 (
            .O(N__28578),
            .I(N__28575));
    Span4Mux_v I__4946 (
            .O(N__28575),
            .I(N__28572));
    Span4Mux_v I__4945 (
            .O(N__28572),
            .I(N__28568));
    CascadeMux I__4944 (
            .O(N__28571),
            .I(N__28565));
    Span4Mux_v I__4943 (
            .O(N__28568),
            .I(N__28561));
    InMux I__4942 (
            .O(N__28565),
            .I(N__28558));
    InMux I__4941 (
            .O(N__28564),
            .I(N__28555));
    Odrv4 I__4940 (
            .O(N__28561),
            .I(pin_out_1));
    LocalMux I__4939 (
            .O(N__28558),
            .I(pin_out_1));
    LocalMux I__4938 (
            .O(N__28555),
            .I(pin_out_1));
    InMux I__4937 (
            .O(N__28548),
            .I(N__28545));
    LocalMux I__4936 (
            .O(N__28545),
            .I(N__28540));
    InMux I__4935 (
            .O(N__28544),
            .I(N__28537));
    InMux I__4934 (
            .O(N__28543),
            .I(N__28534));
    Span4Mux_v I__4933 (
            .O(N__28540),
            .I(N__28530));
    LocalMux I__4932 (
            .O(N__28537),
            .I(N__28527));
    LocalMux I__4931 (
            .O(N__28534),
            .I(N__28524));
    InMux I__4930 (
            .O(N__28533),
            .I(N__28520));
    Span4Mux_v I__4929 (
            .O(N__28530),
            .I(N__28517));
    Span4Mux_v I__4928 (
            .O(N__28527),
            .I(N__28512));
    Span4Mux_v I__4927 (
            .O(N__28524),
            .I(N__28512));
    InMux I__4926 (
            .O(N__28523),
            .I(N__28509));
    LocalMux I__4925 (
            .O(N__28520),
            .I(N__28506));
    Span4Mux_h I__4924 (
            .O(N__28517),
            .I(N__28503));
    Span4Mux_v I__4923 (
            .O(N__28512),
            .I(N__28500));
    LocalMux I__4922 (
            .O(N__28509),
            .I(\nx.bit_ctr_8 ));
    Odrv4 I__4921 (
            .O(N__28506),
            .I(\nx.bit_ctr_8 ));
    Odrv4 I__4920 (
            .O(N__28503),
            .I(\nx.bit_ctr_8 ));
    Odrv4 I__4919 (
            .O(N__28500),
            .I(\nx.bit_ctr_8 ));
    InMux I__4918 (
            .O(N__28491),
            .I(N__28488));
    LocalMux I__4917 (
            .O(N__28488),
            .I(N__28485));
    Span4Mux_h I__4916 (
            .O(N__28485),
            .I(N__28482));
    Odrv4 I__4915 (
            .O(N__28482),
            .I(\nx.n2777 ));
    InMux I__4914 (
            .O(N__28479),
            .I(bfn_7_19_0_));
    InMux I__4913 (
            .O(N__28476),
            .I(N__28469));
    InMux I__4912 (
            .O(N__28475),
            .I(N__28469));
    CascadeMux I__4911 (
            .O(N__28474),
            .I(N__28466));
    LocalMux I__4910 (
            .O(N__28469),
            .I(N__28463));
    InMux I__4909 (
            .O(N__28466),
            .I(N__28460));
    Odrv4 I__4908 (
            .O(N__28463),
            .I(\nx.n1507 ));
    LocalMux I__4907 (
            .O(N__28460),
            .I(\nx.n1507 ));
    CascadeMux I__4906 (
            .O(N__28455),
            .I(N__28452));
    InMux I__4905 (
            .O(N__28452),
            .I(N__28449));
    LocalMux I__4904 (
            .O(N__28449),
            .I(N__28446));
    Odrv4 I__4903 (
            .O(N__28446),
            .I(\nx.n1574 ));
    InMux I__4902 (
            .O(N__28443),
            .I(\nx.n10594 ));
    InMux I__4901 (
            .O(N__28440),
            .I(\nx.n10595 ));
    InMux I__4900 (
            .O(N__28437),
            .I(N__28434));
    LocalMux I__4899 (
            .O(N__28434),
            .I(N__28429));
    InMux I__4898 (
            .O(N__28433),
            .I(N__28426));
    CascadeMux I__4897 (
            .O(N__28432),
            .I(N__28423));
    Span4Mux_h I__4896 (
            .O(N__28429),
            .I(N__28418));
    LocalMux I__4895 (
            .O(N__28426),
            .I(N__28418));
    InMux I__4894 (
            .O(N__28423),
            .I(N__28415));
    Odrv4 I__4893 (
            .O(N__28418),
            .I(\nx.n1505 ));
    LocalMux I__4892 (
            .O(N__28415),
            .I(\nx.n1505 ));
    InMux I__4891 (
            .O(N__28410),
            .I(N__28407));
    LocalMux I__4890 (
            .O(N__28407),
            .I(N__28404));
    Odrv4 I__4889 (
            .O(N__28404),
            .I(\nx.n1572 ));
    InMux I__4888 (
            .O(N__28401),
            .I(\nx.n10596 ));
    CascadeMux I__4887 (
            .O(N__28398),
            .I(N__28394));
    InMux I__4886 (
            .O(N__28397),
            .I(N__28388));
    InMux I__4885 (
            .O(N__28394),
            .I(N__28388));
    CascadeMux I__4884 (
            .O(N__28393),
            .I(N__28385));
    LocalMux I__4883 (
            .O(N__28388),
            .I(N__28382));
    InMux I__4882 (
            .O(N__28385),
            .I(N__28379));
    Span4Mux_h I__4881 (
            .O(N__28382),
            .I(N__28376));
    LocalMux I__4880 (
            .O(N__28379),
            .I(\nx.n1504 ));
    Odrv4 I__4879 (
            .O(N__28376),
            .I(\nx.n1504 ));
    InMux I__4878 (
            .O(N__28371),
            .I(N__28368));
    LocalMux I__4877 (
            .O(N__28368),
            .I(N__28365));
    Odrv4 I__4876 (
            .O(N__28365),
            .I(\nx.n1571 ));
    InMux I__4875 (
            .O(N__28362),
            .I(\nx.n10597 ));
    InMux I__4874 (
            .O(N__28359),
            .I(\nx.n10598 ));
    CascadeMux I__4873 (
            .O(N__28356),
            .I(N__28352));
    InMux I__4872 (
            .O(N__28355),
            .I(N__28348));
    InMux I__4871 (
            .O(N__28352),
            .I(N__28345));
    InMux I__4870 (
            .O(N__28351),
            .I(N__28342));
    LocalMux I__4869 (
            .O(N__28348),
            .I(\nx.n1502 ));
    LocalMux I__4868 (
            .O(N__28345),
            .I(\nx.n1502 ));
    LocalMux I__4867 (
            .O(N__28342),
            .I(\nx.n1502 ));
    InMux I__4866 (
            .O(N__28335),
            .I(N__28332));
    LocalMux I__4865 (
            .O(N__28332),
            .I(N__28329));
    Odrv4 I__4864 (
            .O(N__28329),
            .I(\nx.n1569 ));
    InMux I__4863 (
            .O(N__28326),
            .I(bfn_6_32_0_));
    InMux I__4862 (
            .O(N__28323),
            .I(N__28319));
    CascadeMux I__4861 (
            .O(N__28322),
            .I(N__28316));
    LocalMux I__4860 (
            .O(N__28319),
            .I(N__28313));
    InMux I__4859 (
            .O(N__28316),
            .I(N__28310));
    Span4Mux_v I__4858 (
            .O(N__28313),
            .I(N__28305));
    LocalMux I__4857 (
            .O(N__28310),
            .I(N__28305));
    Odrv4 I__4856 (
            .O(N__28305),
            .I(\nx.n1501 ));
    CascadeMux I__4855 (
            .O(N__28302),
            .I(N__28299));
    InMux I__4854 (
            .O(N__28299),
            .I(N__28296));
    LocalMux I__4853 (
            .O(N__28296),
            .I(N__28293));
    Odrv4 I__4852 (
            .O(N__28293),
            .I(\nx.n1568 ));
    InMux I__4851 (
            .O(N__28290),
            .I(\nx.n10600 ));
    InMux I__4850 (
            .O(N__28287),
            .I(N__28283));
    CascadeMux I__4849 (
            .O(N__28286),
            .I(N__28280));
    LocalMux I__4848 (
            .O(N__28283),
            .I(N__28276));
    InMux I__4847 (
            .O(N__28280),
            .I(N__28273));
    InMux I__4846 (
            .O(N__28279),
            .I(N__28270));
    Odrv4 I__4845 (
            .O(N__28276),
            .I(\nx.n1500 ));
    LocalMux I__4844 (
            .O(N__28273),
            .I(\nx.n1500 ));
    LocalMux I__4843 (
            .O(N__28270),
            .I(\nx.n1500 ));
    CascadeMux I__4842 (
            .O(N__28263),
            .I(N__28260));
    InMux I__4841 (
            .O(N__28260),
            .I(N__28257));
    LocalMux I__4840 (
            .O(N__28257),
            .I(N__28254));
    Odrv4 I__4839 (
            .O(N__28254),
            .I(\nx.n1567 ));
    InMux I__4838 (
            .O(N__28251),
            .I(\nx.n10601 ));
    InMux I__4837 (
            .O(N__28248),
            .I(N__28244));
    CascadeMux I__4836 (
            .O(N__28247),
            .I(N__28240));
    LocalMux I__4835 (
            .O(N__28244),
            .I(N__28237));
    InMux I__4834 (
            .O(N__28243),
            .I(N__28234));
    InMux I__4833 (
            .O(N__28240),
            .I(N__28231));
    Odrv12 I__4832 (
            .O(N__28237),
            .I(\nx.n1409 ));
    LocalMux I__4831 (
            .O(N__28234),
            .I(\nx.n1409 ));
    LocalMux I__4830 (
            .O(N__28231),
            .I(\nx.n1409 ));
    CascadeMux I__4829 (
            .O(N__28224),
            .I(N__28221));
    InMux I__4828 (
            .O(N__28221),
            .I(N__28218));
    LocalMux I__4827 (
            .O(N__28218),
            .I(N__28215));
    Span4Mux_v I__4826 (
            .O(N__28215),
            .I(N__28212));
    Odrv4 I__4825 (
            .O(N__28212),
            .I(\nx.n1476 ));
    InMux I__4824 (
            .O(N__28209),
            .I(N__28204));
    CascadeMux I__4823 (
            .O(N__28208),
            .I(N__28199));
    CascadeMux I__4822 (
            .O(N__28207),
            .I(N__28196));
    LocalMux I__4821 (
            .O(N__28204),
            .I(N__28192));
    CascadeMux I__4820 (
            .O(N__28203),
            .I(N__28189));
    CascadeMux I__4819 (
            .O(N__28202),
            .I(N__28183));
    InMux I__4818 (
            .O(N__28199),
            .I(N__28175));
    InMux I__4817 (
            .O(N__28196),
            .I(N__28175));
    InMux I__4816 (
            .O(N__28195),
            .I(N__28175));
    Span4Mux_h I__4815 (
            .O(N__28192),
            .I(N__28172));
    InMux I__4814 (
            .O(N__28189),
            .I(N__28169));
    InMux I__4813 (
            .O(N__28188),
            .I(N__28162));
    InMux I__4812 (
            .O(N__28187),
            .I(N__28162));
    InMux I__4811 (
            .O(N__28186),
            .I(N__28162));
    InMux I__4810 (
            .O(N__28183),
            .I(N__28157));
    InMux I__4809 (
            .O(N__28182),
            .I(N__28157));
    LocalMux I__4808 (
            .O(N__28175),
            .I(\nx.n1433 ));
    Odrv4 I__4807 (
            .O(N__28172),
            .I(\nx.n1433 ));
    LocalMux I__4806 (
            .O(N__28169),
            .I(\nx.n1433 ));
    LocalMux I__4805 (
            .O(N__28162),
            .I(\nx.n1433 ));
    LocalMux I__4804 (
            .O(N__28157),
            .I(\nx.n1433 ));
    CascadeMux I__4803 (
            .O(N__28146),
            .I(\nx.n1508_cascade_ ));
    InMux I__4802 (
            .O(N__28143),
            .I(N__28140));
    LocalMux I__4801 (
            .O(N__28140),
            .I(\nx.n16_adj_633 ));
    CascadeMux I__4800 (
            .O(N__28137),
            .I(\nx.n1599_cascade_ ));
    InMux I__4799 (
            .O(N__28134),
            .I(bfn_6_31_0_));
    InMux I__4798 (
            .O(N__28131),
            .I(\nx.n10592 ));
    CascadeMux I__4797 (
            .O(N__28128),
            .I(N__28124));
    CascadeMux I__4796 (
            .O(N__28127),
            .I(N__28121));
    InMux I__4795 (
            .O(N__28124),
            .I(N__28118));
    InMux I__4794 (
            .O(N__28121),
            .I(N__28115));
    LocalMux I__4793 (
            .O(N__28118),
            .I(\nx.n1508 ));
    LocalMux I__4792 (
            .O(N__28115),
            .I(\nx.n1508 ));
    InMux I__4791 (
            .O(N__28110),
            .I(N__28107));
    LocalMux I__4790 (
            .O(N__28107),
            .I(N__28104));
    Odrv4 I__4789 (
            .O(N__28104),
            .I(\nx.n1575 ));
    InMux I__4788 (
            .O(N__28101),
            .I(\nx.n10593 ));
    InMux I__4787 (
            .O(N__28098),
            .I(N__28095));
    LocalMux I__4786 (
            .O(N__28095),
            .I(N__28092));
    Odrv4 I__4785 (
            .O(N__28092),
            .I(\nx.n20_adj_634 ));
    CascadeMux I__4784 (
            .O(N__28089),
            .I(\nx.n1532_cascade_ ));
    CascadeMux I__4783 (
            .O(N__28086),
            .I(\nx.n1606_cascade_ ));
    CascadeMux I__4782 (
            .O(N__28083),
            .I(\nx.n22_adj_647_cascade_ ));
    CascadeMux I__4781 (
            .O(N__28080),
            .I(\nx.n1631_cascade_ ));
    InMux I__4780 (
            .O(N__28077),
            .I(N__28074));
    LocalMux I__4779 (
            .O(N__28074),
            .I(\nx.n19_adj_602 ));
    CascadeMux I__4778 (
            .O(N__28071),
            .I(N__28066));
    CascadeMux I__4777 (
            .O(N__28070),
            .I(N__28063));
    InMux I__4776 (
            .O(N__28069),
            .I(N__28060));
    InMux I__4775 (
            .O(N__28066),
            .I(N__28057));
    InMux I__4774 (
            .O(N__28063),
            .I(N__28053));
    LocalMux I__4773 (
            .O(N__28060),
            .I(N__28049));
    LocalMux I__4772 (
            .O(N__28057),
            .I(N__28046));
    InMux I__4771 (
            .O(N__28056),
            .I(N__28043));
    LocalMux I__4770 (
            .O(N__28053),
            .I(N__28040));
    InMux I__4769 (
            .O(N__28052),
            .I(N__28037));
    Span4Mux_v I__4768 (
            .O(N__28049),
            .I(N__28032));
    Span4Mux_v I__4767 (
            .O(N__28046),
            .I(N__28032));
    LocalMux I__4766 (
            .O(N__28043),
            .I(\nx.bit_ctr_26 ));
    Odrv4 I__4765 (
            .O(N__28040),
            .I(\nx.bit_ctr_26 ));
    LocalMux I__4764 (
            .O(N__28037),
            .I(\nx.bit_ctr_26 ));
    Odrv4 I__4763 (
            .O(N__28032),
            .I(\nx.bit_ctr_26 ));
    InMux I__4762 (
            .O(N__28023),
            .I(N__28020));
    LocalMux I__4761 (
            .O(N__28020),
            .I(\nx.n977 ));
    InMux I__4760 (
            .O(N__28017),
            .I(bfn_6_28_0_));
    CascadeMux I__4759 (
            .O(N__28014),
            .I(N__28010));
    InMux I__4758 (
            .O(N__28013),
            .I(N__28007));
    InMux I__4757 (
            .O(N__28010),
            .I(N__28004));
    LocalMux I__4756 (
            .O(N__28007),
            .I(\nx.n7082 ));
    LocalMux I__4755 (
            .O(N__28004),
            .I(\nx.n7082 ));
    CascadeMux I__4754 (
            .O(N__27999),
            .I(N__27996));
    InMux I__4753 (
            .O(N__27996),
            .I(N__27993));
    LocalMux I__4752 (
            .O(N__27993),
            .I(\nx.n976 ));
    InMux I__4751 (
            .O(N__27990),
            .I(\nx.n10474 ));
    CascadeMux I__4750 (
            .O(N__27987),
            .I(N__27984));
    InMux I__4749 (
            .O(N__27984),
            .I(N__27980));
    InMux I__4748 (
            .O(N__27983),
            .I(N__27977));
    LocalMux I__4747 (
            .O(N__27980),
            .I(\nx.n7342 ));
    LocalMux I__4746 (
            .O(N__27977),
            .I(\nx.n7342 ));
    CascadeMux I__4745 (
            .O(N__27972),
            .I(N__27968));
    InMux I__4744 (
            .O(N__27971),
            .I(N__27963));
    InMux I__4743 (
            .O(N__27968),
            .I(N__27963));
    LocalMux I__4742 (
            .O(N__27963),
            .I(\nx.n975 ));
    InMux I__4741 (
            .O(N__27960),
            .I(\nx.n10475 ));
    CascadeMux I__4740 (
            .O(N__27957),
            .I(N__27953));
    InMux I__4739 (
            .O(N__27956),
            .I(N__27950));
    InMux I__4738 (
            .O(N__27953),
            .I(N__27947));
    LocalMux I__4737 (
            .O(N__27950),
            .I(\nx.n974 ));
    LocalMux I__4736 (
            .O(N__27947),
            .I(\nx.n974 ));
    InMux I__4735 (
            .O(N__27942),
            .I(\nx.n10476 ));
    CascadeMux I__4734 (
            .O(N__27939),
            .I(N__27935));
    CascadeMux I__4733 (
            .O(N__27938),
            .I(N__27932));
    InMux I__4732 (
            .O(N__27935),
            .I(N__27928));
    InMux I__4731 (
            .O(N__27932),
            .I(N__27925));
    InMux I__4730 (
            .O(N__27931),
            .I(N__27922));
    LocalMux I__4729 (
            .O(N__27928),
            .I(\nx.n906 ));
    LocalMux I__4728 (
            .O(N__27925),
            .I(\nx.n906 ));
    LocalMux I__4727 (
            .O(N__27922),
            .I(\nx.n906 ));
    InMux I__4726 (
            .O(N__27915),
            .I(N__27912));
    LocalMux I__4725 (
            .O(N__27912),
            .I(\nx.n973 ));
    InMux I__4724 (
            .O(N__27909),
            .I(\nx.n10477 ));
    InMux I__4723 (
            .O(N__27906),
            .I(N__27902));
    InMux I__4722 (
            .O(N__27905),
            .I(N__27899));
    LocalMux I__4721 (
            .O(N__27902),
            .I(\nx.n13064 ));
    LocalMux I__4720 (
            .O(N__27899),
            .I(\nx.n13064 ));
    InMux I__4719 (
            .O(N__27894),
            .I(\nx.n10478 ));
    CascadeMux I__4718 (
            .O(N__27891),
            .I(N__27888));
    InMux I__4717 (
            .O(N__27888),
            .I(N__27885));
    LocalMux I__4716 (
            .O(N__27885),
            .I(N__27881));
    InMux I__4715 (
            .O(N__27884),
            .I(N__27878));
    Odrv4 I__4714 (
            .O(N__27881),
            .I(\nx.n4_adj_596 ));
    LocalMux I__4713 (
            .O(N__27878),
            .I(\nx.n4_adj_596 ));
    InMux I__4712 (
            .O(N__27873),
            .I(N__27866));
    InMux I__4711 (
            .O(N__27872),
            .I(N__27866));
    InMux I__4710 (
            .O(N__27871),
            .I(N__27863));
    LocalMux I__4709 (
            .O(N__27866),
            .I(N__27860));
    LocalMux I__4708 (
            .O(N__27863),
            .I(\nx.n5260 ));
    Odrv4 I__4707 (
            .O(N__27860),
            .I(\nx.n5260 ));
    CascadeMux I__4706 (
            .O(N__27855),
            .I(N__27850));
    InMux I__4705 (
            .O(N__27854),
            .I(N__27845));
    InMux I__4704 (
            .O(N__27853),
            .I(N__27845));
    InMux I__4703 (
            .O(N__27850),
            .I(N__27842));
    LocalMux I__4702 (
            .O(N__27845),
            .I(N__27838));
    LocalMux I__4701 (
            .O(N__27842),
            .I(N__27835));
    InMux I__4700 (
            .O(N__27841),
            .I(N__27832));
    Odrv12 I__4699 (
            .O(N__27838),
            .I(\nx.n11559 ));
    Odrv4 I__4698 (
            .O(N__27835),
            .I(\nx.n11559 ));
    LocalMux I__4697 (
            .O(N__27832),
            .I(\nx.n11559 ));
    CascadeMux I__4696 (
            .O(N__27825),
            .I(N__27820));
    CascadeMux I__4695 (
            .O(N__27824),
            .I(N__27817));
    InMux I__4694 (
            .O(N__27823),
            .I(N__27812));
    InMux I__4693 (
            .O(N__27820),
            .I(N__27803));
    InMux I__4692 (
            .O(N__27817),
            .I(N__27803));
    InMux I__4691 (
            .O(N__27816),
            .I(N__27803));
    InMux I__4690 (
            .O(N__27815),
            .I(N__27803));
    LocalMux I__4689 (
            .O(N__27812),
            .I(\nx.n838 ));
    LocalMux I__4688 (
            .O(N__27803),
            .I(\nx.n838 ));
    CascadeMux I__4687 (
            .O(N__27798),
            .I(N__27795));
    InMux I__4686 (
            .O(N__27795),
            .I(N__27791));
    InMux I__4685 (
            .O(N__27794),
            .I(N__27788));
    LocalMux I__4684 (
            .O(N__27791),
            .I(\nx.n11674 ));
    LocalMux I__4683 (
            .O(N__27788),
            .I(\nx.n11674 ));
    CascadeMux I__4682 (
            .O(N__27783),
            .I(\nx.n1829_cascade_ ));
    CascadeMux I__4681 (
            .O(N__27780),
            .I(\nx.n1906_cascade_ ));
    CascadeMux I__4680 (
            .O(N__27777),
            .I(N__27774));
    InMux I__4679 (
            .O(N__27774),
            .I(N__27771));
    LocalMux I__4678 (
            .O(N__27771),
            .I(\nx.n22_adj_605 ));
    CascadeMux I__4677 (
            .O(N__27768),
            .I(N__27764));
    CascadeMux I__4676 (
            .O(N__27767),
            .I(N__27761));
    InMux I__4675 (
            .O(N__27764),
            .I(N__27758));
    InMux I__4674 (
            .O(N__27761),
            .I(N__27755));
    LocalMux I__4673 (
            .O(N__27758),
            .I(\nx.n1006 ));
    LocalMux I__4672 (
            .O(N__27755),
            .I(\nx.n1006 ));
    CascadeMux I__4671 (
            .O(N__27750),
            .I(\nx.n1804_cascade_ ));
    CascadeMux I__4670 (
            .O(N__27747),
            .I(\nx.n19_cascade_ ));
    InMux I__4669 (
            .O(N__27744),
            .I(N__27741));
    LocalMux I__4668 (
            .O(N__27741),
            .I(\nx.n26_adj_600 ));
    InMux I__4667 (
            .O(N__27738),
            .I(N__27733));
    InMux I__4666 (
            .O(N__27737),
            .I(N__27729));
    CascadeMux I__4665 (
            .O(N__27736),
            .I(N__27725));
    LocalMux I__4664 (
            .O(N__27733),
            .I(N__27720));
    InMux I__4663 (
            .O(N__27732),
            .I(N__27717));
    LocalMux I__4662 (
            .O(N__27729),
            .I(N__27714));
    InMux I__4661 (
            .O(N__27728),
            .I(N__27711));
    InMux I__4660 (
            .O(N__27725),
            .I(N__27704));
    InMux I__4659 (
            .O(N__27724),
            .I(N__27704));
    InMux I__4658 (
            .O(N__27723),
            .I(N__27704));
    Span4Mux_h I__4657 (
            .O(N__27720),
            .I(N__27701));
    LocalMux I__4656 (
            .O(N__27717),
            .I(\nx.bit_ctr_27 ));
    Odrv4 I__4655 (
            .O(N__27714),
            .I(\nx.bit_ctr_27 ));
    LocalMux I__4654 (
            .O(N__27711),
            .I(\nx.bit_ctr_27 ));
    LocalMux I__4653 (
            .O(N__27704),
            .I(\nx.bit_ctr_27 ));
    Odrv4 I__4652 (
            .O(N__27701),
            .I(\nx.bit_ctr_27 ));
    CascadeMux I__4651 (
            .O(N__27690),
            .I(N__27686));
    InMux I__4650 (
            .O(N__27689),
            .I(N__27683));
    InMux I__4649 (
            .O(N__27686),
            .I(N__27679));
    LocalMux I__4648 (
            .O(N__27683),
            .I(N__27675));
    CascadeMux I__4647 (
            .O(N__27682),
            .I(N__27671));
    LocalMux I__4646 (
            .O(N__27679),
            .I(N__27668));
    InMux I__4645 (
            .O(N__27678),
            .I(N__27663));
    Span4Mux_h I__4644 (
            .O(N__27675),
            .I(N__27660));
    InMux I__4643 (
            .O(N__27674),
            .I(N__27655));
    InMux I__4642 (
            .O(N__27671),
            .I(N__27655));
    Span4Mux_v I__4641 (
            .O(N__27668),
            .I(N__27652));
    InMux I__4640 (
            .O(N__27667),
            .I(N__27647));
    InMux I__4639 (
            .O(N__27666),
            .I(N__27647));
    LocalMux I__4638 (
            .O(N__27663),
            .I(\nx.bit_ctr_28 ));
    Odrv4 I__4637 (
            .O(N__27660),
            .I(\nx.bit_ctr_28 ));
    LocalMux I__4636 (
            .O(N__27655),
            .I(\nx.bit_ctr_28 ));
    Odrv4 I__4635 (
            .O(N__27652),
            .I(\nx.bit_ctr_28 ));
    LocalMux I__4634 (
            .O(N__27647),
            .I(\nx.bit_ctr_28 ));
    CascadeMux I__4633 (
            .O(N__27636),
            .I(N__27632));
    InMux I__4632 (
            .O(N__27635),
            .I(N__27628));
    InMux I__4631 (
            .O(N__27632),
            .I(N__27622));
    InMux I__4630 (
            .O(N__27631),
            .I(N__27622));
    LocalMux I__4629 (
            .O(N__27628),
            .I(N__27619));
    InMux I__4628 (
            .O(N__27627),
            .I(N__27616));
    LocalMux I__4627 (
            .O(N__27622),
            .I(\nx.n739 ));
    Odrv4 I__4626 (
            .O(N__27619),
            .I(\nx.n739 ));
    LocalMux I__4625 (
            .O(N__27616),
            .I(\nx.n739 ));
    CascadeMux I__4624 (
            .O(N__27609),
            .I(\nx.n28_adj_660_cascade_ ));
    InMux I__4623 (
            .O(N__27606),
            .I(N__27603));
    LocalMux I__4622 (
            .O(N__27603),
            .I(\nx.n16 ));
    CascadeMux I__4621 (
            .O(N__27600),
            .I(\nx.n1928_cascade_ ));
    CascadeMux I__4620 (
            .O(N__27597),
            .I(\nx.n1908_cascade_ ));
    InMux I__4619 (
            .O(N__27594),
            .I(N__27591));
    LocalMux I__4618 (
            .O(N__27591),
            .I(\nx.n24_adj_648 ));
    InMux I__4617 (
            .O(N__27588),
            .I(N__27585));
    LocalMux I__4616 (
            .O(N__27585),
            .I(\nx.n1877 ));
    InMux I__4615 (
            .O(N__27582),
            .I(bfn_6_24_0_));
    InMux I__4614 (
            .O(N__27579),
            .I(N__27575));
    CascadeMux I__4613 (
            .O(N__27578),
            .I(N__27572));
    LocalMux I__4612 (
            .O(N__27575),
            .I(N__27569));
    InMux I__4611 (
            .O(N__27572),
            .I(N__27566));
    Span4Mux_v I__4610 (
            .O(N__27569),
            .I(N__27563));
    LocalMux I__4609 (
            .O(N__27566),
            .I(\nx.n2885 ));
    Odrv4 I__4608 (
            .O(N__27563),
            .I(\nx.n2885 ));
    InMux I__4607 (
            .O(N__27558),
            .I(N__27555));
    LocalMux I__4606 (
            .O(N__27555),
            .I(\nx.n2858 ));
    CascadeMux I__4605 (
            .O(N__27552),
            .I(\nx.n2791_cascade_ ));
    InMux I__4604 (
            .O(N__27549),
            .I(N__27546));
    LocalMux I__4603 (
            .O(N__27546),
            .I(\nx.n2859 ));
    InMux I__4602 (
            .O(N__27543),
            .I(N__27538));
    InMux I__4601 (
            .O(N__27542),
            .I(N__27535));
    CascadeMux I__4600 (
            .O(N__27541),
            .I(N__27532));
    LocalMux I__4599 (
            .O(N__27538),
            .I(N__27529));
    LocalMux I__4598 (
            .O(N__27535),
            .I(N__27526));
    InMux I__4597 (
            .O(N__27532),
            .I(N__27523));
    Span4Mux_h I__4596 (
            .O(N__27529),
            .I(N__27520));
    Odrv4 I__4595 (
            .O(N__27526),
            .I(\nx.n2891 ));
    LocalMux I__4594 (
            .O(N__27523),
            .I(\nx.n2891 ));
    Odrv4 I__4593 (
            .O(N__27520),
            .I(\nx.n2891 ));
    InMux I__4592 (
            .O(N__27513),
            .I(N__27510));
    LocalMux I__4591 (
            .O(N__27510),
            .I(\nx.n2856 ));
    CascadeMux I__4590 (
            .O(N__27507),
            .I(\nx.n2789_cascade_ ));
    InMux I__4589 (
            .O(N__27504),
            .I(N__27500));
    InMux I__4588 (
            .O(N__27503),
            .I(N__27497));
    LocalMux I__4587 (
            .O(N__27500),
            .I(N__27494));
    LocalMux I__4586 (
            .O(N__27497),
            .I(N__27491));
    Span4Mux_v I__4585 (
            .O(N__27494),
            .I(N__27488));
    Span4Mux_v I__4584 (
            .O(N__27491),
            .I(N__27485));
    Odrv4 I__4583 (
            .O(N__27488),
            .I(\nx.n2995 ));
    Odrv4 I__4582 (
            .O(N__27485),
            .I(\nx.n2995 ));
    CascadeMux I__4581 (
            .O(N__27480),
            .I(N__27477));
    InMux I__4580 (
            .O(N__27477),
            .I(N__27474));
    LocalMux I__4579 (
            .O(N__27474),
            .I(N__27471));
    Span4Mux_h I__4578 (
            .O(N__27471),
            .I(N__27468));
    Odrv4 I__4577 (
            .O(N__27468),
            .I(\nx.n3062 ));
    CascadeMux I__4576 (
            .O(N__27465),
            .I(N__27460));
    CascadeMux I__4575 (
            .O(N__27464),
            .I(N__27453));
    InMux I__4574 (
            .O(N__27463),
            .I(N__27448));
    InMux I__4573 (
            .O(N__27460),
            .I(N__27445));
    InMux I__4572 (
            .O(N__27459),
            .I(N__27442));
    InMux I__4571 (
            .O(N__27458),
            .I(N__27433));
    InMux I__4570 (
            .O(N__27457),
            .I(N__27430));
    InMux I__4569 (
            .O(N__27456),
            .I(N__27423));
    InMux I__4568 (
            .O(N__27453),
            .I(N__27423));
    InMux I__4567 (
            .O(N__27452),
            .I(N__27423));
    CascadeMux I__4566 (
            .O(N__27451),
            .I(N__27416));
    LocalMux I__4565 (
            .O(N__27448),
            .I(N__27412));
    LocalMux I__4564 (
            .O(N__27445),
            .I(N__27407));
    LocalMux I__4563 (
            .O(N__27442),
            .I(N__27407));
    InMux I__4562 (
            .O(N__27441),
            .I(N__27402));
    InMux I__4561 (
            .O(N__27440),
            .I(N__27402));
    CascadeMux I__4560 (
            .O(N__27439),
            .I(N__27396));
    CascadeMux I__4559 (
            .O(N__27438),
            .I(N__27393));
    CascadeMux I__4558 (
            .O(N__27437),
            .I(N__27390));
    CascadeMux I__4557 (
            .O(N__27436),
            .I(N__27384));
    LocalMux I__4556 (
            .O(N__27433),
            .I(N__27377));
    LocalMux I__4555 (
            .O(N__27430),
            .I(N__27377));
    LocalMux I__4554 (
            .O(N__27423),
            .I(N__27377));
    InMux I__4553 (
            .O(N__27422),
            .I(N__27372));
    InMux I__4552 (
            .O(N__27421),
            .I(N__27372));
    InMux I__4551 (
            .O(N__27420),
            .I(N__27363));
    InMux I__4550 (
            .O(N__27419),
            .I(N__27363));
    InMux I__4549 (
            .O(N__27416),
            .I(N__27363));
    InMux I__4548 (
            .O(N__27415),
            .I(N__27363));
    Span4Mux_v I__4547 (
            .O(N__27412),
            .I(N__27360));
    Span4Mux_v I__4546 (
            .O(N__27407),
            .I(N__27355));
    LocalMux I__4545 (
            .O(N__27402),
            .I(N__27355));
    InMux I__4544 (
            .O(N__27401),
            .I(N__27350));
    InMux I__4543 (
            .O(N__27400),
            .I(N__27350));
    InMux I__4542 (
            .O(N__27399),
            .I(N__27339));
    InMux I__4541 (
            .O(N__27396),
            .I(N__27339));
    InMux I__4540 (
            .O(N__27393),
            .I(N__27339));
    InMux I__4539 (
            .O(N__27390),
            .I(N__27339));
    InMux I__4538 (
            .O(N__27389),
            .I(N__27339));
    InMux I__4537 (
            .O(N__27388),
            .I(N__27332));
    InMux I__4536 (
            .O(N__27387),
            .I(N__27332));
    InMux I__4535 (
            .O(N__27384),
            .I(N__27332));
    Span4Mux_h I__4534 (
            .O(N__27377),
            .I(N__27329));
    LocalMux I__4533 (
            .O(N__27372),
            .I(\nx.n3017 ));
    LocalMux I__4532 (
            .O(N__27363),
            .I(\nx.n3017 ));
    Odrv4 I__4531 (
            .O(N__27360),
            .I(\nx.n3017 ));
    Odrv4 I__4530 (
            .O(N__27355),
            .I(\nx.n3017 ));
    LocalMux I__4529 (
            .O(N__27350),
            .I(\nx.n3017 ));
    LocalMux I__4528 (
            .O(N__27339),
            .I(\nx.n3017 ));
    LocalMux I__4527 (
            .O(N__27332),
            .I(\nx.n3017 ));
    Odrv4 I__4526 (
            .O(N__27329),
            .I(\nx.n3017 ));
    InMux I__4525 (
            .O(N__27312),
            .I(N__27308));
    InMux I__4524 (
            .O(N__27311),
            .I(N__27304));
    LocalMux I__4523 (
            .O(N__27308),
            .I(N__27301));
    CascadeMux I__4522 (
            .O(N__27307),
            .I(N__27298));
    LocalMux I__4521 (
            .O(N__27304),
            .I(N__27293));
    Span12Mux_s7_v I__4520 (
            .O(N__27301),
            .I(N__27293));
    InMux I__4519 (
            .O(N__27298),
            .I(N__27290));
    Odrv12 I__4518 (
            .O(N__27293),
            .I(\nx.n3094 ));
    LocalMux I__4517 (
            .O(N__27290),
            .I(\nx.n3094 ));
    InMux I__4516 (
            .O(N__27285),
            .I(N__27281));
    CascadeMux I__4515 (
            .O(N__27284),
            .I(N__27278));
    LocalMux I__4514 (
            .O(N__27281),
            .I(N__27275));
    InMux I__4513 (
            .O(N__27278),
            .I(N__27272));
    Span4Mux_h I__4512 (
            .O(N__27275),
            .I(N__27266));
    LocalMux I__4511 (
            .O(N__27272),
            .I(N__27266));
    InMux I__4510 (
            .O(N__27271),
            .I(N__27263));
    Odrv4 I__4509 (
            .O(N__27266),
            .I(\nx.n2795 ));
    LocalMux I__4508 (
            .O(N__27263),
            .I(\nx.n2795 ));
    CascadeMux I__4507 (
            .O(N__27258),
            .I(N__27255));
    InMux I__4506 (
            .O(N__27255),
            .I(N__27252));
    LocalMux I__4505 (
            .O(N__27252),
            .I(N__27249));
    Odrv4 I__4504 (
            .O(N__27249),
            .I(\nx.n2862 ));
    InMux I__4503 (
            .O(N__27246),
            .I(\nx.n10827 ));
    InMux I__4502 (
            .O(N__27243),
            .I(bfn_6_23_0_));
    InMux I__4501 (
            .O(N__27240),
            .I(\nx.n10829 ));
    InMux I__4500 (
            .O(N__27237),
            .I(\nx.n10830 ));
    InMux I__4499 (
            .O(N__27234),
            .I(\nx.n10831 ));
    InMux I__4498 (
            .O(N__27231),
            .I(\nx.n10832 ));
    InMux I__4497 (
            .O(N__27228),
            .I(\nx.n10833 ));
    InMux I__4496 (
            .O(N__27225),
            .I(\nx.n10834 ));
    InMux I__4495 (
            .O(N__27222),
            .I(\nx.n10835 ));
    InMux I__4494 (
            .O(N__27219),
            .I(\nx.n10819 ));
    CascadeMux I__4493 (
            .O(N__27216),
            .I(N__27212));
    CascadeMux I__4492 (
            .O(N__27215),
            .I(N__27209));
    InMux I__4491 (
            .O(N__27212),
            .I(N__27206));
    InMux I__4490 (
            .O(N__27209),
            .I(N__27203));
    LocalMux I__4489 (
            .O(N__27206),
            .I(N__27199));
    LocalMux I__4488 (
            .O(N__27203),
            .I(N__27196));
    InMux I__4487 (
            .O(N__27202),
            .I(N__27193));
    Odrv4 I__4486 (
            .O(N__27199),
            .I(\nx.n2802 ));
    Odrv12 I__4485 (
            .O(N__27196),
            .I(\nx.n2802 ));
    LocalMux I__4484 (
            .O(N__27193),
            .I(\nx.n2802 ));
    InMux I__4483 (
            .O(N__27186),
            .I(N__27183));
    LocalMux I__4482 (
            .O(N__27183),
            .I(\nx.n2869 ));
    InMux I__4481 (
            .O(N__27180),
            .I(bfn_6_22_0_));
    InMux I__4480 (
            .O(N__27177),
            .I(\nx.n10821 ));
    CascadeMux I__4479 (
            .O(N__27174),
            .I(N__27170));
    InMux I__4478 (
            .O(N__27173),
            .I(N__27167));
    InMux I__4477 (
            .O(N__27170),
            .I(N__27164));
    LocalMux I__4476 (
            .O(N__27167),
            .I(N__27160));
    LocalMux I__4475 (
            .O(N__27164),
            .I(N__27157));
    InMux I__4474 (
            .O(N__27163),
            .I(N__27154));
    Odrv4 I__4473 (
            .O(N__27160),
            .I(\nx.n2800 ));
    Odrv4 I__4472 (
            .O(N__27157),
            .I(\nx.n2800 ));
    LocalMux I__4471 (
            .O(N__27154),
            .I(\nx.n2800 ));
    CascadeMux I__4470 (
            .O(N__27147),
            .I(N__27144));
    InMux I__4469 (
            .O(N__27144),
            .I(N__27141));
    LocalMux I__4468 (
            .O(N__27141),
            .I(N__27138));
    Odrv4 I__4467 (
            .O(N__27138),
            .I(\nx.n2867 ));
    InMux I__4466 (
            .O(N__27135),
            .I(\nx.n10822 ));
    CascadeMux I__4465 (
            .O(N__27132),
            .I(N__27128));
    InMux I__4464 (
            .O(N__27131),
            .I(N__27125));
    InMux I__4463 (
            .O(N__27128),
            .I(N__27122));
    LocalMux I__4462 (
            .O(N__27125),
            .I(N__27116));
    LocalMux I__4461 (
            .O(N__27122),
            .I(N__27116));
    InMux I__4460 (
            .O(N__27121),
            .I(N__27113));
    Odrv4 I__4459 (
            .O(N__27116),
            .I(\nx.n2799 ));
    LocalMux I__4458 (
            .O(N__27113),
            .I(\nx.n2799 ));
    InMux I__4457 (
            .O(N__27108),
            .I(N__27105));
    LocalMux I__4456 (
            .O(N__27105),
            .I(\nx.n2866 ));
    InMux I__4455 (
            .O(N__27102),
            .I(\nx.n10823 ));
    CascadeMux I__4454 (
            .O(N__27099),
            .I(N__27096));
    InMux I__4453 (
            .O(N__27096),
            .I(N__27091));
    InMux I__4452 (
            .O(N__27095),
            .I(N__27088));
    InMux I__4451 (
            .O(N__27094),
            .I(N__27085));
    LocalMux I__4450 (
            .O(N__27091),
            .I(N__27082));
    LocalMux I__4449 (
            .O(N__27088),
            .I(N__27079));
    LocalMux I__4448 (
            .O(N__27085),
            .I(\nx.n2798 ));
    Odrv4 I__4447 (
            .O(N__27082),
            .I(\nx.n2798 ));
    Odrv4 I__4446 (
            .O(N__27079),
            .I(\nx.n2798 ));
    InMux I__4445 (
            .O(N__27072),
            .I(N__27069));
    LocalMux I__4444 (
            .O(N__27069),
            .I(N__27066));
    Odrv4 I__4443 (
            .O(N__27066),
            .I(\nx.n2865 ));
    InMux I__4442 (
            .O(N__27063),
            .I(\nx.n10824 ));
    CascadeMux I__4441 (
            .O(N__27060),
            .I(N__27056));
    InMux I__4440 (
            .O(N__27059),
            .I(N__27053));
    InMux I__4439 (
            .O(N__27056),
            .I(N__27050));
    LocalMux I__4438 (
            .O(N__27053),
            .I(N__27045));
    LocalMux I__4437 (
            .O(N__27050),
            .I(N__27045));
    Odrv4 I__4436 (
            .O(N__27045),
            .I(\nx.n2797 ));
    InMux I__4435 (
            .O(N__27042),
            .I(N__27039));
    LocalMux I__4434 (
            .O(N__27039),
            .I(\nx.n2864 ));
    InMux I__4433 (
            .O(N__27036),
            .I(\nx.n10825 ));
    InMux I__4432 (
            .O(N__27033),
            .I(\nx.n10826 ));
    InMux I__4431 (
            .O(N__27030),
            .I(bfn_6_21_0_));
    CascadeMux I__4430 (
            .O(N__27027),
            .I(N__27024));
    InMux I__4429 (
            .O(N__27024),
            .I(N__27021));
    LocalMux I__4428 (
            .O(N__27021),
            .I(N__27017));
    CascadeMux I__4427 (
            .O(N__27020),
            .I(N__27014));
    Span4Mux_h I__4426 (
            .O(N__27017),
            .I(N__27011));
    InMux I__4425 (
            .O(N__27014),
            .I(N__27008));
    Odrv4 I__4424 (
            .O(N__27011),
            .I(\nx.n2809 ));
    LocalMux I__4423 (
            .O(N__27008),
            .I(\nx.n2809 ));
    InMux I__4422 (
            .O(N__27003),
            .I(N__27000));
    LocalMux I__4421 (
            .O(N__27000),
            .I(N__26997));
    Span12Mux_s11_v I__4420 (
            .O(N__26997),
            .I(N__26994));
    Odrv12 I__4419 (
            .O(N__26994),
            .I(\nx.n2876 ));
    InMux I__4418 (
            .O(N__26991),
            .I(\nx.n10813 ));
    CascadeMux I__4417 (
            .O(N__26988),
            .I(N__26983));
    InMux I__4416 (
            .O(N__26987),
            .I(N__26978));
    InMux I__4415 (
            .O(N__26986),
            .I(N__26978));
    InMux I__4414 (
            .O(N__26983),
            .I(N__26975));
    LocalMux I__4413 (
            .O(N__26978),
            .I(\nx.n2808 ));
    LocalMux I__4412 (
            .O(N__26975),
            .I(\nx.n2808 ));
    CascadeMux I__4411 (
            .O(N__26970),
            .I(N__26967));
    InMux I__4410 (
            .O(N__26967),
            .I(N__26964));
    LocalMux I__4409 (
            .O(N__26964),
            .I(\nx.n2875 ));
    InMux I__4408 (
            .O(N__26961),
            .I(\nx.n10814 ));
    CascadeMux I__4407 (
            .O(N__26958),
            .I(N__26954));
    InMux I__4406 (
            .O(N__26957),
            .I(N__26950));
    InMux I__4405 (
            .O(N__26954),
            .I(N__26947));
    CascadeMux I__4404 (
            .O(N__26953),
            .I(N__26944));
    LocalMux I__4403 (
            .O(N__26950),
            .I(N__26939));
    LocalMux I__4402 (
            .O(N__26947),
            .I(N__26939));
    InMux I__4401 (
            .O(N__26944),
            .I(N__26936));
    Odrv4 I__4400 (
            .O(N__26939),
            .I(\nx.n2807 ));
    LocalMux I__4399 (
            .O(N__26936),
            .I(\nx.n2807 ));
    InMux I__4398 (
            .O(N__26931),
            .I(N__26928));
    LocalMux I__4397 (
            .O(N__26928),
            .I(\nx.n2874 ));
    InMux I__4396 (
            .O(N__26925),
            .I(\nx.n10815 ));
    InMux I__4395 (
            .O(N__26922),
            .I(\nx.n10816 ));
    CascadeMux I__4394 (
            .O(N__26919),
            .I(N__26915));
    CascadeMux I__4393 (
            .O(N__26918),
            .I(N__26912));
    InMux I__4392 (
            .O(N__26915),
            .I(N__26908));
    InMux I__4391 (
            .O(N__26912),
            .I(N__26905));
    InMux I__4390 (
            .O(N__26911),
            .I(N__26902));
    LocalMux I__4389 (
            .O(N__26908),
            .I(N__26897));
    LocalMux I__4388 (
            .O(N__26905),
            .I(N__26897));
    LocalMux I__4387 (
            .O(N__26902),
            .I(\nx.n2805 ));
    Odrv4 I__4386 (
            .O(N__26897),
            .I(\nx.n2805 ));
    InMux I__4385 (
            .O(N__26892),
            .I(N__26889));
    LocalMux I__4384 (
            .O(N__26889),
            .I(\nx.n2872 ));
    InMux I__4383 (
            .O(N__26886),
            .I(\nx.n10817 ));
    InMux I__4382 (
            .O(N__26883),
            .I(\nx.n10818 ));
    InMux I__4381 (
            .O(N__26880),
            .I(N__26877));
    LocalMux I__4380 (
            .O(N__26877),
            .I(\nx.n29_adj_607 ));
    CascadeMux I__4379 (
            .O(N__26874),
            .I(\nx.n37_adj_608_cascade_ ));
    InMux I__4378 (
            .O(N__26871),
            .I(N__26868));
    LocalMux I__4377 (
            .O(N__26868),
            .I(\nx.n40_adj_609 ));
    CascadeMux I__4376 (
            .O(N__26865),
            .I(\nx.n42_cascade_ ));
    CascadeMux I__4375 (
            .O(N__26862),
            .I(\nx.n2720_cascade_ ));
    CascadeMux I__4374 (
            .O(N__26859),
            .I(\nx.n2797_cascade_ ));
    CascadeMux I__4373 (
            .O(N__26856),
            .I(\nx.n2700_cascade_ ));
    CascadeMux I__4372 (
            .O(N__26853),
            .I(\nx.n2801_cascade_ ));
    CascadeMux I__4371 (
            .O(N__26850),
            .I(N__26845));
    InMux I__4370 (
            .O(N__26849),
            .I(N__26842));
    InMux I__4369 (
            .O(N__26848),
            .I(N__26839));
    InMux I__4368 (
            .O(N__26845),
            .I(N__26836));
    LocalMux I__4367 (
            .O(N__26842),
            .I(\nx.n1407 ));
    LocalMux I__4366 (
            .O(N__26839),
            .I(\nx.n1407 ));
    LocalMux I__4365 (
            .O(N__26836),
            .I(\nx.n1407 ));
    CascadeMux I__4364 (
            .O(N__26829),
            .I(N__26826));
    InMux I__4363 (
            .O(N__26826),
            .I(N__26823));
    LocalMux I__4362 (
            .O(N__26823),
            .I(N__26820));
    Odrv4 I__4361 (
            .O(N__26820),
            .I(\nx.n1474 ));
    CascadeMux I__4360 (
            .O(N__26817),
            .I(\nx.n1506_cascade_ ));
    InMux I__4359 (
            .O(N__26814),
            .I(N__26811));
    LocalMux I__4358 (
            .O(N__26811),
            .I(\nx.n18_adj_632 ));
    InMux I__4357 (
            .O(N__26808),
            .I(N__26805));
    LocalMux I__4356 (
            .O(N__26805),
            .I(N__26802));
    Odrv4 I__4355 (
            .O(N__26802),
            .I(\nx.n1475 ));
    CascadeMux I__4354 (
            .O(N__26799),
            .I(N__26796));
    InMux I__4353 (
            .O(N__26796),
            .I(N__26793));
    LocalMux I__4352 (
            .O(N__26793),
            .I(N__26788));
    InMux I__4351 (
            .O(N__26792),
            .I(N__26785));
    CascadeMux I__4350 (
            .O(N__26791),
            .I(N__26782));
    Span4Mux_s2_v I__4349 (
            .O(N__26788),
            .I(N__26779));
    LocalMux I__4348 (
            .O(N__26785),
            .I(N__26776));
    InMux I__4347 (
            .O(N__26782),
            .I(N__26773));
    Odrv4 I__4346 (
            .O(N__26779),
            .I(\nx.n1408 ));
    Odrv4 I__4345 (
            .O(N__26776),
            .I(\nx.n1408 ));
    LocalMux I__4344 (
            .O(N__26773),
            .I(\nx.n1408 ));
    InMux I__4343 (
            .O(N__26766),
            .I(N__26762));
    CascadeMux I__4342 (
            .O(N__26765),
            .I(N__26758));
    LocalMux I__4341 (
            .O(N__26762),
            .I(N__26755));
    InMux I__4340 (
            .O(N__26761),
            .I(N__26752));
    InMux I__4339 (
            .O(N__26758),
            .I(N__26749));
    Odrv4 I__4338 (
            .O(N__26755),
            .I(\nx.n1401 ));
    LocalMux I__4337 (
            .O(N__26752),
            .I(\nx.n1401 ));
    LocalMux I__4336 (
            .O(N__26749),
            .I(\nx.n1401 ));
    InMux I__4335 (
            .O(N__26742),
            .I(N__26739));
    LocalMux I__4334 (
            .O(N__26739),
            .I(N__26736));
    Odrv4 I__4333 (
            .O(N__26736),
            .I(\nx.n1468 ));
    InMux I__4332 (
            .O(N__26733),
            .I(N__26730));
    LocalMux I__4331 (
            .O(N__26730),
            .I(N__26727));
    Span4Mux_s1_v I__4330 (
            .O(N__26727),
            .I(N__26724));
    Odrv4 I__4329 (
            .O(N__26724),
            .I(\nx.n1472 ));
    CascadeMux I__4328 (
            .O(N__26721),
            .I(N__26716));
    InMux I__4327 (
            .O(N__26720),
            .I(N__26713));
    InMux I__4326 (
            .O(N__26719),
            .I(N__26710));
    InMux I__4325 (
            .O(N__26716),
            .I(N__26707));
    LocalMux I__4324 (
            .O(N__26713),
            .I(\nx.n1405 ));
    LocalMux I__4323 (
            .O(N__26710),
            .I(\nx.n1405 ));
    LocalMux I__4322 (
            .O(N__26707),
            .I(\nx.n1405 ));
    InMux I__4321 (
            .O(N__26700),
            .I(N__26697));
    LocalMux I__4320 (
            .O(N__26697),
            .I(N__26694));
    Span4Mux_s1_v I__4319 (
            .O(N__26694),
            .I(N__26691));
    Odrv4 I__4318 (
            .O(N__26691),
            .I(\nx.n1473 ));
    CascadeMux I__4317 (
            .O(N__26688),
            .I(N__26685));
    InMux I__4316 (
            .O(N__26685),
            .I(N__26681));
    CascadeMux I__4315 (
            .O(N__26684),
            .I(N__26678));
    LocalMux I__4314 (
            .O(N__26681),
            .I(N__26674));
    InMux I__4313 (
            .O(N__26678),
            .I(N__26671));
    CascadeMux I__4312 (
            .O(N__26677),
            .I(N__26668));
    Span4Mux_s2_v I__4311 (
            .O(N__26674),
            .I(N__26665));
    LocalMux I__4310 (
            .O(N__26671),
            .I(N__26662));
    InMux I__4309 (
            .O(N__26668),
            .I(N__26659));
    Odrv4 I__4308 (
            .O(N__26665),
            .I(\nx.n1406 ));
    Odrv4 I__4307 (
            .O(N__26662),
            .I(\nx.n1406 ));
    LocalMux I__4306 (
            .O(N__26659),
            .I(\nx.n1406 ));
    CascadeMux I__4305 (
            .O(N__26652),
            .I(N__26648));
    InMux I__4304 (
            .O(N__26651),
            .I(N__26643));
    InMux I__4303 (
            .O(N__26648),
            .I(N__26640));
    InMux I__4302 (
            .O(N__26647),
            .I(N__26637));
    InMux I__4301 (
            .O(N__26646),
            .I(N__26634));
    LocalMux I__4300 (
            .O(N__26643),
            .I(N__26629));
    LocalMux I__4299 (
            .O(N__26640),
            .I(N__26629));
    LocalMux I__4298 (
            .O(N__26637),
            .I(N__26626));
    LocalMux I__4297 (
            .O(N__26634),
            .I(N__26621));
    Span4Mux_v I__4296 (
            .O(N__26629),
            .I(N__26621));
    Span4Mux_v I__4295 (
            .O(N__26626),
            .I(N__26618));
    Odrv4 I__4294 (
            .O(N__26621),
            .I(neopxl_color_15));
    Odrv4 I__4293 (
            .O(N__26618),
            .I(neopxl_color_15));
    CascadeMux I__4292 (
            .O(N__26613),
            .I(\nx.n9618_cascade_ ));
    CascadeMux I__4291 (
            .O(N__26610),
            .I(N__26606));
    InMux I__4290 (
            .O(N__26609),
            .I(N__26603));
    InMux I__4289 (
            .O(N__26606),
            .I(N__26600));
    LocalMux I__4288 (
            .O(N__26603),
            .I(\nx.n608 ));
    LocalMux I__4287 (
            .O(N__26600),
            .I(\nx.n608 ));
    CascadeMux I__4286 (
            .O(N__26595),
            .I(\nx.n11738_cascade_ ));
    InMux I__4285 (
            .O(N__26592),
            .I(N__26586));
    InMux I__4284 (
            .O(N__26591),
            .I(N__26586));
    LocalMux I__4283 (
            .O(N__26586),
            .I(\nx.n708 ));
    CascadeMux I__4282 (
            .O(N__26583),
            .I(\nx.n739_cascade_ ));
    InMux I__4281 (
            .O(N__26580),
            .I(N__26577));
    LocalMux I__4280 (
            .O(N__26577),
            .I(\nx.n11738 ));
    InMux I__4279 (
            .O(N__26574),
            .I(N__26567));
    InMux I__4278 (
            .O(N__26573),
            .I(N__26567));
    InMux I__4277 (
            .O(N__26572),
            .I(N__26564));
    LocalMux I__4276 (
            .O(N__26567),
            .I(\nx.n807 ));
    LocalMux I__4275 (
            .O(N__26564),
            .I(\nx.n807 ));
    CascadeMux I__4274 (
            .O(N__26559),
            .I(N__26554));
    CascadeMux I__4273 (
            .O(N__26558),
            .I(N__26549));
    InMux I__4272 (
            .O(N__26557),
            .I(N__26545));
    InMux I__4271 (
            .O(N__26554),
            .I(N__26542));
    InMux I__4270 (
            .O(N__26553),
            .I(N__26537));
    InMux I__4269 (
            .O(N__26552),
            .I(N__26537));
    InMux I__4268 (
            .O(N__26549),
            .I(N__26532));
    InMux I__4267 (
            .O(N__26548),
            .I(N__26532));
    LocalMux I__4266 (
            .O(N__26545),
            .I(\nx.bit_ctr_31 ));
    LocalMux I__4265 (
            .O(N__26542),
            .I(\nx.bit_ctr_31 ));
    LocalMux I__4264 (
            .O(N__26537),
            .I(\nx.bit_ctr_31 ));
    LocalMux I__4263 (
            .O(N__26532),
            .I(\nx.bit_ctr_31 ));
    CascadeMux I__4262 (
            .O(N__26523),
            .I(N__26519));
    InMux I__4261 (
            .O(N__26522),
            .I(N__26515));
    InMux I__4260 (
            .O(N__26519),
            .I(N__26510));
    InMux I__4259 (
            .O(N__26518),
            .I(N__26510));
    LocalMux I__4258 (
            .O(N__26515),
            .I(\nx.n9618 ));
    LocalMux I__4257 (
            .O(N__26510),
            .I(\nx.n9618 ));
    CascadeMux I__4256 (
            .O(N__26505),
            .I(N__26501));
    InMux I__4255 (
            .O(N__26504),
            .I(N__26494));
    InMux I__4254 (
            .O(N__26501),
            .I(N__26491));
    InMux I__4253 (
            .O(N__26500),
            .I(N__26482));
    InMux I__4252 (
            .O(N__26499),
            .I(N__26482));
    InMux I__4251 (
            .O(N__26498),
            .I(N__26482));
    InMux I__4250 (
            .O(N__26497),
            .I(N__26482));
    LocalMux I__4249 (
            .O(N__26494),
            .I(\nx.bit_ctr_29 ));
    LocalMux I__4248 (
            .O(N__26491),
            .I(\nx.bit_ctr_29 ));
    LocalMux I__4247 (
            .O(N__26482),
            .I(\nx.bit_ctr_29 ));
    CascadeMux I__4246 (
            .O(N__26475),
            .I(\nx.n11771_cascade_ ));
    InMux I__4245 (
            .O(N__26472),
            .I(N__26469));
    LocalMux I__4244 (
            .O(N__26469),
            .I(N__26466));
    Odrv4 I__4243 (
            .O(N__26466),
            .I(\nx.n1470 ));
    CascadeMux I__4242 (
            .O(N__26463),
            .I(N__26459));
    CascadeMux I__4241 (
            .O(N__26462),
            .I(N__26456));
    InMux I__4240 (
            .O(N__26459),
            .I(N__26452));
    InMux I__4239 (
            .O(N__26456),
            .I(N__26449));
    InMux I__4238 (
            .O(N__26455),
            .I(N__26446));
    LocalMux I__4237 (
            .O(N__26452),
            .I(\nx.n1403 ));
    LocalMux I__4236 (
            .O(N__26449),
            .I(\nx.n1403 ));
    LocalMux I__4235 (
            .O(N__26446),
            .I(\nx.n1403 ));
    InMux I__4234 (
            .O(N__26439),
            .I(N__26434));
    CascadeMux I__4233 (
            .O(N__26438),
            .I(N__26429));
    InMux I__4232 (
            .O(N__26437),
            .I(N__26425));
    LocalMux I__4231 (
            .O(N__26434),
            .I(N__26422));
    InMux I__4230 (
            .O(N__26433),
            .I(N__26413));
    InMux I__4229 (
            .O(N__26432),
            .I(N__26413));
    InMux I__4228 (
            .O(N__26429),
            .I(N__26413));
    InMux I__4227 (
            .O(N__26428),
            .I(N__26413));
    LocalMux I__4226 (
            .O(N__26425),
            .I(\nx.bit_ctr_30 ));
    Odrv4 I__4225 (
            .O(N__26422),
            .I(\nx.bit_ctr_30 ));
    LocalMux I__4224 (
            .O(N__26413),
            .I(\nx.bit_ctr_30 ));
    CascadeMux I__4223 (
            .O(N__26406),
            .I(N__26403));
    InMux I__4222 (
            .O(N__26403),
            .I(N__26400));
    LocalMux I__4221 (
            .O(N__26400),
            .I(N__26397));
    Span4Mux_h I__4220 (
            .O(N__26397),
            .I(N__26394));
    Odrv4 I__4219 (
            .O(N__26394),
            .I(\nx.n48_adj_704 ));
    InMux I__4218 (
            .O(N__26391),
            .I(N__26386));
    InMux I__4217 (
            .O(N__26390),
            .I(N__26381));
    InMux I__4216 (
            .O(N__26389),
            .I(N__26381));
    LocalMux I__4215 (
            .O(N__26386),
            .I(N__26378));
    LocalMux I__4214 (
            .O(N__26381),
            .I(\nx.n1008 ));
    Odrv4 I__4213 (
            .O(N__26378),
            .I(\nx.n1008 ));
    CascadeMux I__4212 (
            .O(N__26373),
            .I(\nx.n7084_cascade_ ));
    CascadeMux I__4211 (
            .O(N__26370),
            .I(\nx.n838_cascade_ ));
    CascadeMux I__4210 (
            .O(N__26367),
            .I(\nx.n12595_cascade_ ));
    CascadeMux I__4209 (
            .O(N__26364),
            .I(\nx.n11617_cascade_ ));
    InMux I__4208 (
            .O(N__26361),
            .I(N__26358));
    LocalMux I__4207 (
            .O(N__26358),
            .I(\nx.n1076 ));
    CascadeMux I__4206 (
            .O(N__26355),
            .I(\nx.n1037_cascade_ ));
    CascadeMux I__4205 (
            .O(N__26352),
            .I(N__26348));
    CascadeMux I__4204 (
            .O(N__26351),
            .I(N__26344));
    InMux I__4203 (
            .O(N__26348),
            .I(N__26341));
    InMux I__4202 (
            .O(N__26347),
            .I(N__26338));
    InMux I__4201 (
            .O(N__26344),
            .I(N__26335));
    LocalMux I__4200 (
            .O(N__26341),
            .I(N__26332));
    LocalMux I__4199 (
            .O(N__26338),
            .I(N__26327));
    LocalMux I__4198 (
            .O(N__26335),
            .I(N__26327));
    Span4Mux_h I__4197 (
            .O(N__26332),
            .I(N__26324));
    Span4Mux_h I__4196 (
            .O(N__26327),
            .I(N__26321));
    Odrv4 I__4195 (
            .O(N__26324),
            .I(\nx.n1108 ));
    Odrv4 I__4194 (
            .O(N__26321),
            .I(\nx.n1108 ));
    CascadeMux I__4193 (
            .O(N__26316),
            .I(N__26312));
    InMux I__4192 (
            .O(N__26315),
            .I(N__26309));
    InMux I__4191 (
            .O(N__26312),
            .I(N__26306));
    LocalMux I__4190 (
            .O(N__26309),
            .I(\nx.n1007 ));
    LocalMux I__4189 (
            .O(N__26306),
            .I(\nx.n1007 ));
    InMux I__4188 (
            .O(N__26301),
            .I(N__26298));
    LocalMux I__4187 (
            .O(N__26298),
            .I(N__26295));
    Odrv4 I__4186 (
            .O(N__26295),
            .I(\nx.n1074 ));
    CascadeMux I__4185 (
            .O(N__26292),
            .I(N__26288));
    InMux I__4184 (
            .O(N__26291),
            .I(N__26285));
    InMux I__4183 (
            .O(N__26288),
            .I(N__26281));
    LocalMux I__4182 (
            .O(N__26285),
            .I(N__26278));
    InMux I__4181 (
            .O(N__26284),
            .I(N__26275));
    LocalMux I__4180 (
            .O(N__26281),
            .I(N__26272));
    Span4Mux_h I__4179 (
            .O(N__26278),
            .I(N__26269));
    LocalMux I__4178 (
            .O(N__26275),
            .I(N__26266));
    Span4Mux_h I__4177 (
            .O(N__26272),
            .I(N__26263));
    Span4Mux_s2_v I__4176 (
            .O(N__26269),
            .I(N__26258));
    Span4Mux_h I__4175 (
            .O(N__26266),
            .I(N__26258));
    Odrv4 I__4174 (
            .O(N__26263),
            .I(\nx.n1106 ));
    Odrv4 I__4173 (
            .O(N__26258),
            .I(\nx.n1106 ));
    CascadeMux I__4172 (
            .O(N__26253),
            .I(N__26250));
    InMux I__4171 (
            .O(N__26250),
            .I(N__26246));
    InMux I__4170 (
            .O(N__26249),
            .I(N__26243));
    LocalMux I__4169 (
            .O(N__26246),
            .I(N__26240));
    LocalMux I__4168 (
            .O(N__26243),
            .I(\nx.n1009 ));
    Odrv4 I__4167 (
            .O(N__26240),
            .I(\nx.n1009 ));
    CascadeMux I__4166 (
            .O(N__26235),
            .I(N__26232));
    InMux I__4165 (
            .O(N__26232),
            .I(N__26227));
    InMux I__4164 (
            .O(N__26231),
            .I(N__26224));
    InMux I__4163 (
            .O(N__26230),
            .I(N__26220));
    LocalMux I__4162 (
            .O(N__26227),
            .I(N__26216));
    LocalMux I__4161 (
            .O(N__26224),
            .I(N__26213));
    InMux I__4160 (
            .O(N__26223),
            .I(N__26210));
    LocalMux I__4159 (
            .O(N__26220),
            .I(N__26207));
    InMux I__4158 (
            .O(N__26219),
            .I(N__26204));
    Span4Mux_v I__4157 (
            .O(N__26216),
            .I(N__26199));
    Span4Mux_v I__4156 (
            .O(N__26213),
            .I(N__26199));
    LocalMux I__4155 (
            .O(N__26210),
            .I(N__26196));
    Span4Mux_v I__4154 (
            .O(N__26207),
            .I(N__26193));
    LocalMux I__4153 (
            .O(N__26204),
            .I(\nx.bit_ctr_25 ));
    Odrv4 I__4152 (
            .O(N__26199),
            .I(\nx.bit_ctr_25 ));
    Odrv4 I__4151 (
            .O(N__26196),
            .I(\nx.bit_ctr_25 ));
    Odrv4 I__4150 (
            .O(N__26193),
            .I(\nx.bit_ctr_25 ));
    CascadeMux I__4149 (
            .O(N__26184),
            .I(\nx.n1009_cascade_ ));
    InMux I__4148 (
            .O(N__26181),
            .I(N__26178));
    LocalMux I__4147 (
            .O(N__26178),
            .I(\nx.n7_adj_616 ));
    InMux I__4146 (
            .O(N__26175),
            .I(N__26172));
    LocalMux I__4145 (
            .O(N__26172),
            .I(N__26166));
    InMux I__4144 (
            .O(N__26171),
            .I(N__26163));
    InMux I__4143 (
            .O(N__26170),
            .I(N__26159));
    InMux I__4142 (
            .O(N__26169),
            .I(N__26156));
    Span4Mux_v I__4141 (
            .O(N__26166),
            .I(N__26153));
    LocalMux I__4140 (
            .O(N__26163),
            .I(N__26150));
    InMux I__4139 (
            .O(N__26162),
            .I(N__26147));
    LocalMux I__4138 (
            .O(N__26159),
            .I(\nx.bit_ctr_5 ));
    LocalMux I__4137 (
            .O(N__26156),
            .I(\nx.bit_ctr_5 ));
    Odrv4 I__4136 (
            .O(N__26153),
            .I(\nx.bit_ctr_5 ));
    Odrv12 I__4135 (
            .O(N__26150),
            .I(\nx.bit_ctr_5 ));
    LocalMux I__4134 (
            .O(N__26147),
            .I(\nx.bit_ctr_5 ));
    InMux I__4133 (
            .O(N__26136),
            .I(N__26131));
    InMux I__4132 (
            .O(N__26135),
            .I(N__26128));
    InMux I__4131 (
            .O(N__26134),
            .I(N__26125));
    LocalMux I__4130 (
            .O(N__26131),
            .I(N__26120));
    LocalMux I__4129 (
            .O(N__26128),
            .I(N__26120));
    LocalMux I__4128 (
            .O(N__26125),
            .I(N__26115));
    Span4Mux_v I__4127 (
            .O(N__26120),
            .I(N__26112));
    InMux I__4126 (
            .O(N__26119),
            .I(N__26109));
    InMux I__4125 (
            .O(N__26118),
            .I(N__26106));
    Span4Mux_v I__4124 (
            .O(N__26115),
            .I(N__26103));
    Span4Mux_v I__4123 (
            .O(N__26112),
            .I(N__26100));
    LocalMux I__4122 (
            .O(N__26109),
            .I(\nx.bit_ctr_6 ));
    LocalMux I__4121 (
            .O(N__26106),
            .I(\nx.bit_ctr_6 ));
    Odrv4 I__4120 (
            .O(N__26103),
            .I(\nx.bit_ctr_6 ));
    Odrv4 I__4119 (
            .O(N__26100),
            .I(\nx.bit_ctr_6 ));
    InMux I__4118 (
            .O(N__26091),
            .I(N__26088));
    LocalMux I__4117 (
            .O(N__26088),
            .I(N__26085));
    Odrv12 I__4116 (
            .O(N__26085),
            .I(\nx.n44_adj_708 ));
    CascadeMux I__4115 (
            .O(N__26082),
            .I(N__26079));
    InMux I__4114 (
            .O(N__26079),
            .I(N__26076));
    LocalMux I__4113 (
            .O(N__26076),
            .I(N__26072));
    InMux I__4112 (
            .O(N__26075),
            .I(N__26069));
    Odrv4 I__4111 (
            .O(N__26072),
            .I(\nx.n1005 ));
    LocalMux I__4110 (
            .O(N__26069),
            .I(\nx.n1005 ));
    InMux I__4109 (
            .O(N__26064),
            .I(N__26061));
    LocalMux I__4108 (
            .O(N__26061),
            .I(N__26058));
    Odrv4 I__4107 (
            .O(N__26058),
            .I(\nx.n1072 ));
    CascadeMux I__4106 (
            .O(N__26055),
            .I(\nx.n1005_cascade_ ));
    InMux I__4105 (
            .O(N__26052),
            .I(N__26049));
    LocalMux I__4104 (
            .O(N__26049),
            .I(N__26041));
    InMux I__4103 (
            .O(N__26048),
            .I(N__26038));
    InMux I__4102 (
            .O(N__26047),
            .I(N__26033));
    InMux I__4101 (
            .O(N__26046),
            .I(N__26033));
    InMux I__4100 (
            .O(N__26045),
            .I(N__26028));
    InMux I__4099 (
            .O(N__26044),
            .I(N__26028));
    Span4Mux_h I__4098 (
            .O(N__26041),
            .I(N__26025));
    LocalMux I__4097 (
            .O(N__26038),
            .I(\nx.n1037 ));
    LocalMux I__4096 (
            .O(N__26033),
            .I(\nx.n1037 ));
    LocalMux I__4095 (
            .O(N__26028),
            .I(\nx.n1037 ));
    Odrv4 I__4094 (
            .O(N__26025),
            .I(\nx.n1037 ));
    CascadeMux I__4093 (
            .O(N__26016),
            .I(N__26013));
    InMux I__4092 (
            .O(N__26013),
            .I(N__26008));
    InMux I__4091 (
            .O(N__26012),
            .I(N__26005));
    InMux I__4090 (
            .O(N__26011),
            .I(N__26002));
    LocalMux I__4089 (
            .O(N__26008),
            .I(N__25999));
    LocalMux I__4088 (
            .O(N__26005),
            .I(N__25994));
    LocalMux I__4087 (
            .O(N__26002),
            .I(N__25994));
    Span4Mux_h I__4086 (
            .O(N__25999),
            .I(N__25991));
    Span4Mux_h I__4085 (
            .O(N__25994),
            .I(N__25988));
    Odrv4 I__4084 (
            .O(N__25991),
            .I(\nx.n1104 ));
    Odrv4 I__4083 (
            .O(N__25988),
            .I(\nx.n1104 ));
    InMux I__4082 (
            .O(N__25983),
            .I(\nx.n10472 ));
    InMux I__4081 (
            .O(N__25980),
            .I(\nx.n10473 ));
    CascadeMux I__4080 (
            .O(N__25977),
            .I(N__25973));
    InMux I__4079 (
            .O(N__25976),
            .I(N__25970));
    InMux I__4078 (
            .O(N__25973),
            .I(N__25967));
    LocalMux I__4077 (
            .O(N__25970),
            .I(N__25964));
    LocalMux I__4076 (
            .O(N__25967),
            .I(N__25959));
    Span4Mux_s1_h I__4075 (
            .O(N__25964),
            .I(N__25959));
    Span4Mux_v I__4074 (
            .O(N__25959),
            .I(N__25956));
    Odrv4 I__4073 (
            .O(N__25956),
            .I(\nx.n1103 ));
    InMux I__4072 (
            .O(N__25953),
            .I(N__25950));
    LocalMux I__4071 (
            .O(N__25950),
            .I(N__25947));
    Span4Mux_h I__4070 (
            .O(N__25947),
            .I(N__25944));
    Odrv4 I__4069 (
            .O(N__25944),
            .I(\nx.n46_adj_705 ));
    InMux I__4068 (
            .O(N__25941),
            .I(N__25938));
    LocalMux I__4067 (
            .O(N__25938),
            .I(\nx.n1075 ));
    CascadeMux I__4066 (
            .O(N__25935),
            .I(N__25932));
    InMux I__4065 (
            .O(N__25932),
            .I(N__25927));
    InMux I__4064 (
            .O(N__25931),
            .I(N__25924));
    CascadeMux I__4063 (
            .O(N__25930),
            .I(N__25921));
    LocalMux I__4062 (
            .O(N__25927),
            .I(N__25916));
    LocalMux I__4061 (
            .O(N__25924),
            .I(N__25916));
    InMux I__4060 (
            .O(N__25921),
            .I(N__25913));
    Span4Mux_s3_v I__4059 (
            .O(N__25916),
            .I(N__25908));
    LocalMux I__4058 (
            .O(N__25913),
            .I(N__25908));
    Span4Mux_h I__4057 (
            .O(N__25908),
            .I(N__25905));
    Odrv4 I__4056 (
            .O(N__25905),
            .I(\nx.n1107 ));
    InMux I__4055 (
            .O(N__25902),
            .I(N__25899));
    LocalMux I__4054 (
            .O(N__25899),
            .I(\nx.n1073 ));
    CascadeMux I__4053 (
            .O(N__25896),
            .I(N__25891));
    InMux I__4052 (
            .O(N__25895),
            .I(N__25888));
    InMux I__4051 (
            .O(N__25894),
            .I(N__25885));
    InMux I__4050 (
            .O(N__25891),
            .I(N__25882));
    LocalMux I__4049 (
            .O(N__25888),
            .I(N__25875));
    LocalMux I__4048 (
            .O(N__25885),
            .I(N__25875));
    LocalMux I__4047 (
            .O(N__25882),
            .I(N__25875));
    Span4Mux_v I__4046 (
            .O(N__25875),
            .I(N__25872));
    Odrv4 I__4045 (
            .O(N__25872),
            .I(\nx.n1105 ));
    CascadeMux I__4044 (
            .O(N__25869),
            .I(N__25865));
    InMux I__4043 (
            .O(N__25868),
            .I(N__25862));
    InMux I__4042 (
            .O(N__25865),
            .I(N__25859));
    LocalMux I__4041 (
            .O(N__25862),
            .I(N__25854));
    LocalMux I__4040 (
            .O(N__25859),
            .I(N__25854));
    Span4Mux_v I__4039 (
            .O(N__25854),
            .I(N__25851));
    Odrv4 I__4038 (
            .O(N__25851),
            .I(\nx.n2894 ));
    CascadeMux I__4037 (
            .O(N__25848),
            .I(N__25845));
    InMux I__4036 (
            .O(N__25845),
            .I(N__25842));
    LocalMux I__4035 (
            .O(N__25842),
            .I(N__25838));
    InMux I__4034 (
            .O(N__25841),
            .I(N__25835));
    Span4Mux_h I__4033 (
            .O(N__25838),
            .I(N__25832));
    LocalMux I__4032 (
            .O(N__25835),
            .I(\nx.n2993 ));
    Odrv4 I__4031 (
            .O(N__25832),
            .I(\nx.n2993 ));
    InMux I__4030 (
            .O(N__25827),
            .I(N__25824));
    LocalMux I__4029 (
            .O(N__25824),
            .I(N__25821));
    Span4Mux_h I__4028 (
            .O(N__25821),
            .I(N__25818));
    Odrv4 I__4027 (
            .O(N__25818),
            .I(\nx.n3060 ));
    CascadeMux I__4026 (
            .O(N__25815),
            .I(\nx.n2993_cascade_ ));
    InMux I__4025 (
            .O(N__25812),
            .I(N__25809));
    LocalMux I__4024 (
            .O(N__25809),
            .I(N__25805));
    InMux I__4023 (
            .O(N__25808),
            .I(N__25802));
    Span12Mux_s4_h I__4022 (
            .O(N__25805),
            .I(N__25799));
    LocalMux I__4021 (
            .O(N__25802),
            .I(\nx.n3092 ));
    Odrv12 I__4020 (
            .O(N__25799),
            .I(\nx.n3092 ));
    InMux I__4019 (
            .O(N__25794),
            .I(N__25790));
    InMux I__4018 (
            .O(N__25793),
            .I(N__25787));
    LocalMux I__4017 (
            .O(N__25790),
            .I(N__25784));
    LocalMux I__4016 (
            .O(N__25787),
            .I(N__25780));
    Span4Mux_v I__4015 (
            .O(N__25784),
            .I(N__25777));
    InMux I__4014 (
            .O(N__25783),
            .I(N__25774));
    Span4Mux_h I__4013 (
            .O(N__25780),
            .I(N__25771));
    Odrv4 I__4012 (
            .O(N__25777),
            .I(\nx.n3091 ));
    LocalMux I__4011 (
            .O(N__25774),
            .I(\nx.n3091 ));
    Odrv4 I__4010 (
            .O(N__25771),
            .I(\nx.n3091 ));
    CascadeMux I__4009 (
            .O(N__25764),
            .I(\nx.n3092_cascade_ ));
    InMux I__4008 (
            .O(N__25761),
            .I(N__25758));
    LocalMux I__4007 (
            .O(N__25758),
            .I(N__25755));
    Span4Mux_h I__4006 (
            .O(N__25755),
            .I(N__25752));
    Odrv4 I__4005 (
            .O(N__25752),
            .I(\nx.n46_adj_688 ));
    InMux I__4004 (
            .O(N__25749),
            .I(N__25746));
    LocalMux I__4003 (
            .O(N__25746),
            .I(N__25743));
    Span4Mux_s1_h I__4002 (
            .O(N__25743),
            .I(N__25740));
    Odrv4 I__4001 (
            .O(N__25740),
            .I(\nx.n50 ));
    InMux I__4000 (
            .O(N__25737),
            .I(N__25734));
    LocalMux I__3999 (
            .O(N__25734),
            .I(N__25730));
    InMux I__3998 (
            .O(N__25733),
            .I(N__25726));
    Span4Mux_h I__3997 (
            .O(N__25730),
            .I(N__25723));
    InMux I__3996 (
            .O(N__25729),
            .I(N__25720));
    LocalMux I__3995 (
            .O(N__25726),
            .I(\nx.n3093 ));
    Odrv4 I__3994 (
            .O(N__25723),
            .I(\nx.n3093 ));
    LocalMux I__3993 (
            .O(N__25720),
            .I(\nx.n3093 ));
    InMux I__3992 (
            .O(N__25713),
            .I(N__25710));
    LocalMux I__3991 (
            .O(N__25710),
            .I(\nx.n36_adj_687 ));
    InMux I__3990 (
            .O(N__25707),
            .I(N__25704));
    LocalMux I__3989 (
            .O(N__25704),
            .I(N__25701));
    Span12Mux_s6_v I__3988 (
            .O(N__25701),
            .I(N__25698));
    Odrv12 I__3987 (
            .O(N__25698),
            .I(\nx.n1077 ));
    InMux I__3986 (
            .O(N__25695),
            .I(bfn_5_26_0_));
    InMux I__3985 (
            .O(N__25692),
            .I(\nx.n10468 ));
    InMux I__3984 (
            .O(N__25689),
            .I(\nx.n10469 ));
    InMux I__3983 (
            .O(N__25686),
            .I(\nx.n10470 ));
    InMux I__3982 (
            .O(N__25683),
            .I(\nx.n10471 ));
    InMux I__3981 (
            .O(N__25680),
            .I(N__25677));
    LocalMux I__3980 (
            .O(N__25677),
            .I(\nx.n2959 ));
    InMux I__3979 (
            .O(N__25674),
            .I(\nx.n10854 ));
    CascadeMux I__3978 (
            .O(N__25671),
            .I(N__25668));
    InMux I__3977 (
            .O(N__25668),
            .I(N__25665));
    LocalMux I__3976 (
            .O(N__25665),
            .I(\nx.n2958 ));
    InMux I__3975 (
            .O(N__25662),
            .I(\nx.n10855 ));
    InMux I__3974 (
            .O(N__25659),
            .I(N__25656));
    LocalMux I__3973 (
            .O(N__25656),
            .I(\nx.n2957 ));
    InMux I__3972 (
            .O(N__25653),
            .I(\nx.n10856 ));
    InMux I__3971 (
            .O(N__25650),
            .I(N__25647));
    LocalMux I__3970 (
            .O(N__25647),
            .I(\nx.n2956 ));
    InMux I__3969 (
            .O(N__25644),
            .I(\nx.n10857 ));
    InMux I__3968 (
            .O(N__25641),
            .I(N__25638));
    LocalMux I__3967 (
            .O(N__25638),
            .I(\nx.n2955 ));
    InMux I__3966 (
            .O(N__25635),
            .I(\nx.n10858 ));
    InMux I__3965 (
            .O(N__25632),
            .I(N__25629));
    LocalMux I__3964 (
            .O(N__25629),
            .I(N__25626));
    Odrv4 I__3963 (
            .O(N__25626),
            .I(\nx.n2954 ));
    InMux I__3962 (
            .O(N__25623),
            .I(\nx.n10859 ));
    InMux I__3961 (
            .O(N__25620),
            .I(N__25617));
    LocalMux I__3960 (
            .O(N__25617),
            .I(N__25614));
    Odrv4 I__3959 (
            .O(N__25614),
            .I(\nx.n2953 ));
    InMux I__3958 (
            .O(N__25611),
            .I(bfn_5_25_0_));
    InMux I__3957 (
            .O(N__25608),
            .I(\nx.n10861 ));
    InMux I__3956 (
            .O(N__25605),
            .I(N__25602));
    LocalMux I__3955 (
            .O(N__25602),
            .I(N__25598));
    InMux I__3954 (
            .O(N__25601),
            .I(N__25595));
    Span4Mux_v I__3953 (
            .O(N__25598),
            .I(N__25592));
    LocalMux I__3952 (
            .O(N__25595),
            .I(N__25589));
    Odrv4 I__3951 (
            .O(N__25592),
            .I(\nx.n2984 ));
    Odrv4 I__3950 (
            .O(N__25589),
            .I(\nx.n2984 ));
    InMux I__3949 (
            .O(N__25584),
            .I(N__25581));
    LocalMux I__3948 (
            .O(N__25581),
            .I(\nx.n2961 ));
    CascadeMux I__3947 (
            .O(N__25578),
            .I(N__25575));
    InMux I__3946 (
            .O(N__25575),
            .I(N__25572));
    LocalMux I__3945 (
            .O(N__25572),
            .I(N__25569));
    Odrv4 I__3944 (
            .O(N__25569),
            .I(\nx.n2967 ));
    InMux I__3943 (
            .O(N__25566),
            .I(\nx.n10846 ));
    CascadeMux I__3942 (
            .O(N__25563),
            .I(N__25560));
    InMux I__3941 (
            .O(N__25560),
            .I(N__25556));
    InMux I__3940 (
            .O(N__25559),
            .I(N__25553));
    LocalMux I__3939 (
            .O(N__25556),
            .I(\nx.n2899 ));
    LocalMux I__3938 (
            .O(N__25553),
            .I(\nx.n2899 ));
    InMux I__3937 (
            .O(N__25548),
            .I(N__25545));
    LocalMux I__3936 (
            .O(N__25545),
            .I(\nx.n2966 ));
    InMux I__3935 (
            .O(N__25542),
            .I(\nx.n10847 ));
    CascadeMux I__3934 (
            .O(N__25539),
            .I(N__25535));
    InMux I__3933 (
            .O(N__25538),
            .I(N__25532));
    InMux I__3932 (
            .O(N__25535),
            .I(N__25529));
    LocalMux I__3931 (
            .O(N__25532),
            .I(N__25526));
    LocalMux I__3930 (
            .O(N__25529),
            .I(N__25523));
    Odrv4 I__3929 (
            .O(N__25526),
            .I(\nx.n2898 ));
    Odrv4 I__3928 (
            .O(N__25523),
            .I(\nx.n2898 ));
    CascadeMux I__3927 (
            .O(N__25518),
            .I(N__25515));
    InMux I__3926 (
            .O(N__25515),
            .I(N__25512));
    LocalMux I__3925 (
            .O(N__25512),
            .I(\nx.n2965 ));
    InMux I__3924 (
            .O(N__25509),
            .I(\nx.n10848 ));
    CascadeMux I__3923 (
            .O(N__25506),
            .I(N__25502));
    CascadeMux I__3922 (
            .O(N__25505),
            .I(N__25499));
    InMux I__3921 (
            .O(N__25502),
            .I(N__25496));
    InMux I__3920 (
            .O(N__25499),
            .I(N__25493));
    LocalMux I__3919 (
            .O(N__25496),
            .I(N__25487));
    LocalMux I__3918 (
            .O(N__25493),
            .I(N__25487));
    InMux I__3917 (
            .O(N__25492),
            .I(N__25484));
    Odrv4 I__3916 (
            .O(N__25487),
            .I(\nx.n2897 ));
    LocalMux I__3915 (
            .O(N__25484),
            .I(\nx.n2897 ));
    InMux I__3914 (
            .O(N__25479),
            .I(N__25476));
    LocalMux I__3913 (
            .O(N__25476),
            .I(\nx.n2964 ));
    InMux I__3912 (
            .O(N__25473),
            .I(\nx.n10849 ));
    CascadeMux I__3911 (
            .O(N__25470),
            .I(N__25466));
    InMux I__3910 (
            .O(N__25469),
            .I(N__25463));
    InMux I__3909 (
            .O(N__25466),
            .I(N__25460));
    LocalMux I__3908 (
            .O(N__25463),
            .I(N__25457));
    LocalMux I__3907 (
            .O(N__25460),
            .I(\nx.n2896 ));
    Odrv4 I__3906 (
            .O(N__25457),
            .I(\nx.n2896 ));
    InMux I__3905 (
            .O(N__25452),
            .I(N__25449));
    LocalMux I__3904 (
            .O(N__25449),
            .I(N__25446));
    Odrv4 I__3903 (
            .O(N__25446),
            .I(\nx.n2963 ));
    InMux I__3902 (
            .O(N__25443),
            .I(\nx.n10850 ));
    InMux I__3901 (
            .O(N__25440),
            .I(N__25437));
    LocalMux I__3900 (
            .O(N__25437),
            .I(\nx.n2962 ));
    InMux I__3899 (
            .O(N__25434),
            .I(\nx.n10851 ));
    InMux I__3898 (
            .O(N__25431),
            .I(bfn_5_24_0_));
    InMux I__3897 (
            .O(N__25428),
            .I(N__25425));
    LocalMux I__3896 (
            .O(N__25425),
            .I(\nx.n2960 ));
    InMux I__3895 (
            .O(N__25422),
            .I(\nx.n10853 ));
    CascadeMux I__3894 (
            .O(N__25419),
            .I(N__25416));
    InMux I__3893 (
            .O(N__25416),
            .I(N__25412));
    InMux I__3892 (
            .O(N__25415),
            .I(N__25409));
    LocalMux I__3891 (
            .O(N__25412),
            .I(N__25404));
    LocalMux I__3890 (
            .O(N__25409),
            .I(N__25404));
    Span4Mux_v I__3889 (
            .O(N__25404),
            .I(N__25401));
    Odrv4 I__3888 (
            .O(N__25401),
            .I(\nx.n2908 ));
    InMux I__3887 (
            .O(N__25398),
            .I(N__25395));
    LocalMux I__3886 (
            .O(N__25395),
            .I(N__25392));
    Span4Mux_h I__3885 (
            .O(N__25392),
            .I(N__25389));
    Odrv4 I__3884 (
            .O(N__25389),
            .I(\nx.n2975 ));
    InMux I__3883 (
            .O(N__25386),
            .I(\nx.n10838 ));
    CascadeMux I__3882 (
            .O(N__25383),
            .I(N__25379));
    CascadeMux I__3881 (
            .O(N__25382),
            .I(N__25376));
    InMux I__3880 (
            .O(N__25379),
            .I(N__25373));
    InMux I__3879 (
            .O(N__25376),
            .I(N__25369));
    LocalMux I__3878 (
            .O(N__25373),
            .I(N__25366));
    InMux I__3877 (
            .O(N__25372),
            .I(N__25363));
    LocalMux I__3876 (
            .O(N__25369),
            .I(\nx.n2907 ));
    Odrv4 I__3875 (
            .O(N__25366),
            .I(\nx.n2907 ));
    LocalMux I__3874 (
            .O(N__25363),
            .I(\nx.n2907 ));
    InMux I__3873 (
            .O(N__25356),
            .I(N__25353));
    LocalMux I__3872 (
            .O(N__25353),
            .I(\nx.n2974 ));
    InMux I__3871 (
            .O(N__25350),
            .I(\nx.n10839 ));
    CascadeMux I__3870 (
            .O(N__25347),
            .I(N__25343));
    InMux I__3869 (
            .O(N__25346),
            .I(N__25339));
    InMux I__3868 (
            .O(N__25343),
            .I(N__25336));
    InMux I__3867 (
            .O(N__25342),
            .I(N__25333));
    LocalMux I__3866 (
            .O(N__25339),
            .I(\nx.n2906 ));
    LocalMux I__3865 (
            .O(N__25336),
            .I(\nx.n2906 ));
    LocalMux I__3864 (
            .O(N__25333),
            .I(\nx.n2906 ));
    InMux I__3863 (
            .O(N__25326),
            .I(N__25323));
    LocalMux I__3862 (
            .O(N__25323),
            .I(\nx.n2973 ));
    InMux I__3861 (
            .O(N__25320),
            .I(\nx.n10840 ));
    InMux I__3860 (
            .O(N__25317),
            .I(N__25314));
    LocalMux I__3859 (
            .O(N__25314),
            .I(N__25311));
    Odrv4 I__3858 (
            .O(N__25311),
            .I(\nx.n2972 ));
    InMux I__3857 (
            .O(N__25308),
            .I(\nx.n10841 ));
    InMux I__3856 (
            .O(N__25305),
            .I(\nx.n10842 ));
    CascadeMux I__3855 (
            .O(N__25302),
            .I(N__25299));
    InMux I__3854 (
            .O(N__25299),
            .I(N__25296));
    LocalMux I__3853 (
            .O(N__25296),
            .I(N__25293));
    Odrv4 I__3852 (
            .O(N__25293),
            .I(\nx.n2970 ));
    InMux I__3851 (
            .O(N__25290),
            .I(\nx.n10843 ));
    CascadeMux I__3850 (
            .O(N__25287),
            .I(N__25284));
    InMux I__3849 (
            .O(N__25284),
            .I(N__25281));
    LocalMux I__3848 (
            .O(N__25281),
            .I(N__25278));
    Span4Mux_s2_h I__3847 (
            .O(N__25278),
            .I(N__25275));
    Odrv4 I__3846 (
            .O(N__25275),
            .I(\nx.n2969 ));
    InMux I__3845 (
            .O(N__25272),
            .I(bfn_5_23_0_));
    CascadeMux I__3844 (
            .O(N__25269),
            .I(N__25265));
    InMux I__3843 (
            .O(N__25268),
            .I(N__25262));
    InMux I__3842 (
            .O(N__25265),
            .I(N__25259));
    LocalMux I__3841 (
            .O(N__25262),
            .I(N__25253));
    LocalMux I__3840 (
            .O(N__25259),
            .I(N__25253));
    InMux I__3839 (
            .O(N__25258),
            .I(N__25250));
    Odrv4 I__3838 (
            .O(N__25253),
            .I(\nx.n2901 ));
    LocalMux I__3837 (
            .O(N__25250),
            .I(\nx.n2901 ));
    InMux I__3836 (
            .O(N__25245),
            .I(N__25242));
    LocalMux I__3835 (
            .O(N__25242),
            .I(\nx.n2968 ));
    InMux I__3834 (
            .O(N__25239),
            .I(\nx.n10845 ));
    CascadeMux I__3833 (
            .O(N__25236),
            .I(\nx.n2896_cascade_ ));
    CascadeMux I__3832 (
            .O(N__25233),
            .I(\nx.n2898_cascade_ ));
    CascadeMux I__3831 (
            .O(N__25230),
            .I(\nx.n42_adj_675_cascade_ ));
    InMux I__3830 (
            .O(N__25227),
            .I(N__25224));
    LocalMux I__3829 (
            .O(N__25224),
            .I(\nx.n32_adj_674 ));
    InMux I__3828 (
            .O(N__25221),
            .I(N__25218));
    LocalMux I__3827 (
            .O(N__25218),
            .I(N__25215));
    Odrv4 I__3826 (
            .O(N__25215),
            .I(\nx.n46 ));
    InMux I__3825 (
            .O(N__25212),
            .I(N__25209));
    LocalMux I__3824 (
            .O(N__25209),
            .I(N__25206));
    Span4Mux_v I__3823 (
            .O(N__25206),
            .I(N__25203));
    Odrv4 I__3822 (
            .O(N__25203),
            .I(\nx.n2977 ));
    InMux I__3821 (
            .O(N__25200),
            .I(bfn_5_22_0_));
    CascadeMux I__3820 (
            .O(N__25197),
            .I(N__25194));
    InMux I__3819 (
            .O(N__25194),
            .I(N__25191));
    LocalMux I__3818 (
            .O(N__25191),
            .I(N__25188));
    Span4Mux_h I__3817 (
            .O(N__25188),
            .I(N__25185));
    Odrv4 I__3816 (
            .O(N__25185),
            .I(\nx.n2976 ));
    InMux I__3815 (
            .O(N__25182),
            .I(\nx.n10837 ));
    CascadeMux I__3814 (
            .O(N__25179),
            .I(N__25176));
    InMux I__3813 (
            .O(N__25176),
            .I(N__25172));
    InMux I__3812 (
            .O(N__25175),
            .I(N__25169));
    LocalMux I__3811 (
            .O(N__25172),
            .I(N__25165));
    LocalMux I__3810 (
            .O(N__25169),
            .I(N__25162));
    InMux I__3809 (
            .O(N__25168),
            .I(N__25159));
    Span4Mux_v I__3808 (
            .O(N__25165),
            .I(N__25156));
    Odrv4 I__3807 (
            .O(N__25162),
            .I(timer_20));
    LocalMux I__3806 (
            .O(N__25159),
            .I(timer_20));
    Odrv4 I__3805 (
            .O(N__25156),
            .I(timer_20));
    InMux I__3804 (
            .O(N__25149),
            .I(N__25143));
    InMux I__3803 (
            .O(N__25148),
            .I(N__25143));
    LocalMux I__3802 (
            .O(N__25143),
            .I(neo_pixel_transmitter_t0_20));
    CascadeMux I__3801 (
            .O(N__25140),
            .I(\nx.n2809_cascade_ ));
    CascadeMux I__3800 (
            .O(N__25137),
            .I(\nx.n31_adj_613_cascade_ ));
    InMux I__3799 (
            .O(N__25134),
            .I(N__25131));
    LocalMux I__3798 (
            .O(N__25131),
            .I(\nx.n39_adj_614 ));
    InMux I__3797 (
            .O(N__25128),
            .I(N__25125));
    LocalMux I__3796 (
            .O(N__25125),
            .I(N__25121));
    InMux I__3795 (
            .O(N__25124),
            .I(N__25117));
    Span4Mux_v I__3794 (
            .O(N__25121),
            .I(N__25114));
    InMux I__3793 (
            .O(N__25120),
            .I(N__25111));
    LocalMux I__3792 (
            .O(N__25117),
            .I(N__25108));
    Odrv4 I__3791 (
            .O(N__25114),
            .I(timer_19));
    LocalMux I__3790 (
            .O(N__25111),
            .I(timer_19));
    Odrv12 I__3789 (
            .O(N__25108),
            .I(timer_19));
    InMux I__3788 (
            .O(N__25101),
            .I(N__25098));
    LocalMux I__3787 (
            .O(N__25098),
            .I(N__25095));
    Odrv4 I__3786 (
            .O(N__25095),
            .I(n13171));
    InMux I__3785 (
            .O(N__25092),
            .I(N__25089));
    LocalMux I__3784 (
            .O(N__25089),
            .I(n13170));
    InMux I__3783 (
            .O(N__25086),
            .I(N__25082));
    InMux I__3782 (
            .O(N__25085),
            .I(N__25079));
    LocalMux I__3781 (
            .O(N__25082),
            .I(neo_pixel_transmitter_t0_9));
    LocalMux I__3780 (
            .O(N__25079),
            .I(neo_pixel_transmitter_t0_9));
    InMux I__3779 (
            .O(N__25074),
            .I(N__25071));
    LocalMux I__3778 (
            .O(N__25071),
            .I(N__25068));
    Span4Mux_v I__3777 (
            .O(N__25068),
            .I(N__25065));
    Span4Mux_s2_h I__3776 (
            .O(N__25065),
            .I(N__25062));
    Odrv4 I__3775 (
            .O(N__25062),
            .I(\nx.n24 ));
    InMux I__3774 (
            .O(N__25059),
            .I(N__25055));
    InMux I__3773 (
            .O(N__25058),
            .I(N__25052));
    LocalMux I__3772 (
            .O(N__25055),
            .I(neo_pixel_transmitter_t0_19));
    LocalMux I__3771 (
            .O(N__25052),
            .I(neo_pixel_transmitter_t0_19));
    CascadeMux I__3770 (
            .O(N__25047),
            .I(N__25044));
    InMux I__3769 (
            .O(N__25044),
            .I(N__25041));
    LocalMux I__3768 (
            .O(N__25041),
            .I(N__25038));
    Span4Mux_h I__3767 (
            .O(N__25038),
            .I(N__25035));
    Span4Mux_v I__3766 (
            .O(N__25035),
            .I(N__25032));
    Odrv4 I__3765 (
            .O(N__25032),
            .I(\nx.n14 ));
    InMux I__3764 (
            .O(N__25029),
            .I(N__25026));
    LocalMux I__3763 (
            .O(N__25026),
            .I(neopxl_color_prev_6));
    InMux I__3762 (
            .O(N__25023),
            .I(N__25020));
    LocalMux I__3761 (
            .O(N__25020),
            .I(N__25017));
    Odrv4 I__3760 (
            .O(N__25017),
            .I(neopxl_color_prev_15));
    InMux I__3759 (
            .O(N__25014),
            .I(N__25011));
    LocalMux I__3758 (
            .O(N__25011),
            .I(N__25008));
    Odrv12 I__3757 (
            .O(N__25008),
            .I(n11_adj_775));
    CascadeMux I__3756 (
            .O(N__25005),
            .I(N__25002));
    InMux I__3755 (
            .O(N__25002),
            .I(N__24999));
    LocalMux I__3754 (
            .O(N__24999),
            .I(N__24996));
    Span4Mux_v I__3753 (
            .O(N__24996),
            .I(N__24993));
    Odrv4 I__3752 (
            .O(N__24993),
            .I(neopxl_color_prev_13));
    InMux I__3751 (
            .O(N__24990),
            .I(N__24987));
    LocalMux I__3750 (
            .O(N__24987),
            .I(N__24984));
    Span4Mux_h I__3749 (
            .O(N__24984),
            .I(N__24981));
    Span4Mux_v I__3748 (
            .O(N__24981),
            .I(N__24978));
    Odrv4 I__3747 (
            .O(N__24978),
            .I(\nx.n13_adj_649 ));
    InMux I__3746 (
            .O(N__24975),
            .I(N__24972));
    LocalMux I__3745 (
            .O(N__24972),
            .I(N__24965));
    InMux I__3744 (
            .O(N__24971),
            .I(N__24962));
    InMux I__3743 (
            .O(N__24970),
            .I(N__24959));
    InMux I__3742 (
            .O(N__24969),
            .I(N__24956));
    InMux I__3741 (
            .O(N__24968),
            .I(N__24953));
    Span4Mux_s1_v I__3740 (
            .O(N__24965),
            .I(N__24946));
    LocalMux I__3739 (
            .O(N__24962),
            .I(N__24946));
    LocalMux I__3738 (
            .O(N__24959),
            .I(N__24946));
    LocalMux I__3737 (
            .O(N__24956),
            .I(\nx.bit_ctr_21 ));
    LocalMux I__3736 (
            .O(N__24953),
            .I(\nx.bit_ctr_21 ));
    Odrv4 I__3735 (
            .O(N__24946),
            .I(\nx.bit_ctr_21 ));
    InMux I__3734 (
            .O(N__24939),
            .I(N__24936));
    LocalMux I__3733 (
            .O(N__24936),
            .I(\nx.n1477 ));
    CascadeMux I__3732 (
            .O(N__24933),
            .I(\nx.n1509_cascade_ ));
    InMux I__3731 (
            .O(N__24930),
            .I(N__24927));
    LocalMux I__3730 (
            .O(N__24927),
            .I(\nx.n16_adj_629 ));
    CascadeMux I__3729 (
            .O(N__24924),
            .I(\nx.n18_adj_630_cascade_ ));
    InMux I__3728 (
            .O(N__24921),
            .I(N__24918));
    LocalMux I__3727 (
            .O(N__24918),
            .I(\nx.n13_adj_631 ));
    InMux I__3726 (
            .O(N__24915),
            .I(N__24912));
    LocalMux I__3725 (
            .O(N__24912),
            .I(N__24909));
    Odrv4 I__3724 (
            .O(N__24909),
            .I(\nx.n1469 ));
    CascadeMux I__3723 (
            .O(N__24906),
            .I(\nx.n1433_cascade_ ));
    CascadeMux I__3722 (
            .O(N__24903),
            .I(N__24899));
    InMux I__3721 (
            .O(N__24902),
            .I(N__24895));
    InMux I__3720 (
            .O(N__24899),
            .I(N__24890));
    InMux I__3719 (
            .O(N__24898),
            .I(N__24890));
    LocalMux I__3718 (
            .O(N__24895),
            .I(\nx.n1402 ));
    LocalMux I__3717 (
            .O(N__24890),
            .I(\nx.n1402 ));
    CascadeMux I__3716 (
            .O(N__24885),
            .I(\nx.n1501_cascade_ ));
    InMux I__3715 (
            .O(N__24882),
            .I(N__24879));
    LocalMux I__3714 (
            .O(N__24879),
            .I(\nx.n9672 ));
    InMux I__3713 (
            .O(N__24876),
            .I(N__24873));
    LocalMux I__3712 (
            .O(N__24873),
            .I(N__24869));
    InMux I__3711 (
            .O(N__24872),
            .I(N__24865));
    Span4Mux_h I__3710 (
            .O(N__24869),
            .I(N__24862));
    InMux I__3709 (
            .O(N__24868),
            .I(N__24859));
    LocalMux I__3708 (
            .O(N__24865),
            .I(N__24856));
    Odrv4 I__3707 (
            .O(N__24862),
            .I(timer_22));
    LocalMux I__3706 (
            .O(N__24859),
            .I(timer_22));
    Odrv12 I__3705 (
            .O(N__24856),
            .I(timer_22));
    InMux I__3704 (
            .O(N__24849),
            .I(\nx.n10421 ));
    CEMux I__3703 (
            .O(N__24846),
            .I(N__24841));
    CEMux I__3702 (
            .O(N__24845),
            .I(N__24837));
    CEMux I__3701 (
            .O(N__24844),
            .I(N__24834));
    LocalMux I__3700 (
            .O(N__24841),
            .I(N__24831));
    CEMux I__3699 (
            .O(N__24840),
            .I(N__24828));
    LocalMux I__3698 (
            .O(N__24837),
            .I(N__24825));
    LocalMux I__3697 (
            .O(N__24834),
            .I(N__24822));
    Span4Mux_h I__3696 (
            .O(N__24831),
            .I(N__24817));
    LocalMux I__3695 (
            .O(N__24828),
            .I(N__24817));
    Span4Mux_v I__3694 (
            .O(N__24825),
            .I(N__24814));
    Span4Mux_h I__3693 (
            .O(N__24822),
            .I(N__24811));
    Span4Mux_v I__3692 (
            .O(N__24817),
            .I(N__24808));
    Span4Mux_v I__3691 (
            .O(N__24814),
            .I(N__24805));
    Span4Mux_v I__3690 (
            .O(N__24811),
            .I(N__24802));
    Span4Mux_h I__3689 (
            .O(N__24808),
            .I(N__24799));
    Span4Mux_v I__3688 (
            .O(N__24805),
            .I(N__24796));
    Span4Mux_v I__3687 (
            .O(N__24802),
            .I(N__24793));
    Span4Mux_v I__3686 (
            .O(N__24799),
            .I(N__24790));
    Odrv4 I__3685 (
            .O(N__24796),
            .I(\nx.n7230 ));
    Odrv4 I__3684 (
            .O(N__24793),
            .I(\nx.n7230 ));
    Odrv4 I__3683 (
            .O(N__24790),
            .I(\nx.n7230 ));
    SRMux I__3682 (
            .O(N__24783),
            .I(N__24780));
    LocalMux I__3681 (
            .O(N__24780),
            .I(N__24775));
    SRMux I__3680 (
            .O(N__24779),
            .I(N__24772));
    SRMux I__3679 (
            .O(N__24778),
            .I(N__24769));
    Span4Mux_v I__3678 (
            .O(N__24775),
            .I(N__24765));
    LocalMux I__3677 (
            .O(N__24772),
            .I(N__24760));
    LocalMux I__3676 (
            .O(N__24769),
            .I(N__24760));
    SRMux I__3675 (
            .O(N__24768),
            .I(N__24757));
    Span4Mux_h I__3674 (
            .O(N__24765),
            .I(N__24750));
    Span4Mux_v I__3673 (
            .O(N__24760),
            .I(N__24750));
    LocalMux I__3672 (
            .O(N__24757),
            .I(N__24750));
    Span4Mux_h I__3671 (
            .O(N__24750),
            .I(N__24747));
    Span4Mux_v I__3670 (
            .O(N__24747),
            .I(N__24744));
    Span4Mux_v I__3669 (
            .O(N__24744),
            .I(N__24741));
    Odrv4 I__3668 (
            .O(N__24741),
            .I(\nx.n7411 ));
    InMux I__3667 (
            .O(N__24738),
            .I(N__24735));
    LocalMux I__3666 (
            .O(N__24735),
            .I(N__24730));
    CascadeMux I__3665 (
            .O(N__24734),
            .I(N__24727));
    InMux I__3664 (
            .O(N__24733),
            .I(N__24724));
    Span4Mux_h I__3663 (
            .O(N__24730),
            .I(N__24721));
    InMux I__3662 (
            .O(N__24727),
            .I(N__24718));
    LocalMux I__3661 (
            .O(N__24724),
            .I(N__24715));
    Odrv4 I__3660 (
            .O(N__24721),
            .I(\nx.n1308 ));
    LocalMux I__3659 (
            .O(N__24718),
            .I(\nx.n1308 ));
    Odrv4 I__3658 (
            .O(N__24715),
            .I(\nx.n1308 ));
    CascadeMux I__3657 (
            .O(N__24708),
            .I(N__24705));
    InMux I__3656 (
            .O(N__24705),
            .I(N__24702));
    LocalMux I__3655 (
            .O(N__24702),
            .I(N__24699));
    Odrv4 I__3654 (
            .O(N__24699),
            .I(\nx.n1375 ));
    InMux I__3653 (
            .O(N__24696),
            .I(N__24693));
    LocalMux I__3652 (
            .O(N__24693),
            .I(N__24690));
    Odrv4 I__3651 (
            .O(N__24690),
            .I(\nx.n1373 ));
    InMux I__3650 (
            .O(N__24687),
            .I(N__24684));
    LocalMux I__3649 (
            .O(N__24684),
            .I(N__24680));
    CascadeMux I__3648 (
            .O(N__24683),
            .I(N__24677));
    Span4Mux_s2_v I__3647 (
            .O(N__24680),
            .I(N__24674));
    InMux I__3646 (
            .O(N__24677),
            .I(N__24671));
    Odrv4 I__3645 (
            .O(N__24674),
            .I(\nx.n1306 ));
    LocalMux I__3644 (
            .O(N__24671),
            .I(\nx.n1306 ));
    InMux I__3643 (
            .O(N__24666),
            .I(N__24663));
    LocalMux I__3642 (
            .O(N__24663),
            .I(N__24660));
    Odrv4 I__3641 (
            .O(N__24660),
            .I(\nx.n1371 ));
    CascadeMux I__3640 (
            .O(N__24657),
            .I(N__24654));
    InMux I__3639 (
            .O(N__24654),
            .I(N__24649));
    InMux I__3638 (
            .O(N__24653),
            .I(N__24646));
    InMux I__3637 (
            .O(N__24652),
            .I(N__24643));
    LocalMux I__3636 (
            .O(N__24649),
            .I(\nx.n1304 ));
    LocalMux I__3635 (
            .O(N__24646),
            .I(\nx.n1304 ));
    LocalMux I__3634 (
            .O(N__24643),
            .I(\nx.n1304 ));
    InMux I__3633 (
            .O(N__24636),
            .I(N__24632));
    InMux I__3632 (
            .O(N__24635),
            .I(N__24628));
    LocalMux I__3631 (
            .O(N__24632),
            .I(N__24625));
    CascadeMux I__3630 (
            .O(N__24631),
            .I(N__24622));
    LocalMux I__3629 (
            .O(N__24628),
            .I(N__24619));
    Span4Mux_h I__3628 (
            .O(N__24625),
            .I(N__24616));
    InMux I__3627 (
            .O(N__24622),
            .I(N__24613));
    Span4Mux_h I__3626 (
            .O(N__24619),
            .I(N__24610));
    Odrv4 I__3625 (
            .O(N__24616),
            .I(\nx.n1305 ));
    LocalMux I__3624 (
            .O(N__24613),
            .I(\nx.n1305 ));
    Odrv4 I__3623 (
            .O(N__24610),
            .I(\nx.n1305 ));
    CascadeMux I__3622 (
            .O(N__24603),
            .I(N__24600));
    InMux I__3621 (
            .O(N__24600),
            .I(N__24597));
    LocalMux I__3620 (
            .O(N__24597),
            .I(N__24594));
    Odrv4 I__3619 (
            .O(N__24594),
            .I(\nx.n1372 ));
    CascadeMux I__3618 (
            .O(N__24591),
            .I(N__24582));
    InMux I__3617 (
            .O(N__24590),
            .I(N__24577));
    InMux I__3616 (
            .O(N__24589),
            .I(N__24572));
    InMux I__3615 (
            .O(N__24588),
            .I(N__24572));
    InMux I__3614 (
            .O(N__24587),
            .I(N__24567));
    InMux I__3613 (
            .O(N__24586),
            .I(N__24567));
    InMux I__3612 (
            .O(N__24585),
            .I(N__24558));
    InMux I__3611 (
            .O(N__24582),
            .I(N__24558));
    InMux I__3610 (
            .O(N__24581),
            .I(N__24558));
    InMux I__3609 (
            .O(N__24580),
            .I(N__24558));
    LocalMux I__3608 (
            .O(N__24577),
            .I(N__24553));
    LocalMux I__3607 (
            .O(N__24572),
            .I(N__24553));
    LocalMux I__3606 (
            .O(N__24567),
            .I(\nx.n1334 ));
    LocalMux I__3605 (
            .O(N__24558),
            .I(\nx.n1334 ));
    Odrv4 I__3604 (
            .O(N__24553),
            .I(\nx.n1334 ));
    CascadeMux I__3603 (
            .O(N__24546),
            .I(\nx.n1404_cascade_ ));
    InMux I__3602 (
            .O(N__24543),
            .I(N__24538));
    InMux I__3601 (
            .O(N__24542),
            .I(N__24535));
    InMux I__3600 (
            .O(N__24541),
            .I(N__24530));
    LocalMux I__3599 (
            .O(N__24538),
            .I(N__24527));
    LocalMux I__3598 (
            .O(N__24535),
            .I(N__24524));
    InMux I__3597 (
            .O(N__24534),
            .I(N__24521));
    InMux I__3596 (
            .O(N__24533),
            .I(N__24518));
    LocalMux I__3595 (
            .O(N__24530),
            .I(N__24513));
    Span4Mux_s3_h I__3594 (
            .O(N__24527),
            .I(N__24513));
    Span4Mux_s3_h I__3593 (
            .O(N__24524),
            .I(N__24510));
    LocalMux I__3592 (
            .O(N__24521),
            .I(\nx.bit_ctr_23 ));
    LocalMux I__3591 (
            .O(N__24518),
            .I(\nx.bit_ctr_23 ));
    Odrv4 I__3590 (
            .O(N__24513),
            .I(\nx.bit_ctr_23 ));
    Odrv4 I__3589 (
            .O(N__24510),
            .I(\nx.bit_ctr_23 ));
    InMux I__3588 (
            .O(N__24501),
            .I(N__24498));
    LocalMux I__3587 (
            .O(N__24498),
            .I(N__24495));
    Span4Mux_h I__3586 (
            .O(N__24495),
            .I(N__24492));
    Odrv4 I__3585 (
            .O(N__24492),
            .I(\nx.n47_adj_706 ));
    CascadeMux I__3584 (
            .O(N__24489),
            .I(N__24485));
    InMux I__3583 (
            .O(N__24488),
            .I(N__24482));
    InMux I__3582 (
            .O(N__24485),
            .I(N__24479));
    LocalMux I__3581 (
            .O(N__24482),
            .I(\nx.n1404 ));
    LocalMux I__3580 (
            .O(N__24479),
            .I(\nx.n1404 ));
    InMux I__3579 (
            .O(N__24474),
            .I(N__24471));
    LocalMux I__3578 (
            .O(N__24471),
            .I(\nx.n1471 ));
    InMux I__3577 (
            .O(N__24468),
            .I(\nx.n10412 ));
    InMux I__3576 (
            .O(N__24465),
            .I(\nx.n10413 ));
    CascadeMux I__3575 (
            .O(N__24462),
            .I(N__24457));
    InMux I__3574 (
            .O(N__24461),
            .I(N__24451));
    InMux I__3573 (
            .O(N__24460),
            .I(N__24451));
    InMux I__3572 (
            .O(N__24457),
            .I(N__24448));
    InMux I__3571 (
            .O(N__24456),
            .I(N__24445));
    LocalMux I__3570 (
            .O(N__24451),
            .I(N__24441));
    LocalMux I__3569 (
            .O(N__24448),
            .I(N__24436));
    LocalMux I__3568 (
            .O(N__24445),
            .I(N__24436));
    InMux I__3567 (
            .O(N__24444),
            .I(N__24433));
    Span4Mux_s1_h I__3566 (
            .O(N__24441),
            .I(N__24428));
    Span4Mux_v I__3565 (
            .O(N__24436),
            .I(N__24428));
    LocalMux I__3564 (
            .O(N__24433),
            .I(\nx.bit_ctr_24 ));
    Odrv4 I__3563 (
            .O(N__24428),
            .I(\nx.bit_ctr_24 ));
    InMux I__3562 (
            .O(N__24423),
            .I(bfn_4_30_0_));
    InMux I__3561 (
            .O(N__24420),
            .I(\nx.n10415 ));
    InMux I__3560 (
            .O(N__24417),
            .I(\nx.n10416 ));
    InMux I__3559 (
            .O(N__24414),
            .I(\nx.n10417 ));
    InMux I__3558 (
            .O(N__24411),
            .I(\nx.n10418 ));
    InMux I__3557 (
            .O(N__24408),
            .I(\nx.n10419 ));
    InMux I__3556 (
            .O(N__24405),
            .I(\nx.n10420 ));
    InMux I__3555 (
            .O(N__24402),
            .I(\nx.n10403 ));
    InMux I__3554 (
            .O(N__24399),
            .I(\nx.n10404 ));
    InMux I__3553 (
            .O(N__24396),
            .I(\nx.n10405 ));
    InMux I__3552 (
            .O(N__24393),
            .I(bfn_4_29_0_));
    InMux I__3551 (
            .O(N__24390),
            .I(\nx.n10407 ));
    InMux I__3550 (
            .O(N__24387),
            .I(\nx.n10408 ));
    InMux I__3549 (
            .O(N__24384),
            .I(\nx.n10409 ));
    InMux I__3548 (
            .O(N__24381),
            .I(\nx.n10410 ));
    InMux I__3547 (
            .O(N__24378),
            .I(\nx.n10411 ));
    InMux I__3546 (
            .O(N__24375),
            .I(N__24371));
    InMux I__3545 (
            .O(N__24374),
            .I(N__24366));
    LocalMux I__3544 (
            .O(N__24371),
            .I(N__24363));
    InMux I__3543 (
            .O(N__24370),
            .I(N__24360));
    InMux I__3542 (
            .O(N__24369),
            .I(N__24357));
    LocalMux I__3541 (
            .O(N__24366),
            .I(N__24353));
    Span4Mux_v I__3540 (
            .O(N__24363),
            .I(N__24350));
    LocalMux I__3539 (
            .O(N__24360),
            .I(N__24345));
    LocalMux I__3538 (
            .O(N__24357),
            .I(N__24345));
    InMux I__3537 (
            .O(N__24356),
            .I(N__24342));
    Span4Mux_v I__3536 (
            .O(N__24353),
            .I(N__24335));
    Span4Mux_s1_h I__3535 (
            .O(N__24350),
            .I(N__24335));
    Span4Mux_v I__3534 (
            .O(N__24345),
            .I(N__24335));
    LocalMux I__3533 (
            .O(N__24342),
            .I(\nx.bit_ctr_4 ));
    Odrv4 I__3532 (
            .O(N__24335),
            .I(\nx.bit_ctr_4 ));
    InMux I__3531 (
            .O(N__24330),
            .I(\nx.n10394 ));
    InMux I__3530 (
            .O(N__24327),
            .I(\nx.n10395 ));
    InMux I__3529 (
            .O(N__24324),
            .I(\nx.n10396 ));
    InMux I__3528 (
            .O(N__24321),
            .I(\nx.n10397 ));
    InMux I__3527 (
            .O(N__24318),
            .I(bfn_4_28_0_));
    InMux I__3526 (
            .O(N__24315),
            .I(\nx.n10399 ));
    InMux I__3525 (
            .O(N__24312),
            .I(\nx.n10400 ));
    InMux I__3524 (
            .O(N__24309),
            .I(\nx.n10401 ));
    InMux I__3523 (
            .O(N__24306),
            .I(\nx.n10402 ));
    InMux I__3522 (
            .O(N__24303),
            .I(N__24300));
    LocalMux I__3521 (
            .O(N__24300),
            .I(N__24297));
    Span4Mux_h I__3520 (
            .O(N__24297),
            .I(N__24294));
    Odrv4 I__3519 (
            .O(N__24294),
            .I(\nx.n3157 ));
    CascadeMux I__3518 (
            .O(N__24291),
            .I(\nx.n12361_cascade_ ));
    CascadeMux I__3517 (
            .O(N__24288),
            .I(N__24285));
    InMux I__3516 (
            .O(N__24285),
            .I(N__24282));
    LocalMux I__3515 (
            .O(N__24282),
            .I(N__24278));
    InMux I__3514 (
            .O(N__24281),
            .I(N__24274));
    Span4Mux_v I__3513 (
            .O(N__24278),
            .I(N__24271));
    InMux I__3512 (
            .O(N__24277),
            .I(N__24268));
    LocalMux I__3511 (
            .O(N__24274),
            .I(\nx.n3090 ));
    Odrv4 I__3510 (
            .O(N__24271),
            .I(\nx.n3090 ));
    LocalMux I__3509 (
            .O(N__24268),
            .I(\nx.n3090 ));
    InMux I__3508 (
            .O(N__24261),
            .I(N__24258));
    LocalMux I__3507 (
            .O(N__24258),
            .I(N__24255));
    Span4Mux_h I__3506 (
            .O(N__24255),
            .I(N__24252));
    Odrv4 I__3505 (
            .O(N__24252),
            .I(\nx.n3156 ));
    CascadeMux I__3504 (
            .O(N__24249),
            .I(\nx.n12363_cascade_ ));
    CascadeMux I__3503 (
            .O(N__24246),
            .I(N__24243));
    InMux I__3502 (
            .O(N__24243),
            .I(N__24231));
    InMux I__3501 (
            .O(N__24242),
            .I(N__24218));
    InMux I__3500 (
            .O(N__24241),
            .I(N__24218));
    InMux I__3499 (
            .O(N__24240),
            .I(N__24218));
    InMux I__3498 (
            .O(N__24239),
            .I(N__24218));
    InMux I__3497 (
            .O(N__24238),
            .I(N__24218));
    InMux I__3496 (
            .O(N__24237),
            .I(N__24218));
    CascadeMux I__3495 (
            .O(N__24236),
            .I(N__24215));
    CascadeMux I__3494 (
            .O(N__24235),
            .I(N__24210));
    InMux I__3493 (
            .O(N__24234),
            .I(N__24204));
    LocalMux I__3492 (
            .O(N__24231),
            .I(N__24201));
    LocalMux I__3491 (
            .O(N__24218),
            .I(N__24198));
    InMux I__3490 (
            .O(N__24215),
            .I(N__24195));
    InMux I__3489 (
            .O(N__24214),
            .I(N__24190));
    InMux I__3488 (
            .O(N__24213),
            .I(N__24190));
    InMux I__3487 (
            .O(N__24210),
            .I(N__24185));
    InMux I__3486 (
            .O(N__24209),
            .I(N__24185));
    CascadeMux I__3485 (
            .O(N__24208),
            .I(N__24182));
    CascadeMux I__3484 (
            .O(N__24207),
            .I(N__24178));
    LocalMux I__3483 (
            .O(N__24204),
            .I(N__24164));
    Span4Mux_v I__3482 (
            .O(N__24201),
            .I(N__24157));
    Span4Mux_v I__3481 (
            .O(N__24198),
            .I(N__24157));
    LocalMux I__3480 (
            .O(N__24195),
            .I(N__24157));
    LocalMux I__3479 (
            .O(N__24190),
            .I(N__24152));
    LocalMux I__3478 (
            .O(N__24185),
            .I(N__24152));
    InMux I__3477 (
            .O(N__24182),
            .I(N__24137));
    InMux I__3476 (
            .O(N__24181),
            .I(N__24137));
    InMux I__3475 (
            .O(N__24178),
            .I(N__24137));
    InMux I__3474 (
            .O(N__24177),
            .I(N__24137));
    InMux I__3473 (
            .O(N__24176),
            .I(N__24137));
    InMux I__3472 (
            .O(N__24175),
            .I(N__24137));
    InMux I__3471 (
            .O(N__24174),
            .I(N__24137));
    InMux I__3470 (
            .O(N__24173),
            .I(N__24132));
    InMux I__3469 (
            .O(N__24172),
            .I(N__24132));
    InMux I__3468 (
            .O(N__24171),
            .I(N__24127));
    InMux I__3467 (
            .O(N__24170),
            .I(N__24127));
    InMux I__3466 (
            .O(N__24169),
            .I(N__24120));
    InMux I__3465 (
            .O(N__24168),
            .I(N__24120));
    InMux I__3464 (
            .O(N__24167),
            .I(N__24120));
    Odrv4 I__3463 (
            .O(N__24164),
            .I(\nx.n3116 ));
    Odrv4 I__3462 (
            .O(N__24157),
            .I(\nx.n3116 ));
    Odrv4 I__3461 (
            .O(N__24152),
            .I(\nx.n3116 ));
    LocalMux I__3460 (
            .O(N__24137),
            .I(\nx.n3116 ));
    LocalMux I__3459 (
            .O(N__24132),
            .I(\nx.n3116 ));
    LocalMux I__3458 (
            .O(N__24127),
            .I(\nx.n3116 ));
    LocalMux I__3457 (
            .O(N__24120),
            .I(\nx.n3116 ));
    InMux I__3456 (
            .O(N__24105),
            .I(N__24102));
    LocalMux I__3455 (
            .O(N__24102),
            .I(N__24098));
    InMux I__3454 (
            .O(N__24101),
            .I(N__24095));
    Span4Mux_v I__3453 (
            .O(N__24098),
            .I(N__24092));
    LocalMux I__3452 (
            .O(N__24095),
            .I(\nx.n3088 ));
    Odrv4 I__3451 (
            .O(N__24092),
            .I(\nx.n3088 ));
    CascadeMux I__3450 (
            .O(N__24087),
            .I(\nx.n12365_cascade_ ));
    InMux I__3449 (
            .O(N__24084),
            .I(N__24081));
    LocalMux I__3448 (
            .O(N__24081),
            .I(N__24078));
    Span4Mux_h I__3447 (
            .O(N__24078),
            .I(N__24075));
    Odrv4 I__3446 (
            .O(N__24075),
            .I(\nx.n3155 ));
    InMux I__3445 (
            .O(N__24072),
            .I(N__24069));
    LocalMux I__3444 (
            .O(N__24069),
            .I(N__24066));
    Span4Mux_s1_h I__3443 (
            .O(N__24066),
            .I(N__24063));
    Span4Mux_v I__3442 (
            .O(N__24063),
            .I(N__24060));
    Odrv4 I__3441 (
            .O(N__24060),
            .I(\nx.n12367 ));
    CascadeMux I__3440 (
            .O(N__24057),
            .I(N__24054));
    InMux I__3439 (
            .O(N__24054),
            .I(N__24050));
    InMux I__3438 (
            .O(N__24053),
            .I(N__24047));
    LocalMux I__3437 (
            .O(N__24050),
            .I(N__24044));
    LocalMux I__3436 (
            .O(N__24047),
            .I(N__24040));
    Span4Mux_v I__3435 (
            .O(N__24044),
            .I(N__24037));
    InMux I__3434 (
            .O(N__24043),
            .I(N__24034));
    Odrv4 I__3433 (
            .O(N__24040),
            .I(\nx.n2990 ));
    Odrv4 I__3432 (
            .O(N__24037),
            .I(\nx.n2990 ));
    LocalMux I__3431 (
            .O(N__24034),
            .I(\nx.n2990 ));
    CascadeMux I__3430 (
            .O(N__24027),
            .I(N__24024));
    InMux I__3429 (
            .O(N__24024),
            .I(N__24021));
    LocalMux I__3428 (
            .O(N__24021),
            .I(N__24018));
    Odrv4 I__3427 (
            .O(N__24018),
            .I(\nx.n3057 ));
    InMux I__3426 (
            .O(N__24015),
            .I(N__24011));
    InMux I__3425 (
            .O(N__24014),
            .I(N__24008));
    LocalMux I__3424 (
            .O(N__24011),
            .I(N__24005));
    LocalMux I__3423 (
            .O(N__24008),
            .I(N__23999));
    Span4Mux_s3_h I__3422 (
            .O(N__24005),
            .I(N__23999));
    InMux I__3421 (
            .O(N__24004),
            .I(N__23996));
    Odrv4 I__3420 (
            .O(N__23999),
            .I(\nx.n3089 ));
    LocalMux I__3419 (
            .O(N__23996),
            .I(\nx.n3089 ));
    InMux I__3418 (
            .O(N__23991),
            .I(N__23986));
    InMux I__3417 (
            .O(N__23990),
            .I(N__23983));
    InMux I__3416 (
            .O(N__23989),
            .I(N__23980));
    LocalMux I__3415 (
            .O(N__23986),
            .I(N__23976));
    LocalMux I__3414 (
            .O(N__23983),
            .I(N__23971));
    LocalMux I__3413 (
            .O(N__23980),
            .I(N__23971));
    InMux I__3412 (
            .O(N__23979),
            .I(N__23968));
    Span4Mux_v I__3411 (
            .O(N__23976),
            .I(N__23963));
    Span4Mux_v I__3410 (
            .O(N__23971),
            .I(N__23963));
    LocalMux I__3409 (
            .O(N__23968),
            .I(N__23960));
    Span4Mux_v I__3408 (
            .O(N__23963),
            .I(N__23956));
    Span12Mux_v I__3407 (
            .O(N__23960),
            .I(N__23953));
    InMux I__3406 (
            .O(N__23959),
            .I(N__23950));
    Odrv4 I__3405 (
            .O(N__23956),
            .I(\nx.bit_ctr_0 ));
    Odrv12 I__3404 (
            .O(N__23953),
            .I(\nx.bit_ctr_0 ));
    LocalMux I__3403 (
            .O(N__23950),
            .I(\nx.bit_ctr_0 ));
    InMux I__3402 (
            .O(N__23943),
            .I(bfn_4_27_0_));
    CascadeMux I__3401 (
            .O(N__23940),
            .I(N__23937));
    InMux I__3400 (
            .O(N__23937),
            .I(N__23934));
    LocalMux I__3399 (
            .O(N__23934),
            .I(N__23931));
    Span4Mux_s3_h I__3398 (
            .O(N__23931),
            .I(N__23928));
    Span4Mux_v I__3397 (
            .O(N__23928),
            .I(N__23924));
    InMux I__3396 (
            .O(N__23927),
            .I(N__23921));
    Odrv4 I__3395 (
            .O(N__23924),
            .I(\nx.bit_ctr_1 ));
    LocalMux I__3394 (
            .O(N__23921),
            .I(\nx.bit_ctr_1 ));
    InMux I__3393 (
            .O(N__23916),
            .I(\nx.n10391 ));
    InMux I__3392 (
            .O(N__23913),
            .I(N__23910));
    LocalMux I__3391 (
            .O(N__23910),
            .I(N__23907));
    Span4Mux_v I__3390 (
            .O(N__23907),
            .I(N__23904));
    Span4Mux_v I__3389 (
            .O(N__23904),
            .I(N__23900));
    InMux I__3388 (
            .O(N__23903),
            .I(N__23897));
    Odrv4 I__3387 (
            .O(N__23900),
            .I(\nx.bit_ctr_2 ));
    LocalMux I__3386 (
            .O(N__23897),
            .I(\nx.bit_ctr_2 ));
    InMux I__3385 (
            .O(N__23892),
            .I(\nx.n10392 ));
    InMux I__3384 (
            .O(N__23889),
            .I(N__23882));
    InMux I__3383 (
            .O(N__23888),
            .I(N__23882));
    InMux I__3382 (
            .O(N__23887),
            .I(N__23879));
    LocalMux I__3381 (
            .O(N__23882),
            .I(N__23874));
    LocalMux I__3380 (
            .O(N__23879),
            .I(N__23871));
    InMux I__3379 (
            .O(N__23878),
            .I(N__23868));
    InMux I__3378 (
            .O(N__23877),
            .I(N__23865));
    Span4Mux_v I__3377 (
            .O(N__23874),
            .I(N__23858));
    Span4Mux_v I__3376 (
            .O(N__23871),
            .I(N__23858));
    LocalMux I__3375 (
            .O(N__23868),
            .I(N__23858));
    LocalMux I__3374 (
            .O(N__23865),
            .I(N__23853));
    Span4Mux_v I__3373 (
            .O(N__23858),
            .I(N__23853));
    Odrv4 I__3372 (
            .O(N__23853),
            .I(\nx.bit_ctr_3 ));
    InMux I__3371 (
            .O(N__23850),
            .I(\nx.n10393 ));
    CascadeMux I__3370 (
            .O(N__23847),
            .I(N__23843));
    CascadeMux I__3369 (
            .O(N__23846),
            .I(N__23840));
    InMux I__3368 (
            .O(N__23843),
            .I(N__23837));
    InMux I__3367 (
            .O(N__23840),
            .I(N__23834));
    LocalMux I__3366 (
            .O(N__23837),
            .I(N__23829));
    LocalMux I__3365 (
            .O(N__23834),
            .I(N__23829));
    Span4Mux_v I__3364 (
            .O(N__23829),
            .I(N__23825));
    InMux I__3363 (
            .O(N__23828),
            .I(N__23822));
    Odrv4 I__3362 (
            .O(N__23825),
            .I(\nx.n2992 ));
    LocalMux I__3361 (
            .O(N__23822),
            .I(\nx.n2992 ));
    CascadeMux I__3360 (
            .O(N__23817),
            .I(N__23814));
    InMux I__3359 (
            .O(N__23814),
            .I(N__23810));
    CascadeMux I__3358 (
            .O(N__23813),
            .I(N__23807));
    LocalMux I__3357 (
            .O(N__23810),
            .I(N__23804));
    InMux I__3356 (
            .O(N__23807),
            .I(N__23800));
    Span4Mux_v I__3355 (
            .O(N__23804),
            .I(N__23797));
    InMux I__3354 (
            .O(N__23803),
            .I(N__23794));
    LocalMux I__3353 (
            .O(N__23800),
            .I(\nx.n2989 ));
    Odrv4 I__3352 (
            .O(N__23797),
            .I(\nx.n2989 ));
    LocalMux I__3351 (
            .O(N__23794),
            .I(\nx.n2989 ));
    InMux I__3350 (
            .O(N__23787),
            .I(N__23784));
    LocalMux I__3349 (
            .O(N__23784),
            .I(N__23781));
    Odrv4 I__3348 (
            .O(N__23781),
            .I(\nx.n3056 ));
    CascadeMux I__3347 (
            .O(N__23778),
            .I(N__23773));
    CascadeMux I__3346 (
            .O(N__23777),
            .I(N__23770));
    InMux I__3345 (
            .O(N__23776),
            .I(N__23767));
    InMux I__3344 (
            .O(N__23773),
            .I(N__23764));
    InMux I__3343 (
            .O(N__23770),
            .I(N__23761));
    LocalMux I__3342 (
            .O(N__23767),
            .I(N__23758));
    LocalMux I__3341 (
            .O(N__23764),
            .I(\nx.n3104 ));
    LocalMux I__3340 (
            .O(N__23761),
            .I(\nx.n3104 ));
    Odrv4 I__3339 (
            .O(N__23758),
            .I(\nx.n3104 ));
    CascadeMux I__3338 (
            .O(N__23751),
            .I(\nx.n3088_cascade_ ));
    InMux I__3337 (
            .O(N__23748),
            .I(N__23745));
    LocalMux I__3336 (
            .O(N__23745),
            .I(N__23742));
    Odrv4 I__3335 (
            .O(N__23742),
            .I(\nx.n44_adj_690 ));
    InMux I__3334 (
            .O(N__23739),
            .I(N__23736));
    LocalMux I__3333 (
            .O(N__23736),
            .I(N__23733));
    Odrv4 I__3332 (
            .O(N__23733),
            .I(\nx.n3061 ));
    CascadeMux I__3331 (
            .O(N__23730),
            .I(N__23726));
    InMux I__3330 (
            .O(N__23729),
            .I(N__23723));
    InMux I__3329 (
            .O(N__23726),
            .I(N__23720));
    LocalMux I__3328 (
            .O(N__23723),
            .I(N__23717));
    LocalMux I__3327 (
            .O(N__23720),
            .I(N__23712));
    Span4Mux_v I__3326 (
            .O(N__23717),
            .I(N__23712));
    Odrv4 I__3325 (
            .O(N__23712),
            .I(\nx.n2994 ));
    CascadeMux I__3324 (
            .O(N__23709),
            .I(N__23706));
    InMux I__3323 (
            .O(N__23706),
            .I(N__23702));
    InMux I__3322 (
            .O(N__23705),
            .I(N__23699));
    LocalMux I__3321 (
            .O(N__23702),
            .I(N__23696));
    LocalMux I__3320 (
            .O(N__23699),
            .I(N__23690));
    Span4Mux_v I__3319 (
            .O(N__23696),
            .I(N__23690));
    InMux I__3318 (
            .O(N__23695),
            .I(N__23687));
    Odrv4 I__3317 (
            .O(N__23690),
            .I(\nx.n2991 ));
    LocalMux I__3316 (
            .O(N__23687),
            .I(\nx.n2991 ));
    InMux I__3315 (
            .O(N__23682),
            .I(N__23679));
    LocalMux I__3314 (
            .O(N__23679),
            .I(N__23676));
    Odrv4 I__3313 (
            .O(N__23676),
            .I(\nx.n3058 ));
    InMux I__3312 (
            .O(N__23673),
            .I(N__23670));
    LocalMux I__3311 (
            .O(N__23670),
            .I(N__23667));
    Span4Mux_h I__3310 (
            .O(N__23667),
            .I(N__23664));
    Odrv4 I__3309 (
            .O(N__23664),
            .I(\nx.n3161 ));
    InMux I__3308 (
            .O(N__23661),
            .I(N__23658));
    LocalMux I__3307 (
            .O(N__23658),
            .I(N__23655));
    Odrv4 I__3306 (
            .O(N__23655),
            .I(\nx.n12353 ));
    CascadeMux I__3305 (
            .O(N__23652),
            .I(N__23649));
    InMux I__3304 (
            .O(N__23649),
            .I(N__23646));
    LocalMux I__3303 (
            .O(N__23646),
            .I(N__23643));
    Span4Mux_h I__3302 (
            .O(N__23643),
            .I(N__23640));
    Odrv4 I__3301 (
            .O(N__23640),
            .I(\nx.n3160 ));
    InMux I__3300 (
            .O(N__23637),
            .I(N__23634));
    LocalMux I__3299 (
            .O(N__23634),
            .I(\nx.n12355 ));
    CascadeMux I__3298 (
            .O(N__23631),
            .I(\nx.n12357_cascade_ ));
    InMux I__3297 (
            .O(N__23628),
            .I(N__23625));
    LocalMux I__3296 (
            .O(N__23625),
            .I(N__23622));
    Span4Mux_v I__3295 (
            .O(N__23622),
            .I(N__23619));
    Odrv4 I__3294 (
            .O(N__23619),
            .I(\nx.n3159 ));
    InMux I__3293 (
            .O(N__23616),
            .I(N__23613));
    LocalMux I__3292 (
            .O(N__23613),
            .I(N__23610));
    Span4Mux_v I__3291 (
            .O(N__23610),
            .I(N__23607));
    Odrv4 I__3290 (
            .O(N__23607),
            .I(\nx.n3158 ));
    CascadeMux I__3289 (
            .O(N__23604),
            .I(\nx.n12359_cascade_ ));
    CascadeMux I__3288 (
            .O(N__23601),
            .I(N__23596));
    InMux I__3287 (
            .O(N__23600),
            .I(N__23591));
    InMux I__3286 (
            .O(N__23599),
            .I(N__23591));
    InMux I__3285 (
            .O(N__23596),
            .I(N__23588));
    LocalMux I__3284 (
            .O(N__23591),
            .I(N__23585));
    LocalMux I__3283 (
            .O(N__23588),
            .I(N__23582));
    Odrv4 I__3282 (
            .O(N__23585),
            .I(\nx.n3004 ));
    Odrv4 I__3281 (
            .O(N__23582),
            .I(\nx.n3004 ));
    CascadeMux I__3280 (
            .O(N__23577),
            .I(N__23573));
    InMux I__3279 (
            .O(N__23576),
            .I(N__23570));
    InMux I__3278 (
            .O(N__23573),
            .I(N__23567));
    LocalMux I__3277 (
            .O(N__23570),
            .I(N__23564));
    LocalMux I__3276 (
            .O(N__23567),
            .I(N__23561));
    Span4Mux_s3_h I__3275 (
            .O(N__23564),
            .I(N__23558));
    Span4Mux_v I__3274 (
            .O(N__23561),
            .I(N__23555));
    Odrv4 I__3273 (
            .O(N__23558),
            .I(\nx.n2988 ));
    Odrv4 I__3272 (
            .O(N__23555),
            .I(\nx.n2988 ));
    CascadeMux I__3271 (
            .O(N__23550),
            .I(\nx.n2988_cascade_ ));
    InMux I__3270 (
            .O(N__23547),
            .I(N__23544));
    LocalMux I__3269 (
            .O(N__23544),
            .I(N__23541));
    Odrv4 I__3268 (
            .O(N__23541),
            .I(\nx.n41_adj_686 ));
    CascadeMux I__3267 (
            .O(N__23538),
            .I(\nx.n2994_cascade_ ));
    CascadeMux I__3266 (
            .O(N__23535),
            .I(N__23531));
    CascadeMux I__3265 (
            .O(N__23534),
            .I(N__23528));
    InMux I__3264 (
            .O(N__23531),
            .I(N__23525));
    InMux I__3263 (
            .O(N__23528),
            .I(N__23522));
    LocalMux I__3262 (
            .O(N__23525),
            .I(N__23518));
    LocalMux I__3261 (
            .O(N__23522),
            .I(N__23515));
    InMux I__3260 (
            .O(N__23521),
            .I(N__23512));
    Span4Mux_v I__3259 (
            .O(N__23518),
            .I(N__23509));
    Odrv4 I__3258 (
            .O(N__23515),
            .I(\nx.n3002 ));
    LocalMux I__3257 (
            .O(N__23512),
            .I(\nx.n3002 ));
    Odrv4 I__3256 (
            .O(N__23509),
            .I(\nx.n3002 ));
    InMux I__3255 (
            .O(N__23502),
            .I(N__23499));
    LocalMux I__3254 (
            .O(N__23499),
            .I(N__23496));
    Odrv4 I__3253 (
            .O(N__23496),
            .I(\nx.n42_adj_684 ));
    InMux I__3252 (
            .O(N__23493),
            .I(N__23489));
    InMux I__3251 (
            .O(N__23492),
            .I(N__23486));
    LocalMux I__3250 (
            .O(N__23489),
            .I(N__23482));
    LocalMux I__3249 (
            .O(N__23486),
            .I(N__23479));
    CascadeMux I__3248 (
            .O(N__23485),
            .I(N__23476));
    Span4Mux_s3_h I__3247 (
            .O(N__23482),
            .I(N__23471));
    Span4Mux_h I__3246 (
            .O(N__23479),
            .I(N__23471));
    InMux I__3245 (
            .O(N__23476),
            .I(N__23468));
    Odrv4 I__3244 (
            .O(N__23471),
            .I(\nx.n3009 ));
    LocalMux I__3243 (
            .O(N__23468),
            .I(\nx.n3009 ));
    CascadeMux I__3242 (
            .O(N__23463),
            .I(\nx.n2985_cascade_ ));
    CascadeMux I__3241 (
            .O(N__23460),
            .I(N__23457));
    InMux I__3240 (
            .O(N__23457),
            .I(N__23453));
    InMux I__3239 (
            .O(N__23456),
            .I(N__23450));
    LocalMux I__3238 (
            .O(N__23453),
            .I(N__23447));
    LocalMux I__3237 (
            .O(N__23450),
            .I(N__23444));
    Span4Mux_s3_h I__3236 (
            .O(N__23447),
            .I(N__23440));
    Sp12to4 I__3235 (
            .O(N__23444),
            .I(N__23437));
    InMux I__3234 (
            .O(N__23443),
            .I(N__23434));
    Odrv4 I__3233 (
            .O(N__23440),
            .I(\nx.n2986 ));
    Odrv12 I__3232 (
            .O(N__23437),
            .I(\nx.n2986 ));
    LocalMux I__3231 (
            .O(N__23434),
            .I(\nx.n2986 ));
    InMux I__3230 (
            .O(N__23427),
            .I(N__23424));
    LocalMux I__3229 (
            .O(N__23424),
            .I(N__23421));
    Span4Mux_s3_h I__3228 (
            .O(N__23421),
            .I(N__23418));
    Odrv4 I__3227 (
            .O(N__23418),
            .I(\nx.n40_adj_683 ));
    CascadeMux I__3226 (
            .O(N__23415),
            .I(N__23412));
    InMux I__3225 (
            .O(N__23412),
            .I(N__23409));
    LocalMux I__3224 (
            .O(N__23409),
            .I(N__23406));
    Odrv4 I__3223 (
            .O(N__23406),
            .I(\nx.n43_adj_677 ));
    InMux I__3222 (
            .O(N__23403),
            .I(N__23400));
    LocalMux I__3221 (
            .O(N__23400),
            .I(\nx.n40_adj_678 ));
    CascadeMux I__3220 (
            .O(N__23397),
            .I(\nx.n47_cascade_ ));
    CascadeMux I__3219 (
            .O(N__23394),
            .I(\nx.n2918_cascade_ ));
    CascadeMux I__3218 (
            .O(N__23391),
            .I(N__23387));
    InMux I__3217 (
            .O(N__23390),
            .I(N__23383));
    InMux I__3216 (
            .O(N__23387),
            .I(N__23380));
    InMux I__3215 (
            .O(N__23386),
            .I(N__23377));
    LocalMux I__3214 (
            .O(N__23383),
            .I(N__23372));
    LocalMux I__3213 (
            .O(N__23380),
            .I(N__23372));
    LocalMux I__3212 (
            .O(N__23377),
            .I(N__23369));
    Span4Mux_v I__3211 (
            .O(N__23372),
            .I(N__23366));
    Odrv4 I__3210 (
            .O(N__23369),
            .I(\nx.n3000 ));
    Odrv4 I__3209 (
            .O(N__23366),
            .I(\nx.n3000 ));
    InMux I__3208 (
            .O(N__23361),
            .I(N__23358));
    LocalMux I__3207 (
            .O(N__23358),
            .I(\nx.n38_adj_676 ));
    CascadeMux I__3206 (
            .O(N__23355),
            .I(N__23351));
    CascadeMux I__3205 (
            .O(N__23354),
            .I(N__23348));
    InMux I__3204 (
            .O(N__23351),
            .I(N__23344));
    InMux I__3203 (
            .O(N__23348),
            .I(N__23341));
    InMux I__3202 (
            .O(N__23347),
            .I(N__23338));
    LocalMux I__3201 (
            .O(N__23344),
            .I(N__23335));
    LocalMux I__3200 (
            .O(N__23341),
            .I(N__23332));
    LocalMux I__3199 (
            .O(N__23338),
            .I(N__23329));
    Span12Mux_s3_h I__3198 (
            .O(N__23335),
            .I(N__23326));
    Odrv4 I__3197 (
            .O(N__23332),
            .I(\nx.n2996 ));
    Odrv4 I__3196 (
            .O(N__23329),
            .I(\nx.n2996 ));
    Odrv12 I__3195 (
            .O(N__23326),
            .I(\nx.n2996 ));
    InMux I__3194 (
            .O(N__23319),
            .I(N__23315));
    CascadeMux I__3193 (
            .O(N__23318),
            .I(N__23312));
    LocalMux I__3192 (
            .O(N__23315),
            .I(N__23308));
    InMux I__3191 (
            .O(N__23312),
            .I(N__23305));
    CascadeMux I__3190 (
            .O(N__23311),
            .I(N__23302));
    Span4Mux_s3_h I__3189 (
            .O(N__23308),
            .I(N__23297));
    LocalMux I__3188 (
            .O(N__23305),
            .I(N__23297));
    InMux I__3187 (
            .O(N__23302),
            .I(N__23294));
    Span4Mux_v I__3186 (
            .O(N__23297),
            .I(N__23291));
    LocalMux I__3185 (
            .O(N__23294),
            .I(N__23288));
    Odrv4 I__3184 (
            .O(N__23291),
            .I(\nx.n2997 ));
    Odrv4 I__3183 (
            .O(N__23288),
            .I(\nx.n2997 ));
    CascadeMux I__3182 (
            .O(N__23283),
            .I(N__23279));
    CascadeMux I__3181 (
            .O(N__23282),
            .I(N__23276));
    InMux I__3180 (
            .O(N__23279),
            .I(N__23273));
    InMux I__3179 (
            .O(N__23276),
            .I(N__23270));
    LocalMux I__3178 (
            .O(N__23273),
            .I(N__23267));
    LocalMux I__3177 (
            .O(N__23270),
            .I(N__23264));
    Span4Mux_h I__3176 (
            .O(N__23267),
            .I(N__23260));
    Span4Mux_v I__3175 (
            .O(N__23264),
            .I(N__23257));
    InMux I__3174 (
            .O(N__23263),
            .I(N__23254));
    Odrv4 I__3173 (
            .O(N__23260),
            .I(\nx.n2987 ));
    Odrv4 I__3172 (
            .O(N__23257),
            .I(\nx.n2987 ));
    LocalMux I__3171 (
            .O(N__23254),
            .I(\nx.n2987 ));
    CascadeMux I__3170 (
            .O(N__23247),
            .I(N__23243));
    InMux I__3169 (
            .O(N__23246),
            .I(N__23240));
    InMux I__3168 (
            .O(N__23243),
            .I(N__23237));
    LocalMux I__3167 (
            .O(N__23240),
            .I(N__23234));
    LocalMux I__3166 (
            .O(N__23237),
            .I(N__23230));
    Span12Mux_s3_h I__3165 (
            .O(N__23234),
            .I(N__23227));
    InMux I__3164 (
            .O(N__23233),
            .I(N__23224));
    Span4Mux_v I__3163 (
            .O(N__23230),
            .I(N__23221));
    Odrv12 I__3162 (
            .O(N__23227),
            .I(\nx.n3005 ));
    LocalMux I__3161 (
            .O(N__23224),
            .I(\nx.n3005 ));
    Odrv4 I__3160 (
            .O(N__23221),
            .I(\nx.n3005 ));
    InMux I__3159 (
            .O(N__23214),
            .I(N__23210));
    InMux I__3158 (
            .O(N__23213),
            .I(N__23207));
    LocalMux I__3157 (
            .O(N__23210),
            .I(N__23202));
    LocalMux I__3156 (
            .O(N__23207),
            .I(N__23202));
    Odrv4 I__3155 (
            .O(N__23202),
            .I(neo_pixel_transmitter_t0_7));
    InMux I__3154 (
            .O(N__23199),
            .I(N__23196));
    LocalMux I__3153 (
            .O(N__23196),
            .I(\nx.n26 ));
    CascadeMux I__3152 (
            .O(N__23193),
            .I(N__23189));
    InMux I__3151 (
            .O(N__23192),
            .I(N__23186));
    InMux I__3150 (
            .O(N__23189),
            .I(N__23183));
    LocalMux I__3149 (
            .O(N__23186),
            .I(N__23179));
    LocalMux I__3148 (
            .O(N__23183),
            .I(N__23176));
    InMux I__3147 (
            .O(N__23182),
            .I(N__23173));
    Span4Mux_s3_h I__3146 (
            .O(N__23179),
            .I(N__23168));
    Span4Mux_v I__3145 (
            .O(N__23176),
            .I(N__23168));
    LocalMux I__3144 (
            .O(N__23173),
            .I(\nx.n3006 ));
    Odrv4 I__3143 (
            .O(N__23168),
            .I(\nx.n3006 ));
    CascadeMux I__3142 (
            .O(N__23163),
            .I(\nx.n2899_cascade_ ));
    CascadeMux I__3141 (
            .O(N__23160),
            .I(N__23156));
    InMux I__3140 (
            .O(N__23159),
            .I(N__23153));
    InMux I__3139 (
            .O(N__23156),
            .I(N__23150));
    LocalMux I__3138 (
            .O(N__23153),
            .I(N__23147));
    LocalMux I__3137 (
            .O(N__23150),
            .I(N__23144));
    Span4Mux_s3_h I__3136 (
            .O(N__23147),
            .I(N__23138));
    Span4Mux_v I__3135 (
            .O(N__23144),
            .I(N__23138));
    InMux I__3134 (
            .O(N__23143),
            .I(N__23135));
    Odrv4 I__3133 (
            .O(N__23138),
            .I(\nx.n2998 ));
    LocalMux I__3132 (
            .O(N__23135),
            .I(\nx.n2998 ));
    CascadeMux I__3131 (
            .O(N__23130),
            .I(\nx.n2894_cascade_ ));
    CascadeMux I__3130 (
            .O(N__23127),
            .I(N__23123));
    CascadeMux I__3129 (
            .O(N__23126),
            .I(N__23120));
    InMux I__3128 (
            .O(N__23123),
            .I(N__23117));
    InMux I__3127 (
            .O(N__23120),
            .I(N__23114));
    LocalMux I__3126 (
            .O(N__23117),
            .I(N__23111));
    LocalMux I__3125 (
            .O(N__23114),
            .I(N__23108));
    Span12Mux_s3_h I__3124 (
            .O(N__23111),
            .I(N__23105));
    Span4Mux_v I__3123 (
            .O(N__23108),
            .I(N__23102));
    Odrv12 I__3122 (
            .O(N__23105),
            .I(\nx.n2985 ));
    Odrv4 I__3121 (
            .O(N__23102),
            .I(\nx.n2985 ));
    CascadeMux I__3120 (
            .O(N__23097),
            .I(N__23094));
    InMux I__3119 (
            .O(N__23094),
            .I(N__23091));
    LocalMux I__3118 (
            .O(N__23091),
            .I(N__23088));
    Span4Mux_v I__3117 (
            .O(N__23088),
            .I(N__23085));
    Span4Mux_h I__3116 (
            .O(N__23085),
            .I(N__23082));
    Odrv4 I__3115 (
            .O(N__23082),
            .I(\nx.n5 ));
    CascadeMux I__3114 (
            .O(N__23079),
            .I(N__23076));
    InMux I__3113 (
            .O(N__23076),
            .I(N__23070));
    InMux I__3112 (
            .O(N__23075),
            .I(N__23070));
    LocalMux I__3111 (
            .O(N__23070),
            .I(neo_pixel_transmitter_t0_25));
    InMux I__3110 (
            .O(N__23067),
            .I(N__23064));
    LocalMux I__3109 (
            .O(N__23064),
            .I(N__23061));
    Span4Mux_v I__3108 (
            .O(N__23061),
            .I(N__23058));
    Odrv4 I__3107 (
            .O(N__23058),
            .I(\nx.n8 ));
    InMux I__3106 (
            .O(N__23055),
            .I(N__23049));
    InMux I__3105 (
            .O(N__23054),
            .I(N__23049));
    LocalMux I__3104 (
            .O(N__23049),
            .I(neo_pixel_transmitter_t0_18));
    InMux I__3103 (
            .O(N__23046),
            .I(N__23043));
    LocalMux I__3102 (
            .O(N__23043),
            .I(N__23040));
    Span4Mux_v I__3101 (
            .O(N__23040),
            .I(N__23037));
    Odrv4 I__3100 (
            .O(N__23037),
            .I(\nx.n15 ));
    InMux I__3099 (
            .O(N__23034),
            .I(N__23031));
    LocalMux I__3098 (
            .O(N__23031),
            .I(N__23026));
    InMux I__3097 (
            .O(N__23030),
            .I(N__23023));
    InMux I__3096 (
            .O(N__23029),
            .I(N__23020));
    Span12Mux_s8_v I__3095 (
            .O(N__23026),
            .I(N__23017));
    LocalMux I__3094 (
            .O(N__23023),
            .I(timer_28));
    LocalMux I__3093 (
            .O(N__23020),
            .I(timer_28));
    Odrv12 I__3092 (
            .O(N__23017),
            .I(timer_28));
    CascadeMux I__3091 (
            .O(N__23010),
            .I(N__23007));
    InMux I__3090 (
            .O(N__23007),
            .I(N__23001));
    InMux I__3089 (
            .O(N__23006),
            .I(N__23001));
    LocalMux I__3088 (
            .O(N__23001),
            .I(neo_pixel_transmitter_t0_28));
    CascadeMux I__3087 (
            .O(N__22998),
            .I(\nx.n2995_cascade_ ));
    InMux I__3086 (
            .O(N__22995),
            .I(N__22992));
    LocalMux I__3085 (
            .O(N__22992),
            .I(\nx.n44_adj_681 ));
    CascadeMux I__3084 (
            .O(N__22989),
            .I(\nx.n33_adj_682_cascade_ ));
    InMux I__3083 (
            .O(N__22986),
            .I(N__22983));
    LocalMux I__3082 (
            .O(N__22983),
            .I(N__22980));
    Span4Mux_s3_h I__3081 (
            .O(N__22980),
            .I(N__22977));
    Odrv4 I__3080 (
            .O(N__22977),
            .I(\nx.n48 ));
    CascadeMux I__3079 (
            .O(N__22974),
            .I(N__22971));
    InMux I__3078 (
            .O(N__22971),
            .I(N__22966));
    InMux I__3077 (
            .O(N__22970),
            .I(N__22963));
    InMux I__3076 (
            .O(N__22969),
            .I(N__22960));
    LocalMux I__3075 (
            .O(N__22966),
            .I(N__22957));
    LocalMux I__3074 (
            .O(N__22963),
            .I(timer_21));
    LocalMux I__3073 (
            .O(N__22960),
            .I(timer_21));
    Odrv12 I__3072 (
            .O(N__22957),
            .I(timer_21));
    CascadeMux I__3071 (
            .O(N__22950),
            .I(N__22947));
    InMux I__3070 (
            .O(N__22947),
            .I(N__22944));
    LocalMux I__3069 (
            .O(N__22944),
            .I(N__22939));
    InMux I__3068 (
            .O(N__22943),
            .I(N__22936));
    InMux I__3067 (
            .O(N__22942),
            .I(N__22933));
    Span4Mux_v I__3066 (
            .O(N__22939),
            .I(N__22930));
    LocalMux I__3065 (
            .O(N__22936),
            .I(timer_13));
    LocalMux I__3064 (
            .O(N__22933),
            .I(timer_13));
    Odrv4 I__3063 (
            .O(N__22930),
            .I(timer_13));
    InMux I__3062 (
            .O(N__22923),
            .I(N__22919));
    InMux I__3061 (
            .O(N__22922),
            .I(N__22916));
    LocalMux I__3060 (
            .O(N__22919),
            .I(neo_pixel_transmitter_t0_11));
    LocalMux I__3059 (
            .O(N__22916),
            .I(neo_pixel_transmitter_t0_11));
    InMux I__3058 (
            .O(N__22911),
            .I(N__22908));
    LocalMux I__3057 (
            .O(N__22908),
            .I(N__22905));
    Span4Mux_h I__3056 (
            .O(N__22905),
            .I(N__22902));
    Odrv4 I__3055 (
            .O(N__22902),
            .I(\nx.n22_adj_618 ));
    InMux I__3054 (
            .O(N__22899),
            .I(N__22893));
    InMux I__3053 (
            .O(N__22898),
            .I(N__22893));
    LocalMux I__3052 (
            .O(N__22893),
            .I(neo_pixel_transmitter_t0_13));
    InMux I__3051 (
            .O(N__22890),
            .I(N__22887));
    LocalMux I__3050 (
            .O(N__22887),
            .I(N__22884));
    Odrv4 I__3049 (
            .O(N__22884),
            .I(\nx.n20 ));
    CascadeMux I__3048 (
            .O(N__22881),
            .I(N__22878));
    InMux I__3047 (
            .O(N__22878),
            .I(N__22874));
    InMux I__3046 (
            .O(N__22877),
            .I(N__22871));
    LocalMux I__3045 (
            .O(N__22874),
            .I(N__22867));
    LocalMux I__3044 (
            .O(N__22871),
            .I(N__22864));
    InMux I__3043 (
            .O(N__22870),
            .I(N__22861));
    Span4Mux_v I__3042 (
            .O(N__22867),
            .I(N__22858));
    Odrv4 I__3041 (
            .O(N__22864),
            .I(timer_7));
    LocalMux I__3040 (
            .O(N__22861),
            .I(timer_7));
    Odrv4 I__3039 (
            .O(N__22858),
            .I(timer_7));
    InMux I__3038 (
            .O(N__22851),
            .I(N__22848));
    LocalMux I__3037 (
            .O(N__22848),
            .I(N__22845));
    Span4Mux_s3_h I__3036 (
            .O(N__22845),
            .I(N__22842));
    Odrv4 I__3035 (
            .O(N__22842),
            .I(\nx.n13159 ));
    CascadeMux I__3034 (
            .O(N__22839),
            .I(N__22836));
    InMux I__3033 (
            .O(N__22836),
            .I(N__22830));
    InMux I__3032 (
            .O(N__22835),
            .I(N__22830));
    LocalMux I__3031 (
            .O(N__22830),
            .I(neo_pixel_transmitter_t0_21));
    InMux I__3030 (
            .O(N__22827),
            .I(N__22824));
    LocalMux I__3029 (
            .O(N__22824),
            .I(N__22821));
    Span4Mux_v I__3028 (
            .O(N__22821),
            .I(N__22818));
    Odrv4 I__3027 (
            .O(N__22818),
            .I(\nx.n12 ));
    CascadeMux I__3026 (
            .O(N__22815),
            .I(N__22812));
    InMux I__3025 (
            .O(N__22812),
            .I(N__22809));
    LocalMux I__3024 (
            .O(N__22809),
            .I(N__22804));
    InMux I__3023 (
            .O(N__22808),
            .I(N__22801));
    InMux I__3022 (
            .O(N__22807),
            .I(N__22798));
    Span4Mux_v I__3021 (
            .O(N__22804),
            .I(N__22795));
    LocalMux I__3020 (
            .O(N__22801),
            .I(timer_25));
    LocalMux I__3019 (
            .O(N__22798),
            .I(timer_25));
    Odrv4 I__3018 (
            .O(N__22795),
            .I(timer_25));
    CascadeMux I__3017 (
            .O(N__22788),
            .I(N__22785));
    InMux I__3016 (
            .O(N__22785),
            .I(N__22780));
    InMux I__3015 (
            .O(N__22784),
            .I(N__22777));
    InMux I__3014 (
            .O(N__22783),
            .I(N__22774));
    LocalMux I__3013 (
            .O(N__22780),
            .I(N__22771));
    LocalMux I__3012 (
            .O(N__22777),
            .I(timer_18));
    LocalMux I__3011 (
            .O(N__22774),
            .I(timer_18));
    Odrv12 I__3010 (
            .O(N__22771),
            .I(timer_18));
    InMux I__3009 (
            .O(N__22764),
            .I(N__22761));
    LocalMux I__3008 (
            .O(N__22761),
            .I(N__22758));
    Span4Mux_v I__3007 (
            .O(N__22758),
            .I(N__22755));
    Odrv4 I__3006 (
            .O(N__22755),
            .I(\nx.n31_adj_650 ));
    CascadeMux I__3005 (
            .O(N__22752),
            .I(N__22749));
    InMux I__3004 (
            .O(N__22749),
            .I(N__22746));
    LocalMux I__3003 (
            .O(N__22746),
            .I(N__22743));
    Span4Mux_v I__3002 (
            .O(N__22743),
            .I(N__22740));
    Odrv4 I__3001 (
            .O(N__22740),
            .I(\nx.n16_adj_661 ));
    InMux I__3000 (
            .O(N__22737),
            .I(N__22733));
    InMux I__2999 (
            .O(N__22736),
            .I(N__22730));
    LocalMux I__2998 (
            .O(N__22733),
            .I(N__22726));
    LocalMux I__2997 (
            .O(N__22730),
            .I(N__22723));
    InMux I__2996 (
            .O(N__22729),
            .I(N__22720));
    Span4Mux_v I__2995 (
            .O(N__22726),
            .I(N__22717));
    Odrv4 I__2994 (
            .O(N__22723),
            .I(timer_17));
    LocalMux I__2993 (
            .O(N__22720),
            .I(timer_17));
    Odrv4 I__2992 (
            .O(N__22717),
            .I(timer_17));
    CascadeMux I__2991 (
            .O(N__22710),
            .I(N__22707));
    InMux I__2990 (
            .O(N__22707),
            .I(N__22701));
    InMux I__2989 (
            .O(N__22706),
            .I(N__22701));
    LocalMux I__2988 (
            .O(N__22701),
            .I(neo_pixel_transmitter_t0_17));
    CascadeMux I__2987 (
            .O(N__22698),
            .I(N__22695));
    InMux I__2986 (
            .O(N__22695),
            .I(N__22690));
    InMux I__2985 (
            .O(N__22694),
            .I(N__22687));
    InMux I__2984 (
            .O(N__22693),
            .I(N__22684));
    LocalMux I__2983 (
            .O(N__22690),
            .I(N__22681));
    LocalMux I__2982 (
            .O(N__22687),
            .I(timer_2));
    LocalMux I__2981 (
            .O(N__22684),
            .I(timer_2));
    Odrv12 I__2980 (
            .O(N__22681),
            .I(timer_2));
    InMux I__2979 (
            .O(N__22674),
            .I(N__22670));
    InMux I__2978 (
            .O(N__22673),
            .I(N__22667));
    LocalMux I__2977 (
            .O(N__22670),
            .I(neo_pixel_transmitter_t0_2));
    LocalMux I__2976 (
            .O(N__22667),
            .I(neo_pixel_transmitter_t0_2));
    InMux I__2975 (
            .O(N__22662),
            .I(N__22658));
    InMux I__2974 (
            .O(N__22661),
            .I(N__22655));
    LocalMux I__2973 (
            .O(N__22658),
            .I(N__22651));
    LocalMux I__2972 (
            .O(N__22655),
            .I(N__22648));
    InMux I__2971 (
            .O(N__22654),
            .I(N__22645));
    Span4Mux_v I__2970 (
            .O(N__22651),
            .I(N__22642));
    Odrv4 I__2969 (
            .O(N__22648),
            .I(timer_29));
    LocalMux I__2968 (
            .O(N__22645),
            .I(timer_29));
    Odrv4 I__2967 (
            .O(N__22642),
            .I(timer_29));
    CascadeMux I__2966 (
            .O(N__22635),
            .I(N__22632));
    InMux I__2965 (
            .O(N__22632),
            .I(N__22627));
    InMux I__2964 (
            .O(N__22631),
            .I(N__22624));
    InMux I__2963 (
            .O(N__22630),
            .I(N__22621));
    LocalMux I__2962 (
            .O(N__22627),
            .I(N__22618));
    LocalMux I__2961 (
            .O(N__22624),
            .I(timer_9));
    LocalMux I__2960 (
            .O(N__22621),
            .I(timer_9));
    Odrv12 I__2959 (
            .O(N__22618),
            .I(timer_9));
    InMux I__2958 (
            .O(N__22611),
            .I(N__22607));
    InMux I__2957 (
            .O(N__22610),
            .I(N__22604));
    LocalMux I__2956 (
            .O(N__22607),
            .I(N__22601));
    LocalMux I__2955 (
            .O(N__22604),
            .I(neo_pixel_transmitter_t0_10));
    Odrv4 I__2954 (
            .O(N__22601),
            .I(neo_pixel_transmitter_t0_10));
    InMux I__2953 (
            .O(N__22596),
            .I(N__22593));
    LocalMux I__2952 (
            .O(N__22593),
            .I(N__22590));
    Span4Mux_v I__2951 (
            .O(N__22590),
            .I(N__22587));
    Odrv4 I__2950 (
            .O(N__22587),
            .I(\nx.n23_adj_617 ));
    InMux I__2949 (
            .O(N__22584),
            .I(N__22578));
    InMux I__2948 (
            .O(N__22583),
            .I(N__22578));
    LocalMux I__2947 (
            .O(N__22578),
            .I(neo_pixel_transmitter_t0_29));
    CascadeMux I__2946 (
            .O(N__22575),
            .I(N__22572));
    InMux I__2945 (
            .O(N__22572),
            .I(N__22569));
    LocalMux I__2944 (
            .O(N__22569),
            .I(N__22566));
    Span4Mux_s3_h I__2943 (
            .O(N__22566),
            .I(N__22563));
    Span4Mux_v I__2942 (
            .O(N__22563),
            .I(N__22560));
    Odrv4 I__2941 (
            .O(N__22560),
            .I(\nx.n4 ));
    CascadeMux I__2940 (
            .O(N__22557),
            .I(N__22554));
    InMux I__2939 (
            .O(N__22554),
            .I(N__22549));
    InMux I__2938 (
            .O(N__22553),
            .I(N__22546));
    InMux I__2937 (
            .O(N__22552),
            .I(N__22543));
    LocalMux I__2936 (
            .O(N__22549),
            .I(N__22540));
    LocalMux I__2935 (
            .O(N__22546),
            .I(timer_11));
    LocalMux I__2934 (
            .O(N__22543),
            .I(timer_11));
    Odrv12 I__2933 (
            .O(N__22540),
            .I(timer_11));
    InMux I__2932 (
            .O(N__22533),
            .I(\nx.n10588 ));
    InMux I__2931 (
            .O(N__22530),
            .I(bfn_3_32_0_));
    InMux I__2930 (
            .O(N__22527),
            .I(\nx.n10590 ));
    InMux I__2929 (
            .O(N__22524),
            .I(\nx.n10591 ));
    InMux I__2928 (
            .O(N__22521),
            .I(N__22518));
    LocalMux I__2927 (
            .O(N__22518),
            .I(N__22513));
    CascadeMux I__2926 (
            .O(N__22517),
            .I(N__22510));
    CascadeMux I__2925 (
            .O(N__22516),
            .I(N__22507));
    Span4Mux_s2_v I__2924 (
            .O(N__22513),
            .I(N__22504));
    InMux I__2923 (
            .O(N__22510),
            .I(N__22501));
    InMux I__2922 (
            .O(N__22507),
            .I(N__22498));
    Odrv4 I__2921 (
            .O(N__22504),
            .I(\nx.n1303 ));
    LocalMux I__2920 (
            .O(N__22501),
            .I(\nx.n1303 ));
    LocalMux I__2919 (
            .O(N__22498),
            .I(\nx.n1303 ));
    CascadeMux I__2918 (
            .O(N__22491),
            .I(N__22488));
    InMux I__2917 (
            .O(N__22488),
            .I(N__22485));
    LocalMux I__2916 (
            .O(N__22485),
            .I(\nx.n1370 ));
    InMux I__2915 (
            .O(N__22482),
            .I(N__22476));
    InMux I__2914 (
            .O(N__22481),
            .I(N__22476));
    LocalMux I__2913 (
            .O(N__22476),
            .I(\nx.n1400 ));
    CascadeMux I__2912 (
            .O(N__22473),
            .I(N__22470));
    InMux I__2911 (
            .O(N__22470),
            .I(N__22467));
    LocalMux I__2910 (
            .O(N__22467),
            .I(N__22464));
    Span4Mux_v I__2909 (
            .O(N__22464),
            .I(N__22461));
    Span4Mux_v I__2908 (
            .O(N__22461),
            .I(N__22458));
    Odrv4 I__2907 (
            .O(N__22458),
            .I(\nx.n3 ));
    InMux I__2906 (
            .O(N__22455),
            .I(N__22451));
    InMux I__2905 (
            .O(N__22454),
            .I(N__22448));
    LocalMux I__2904 (
            .O(N__22451),
            .I(N__22445));
    LocalMux I__2903 (
            .O(N__22448),
            .I(N__22441));
    Span4Mux_v I__2902 (
            .O(N__22445),
            .I(N__22438));
    InMux I__2901 (
            .O(N__22444),
            .I(N__22435));
    Span4Mux_v I__2900 (
            .O(N__22441),
            .I(N__22432));
    Odrv4 I__2899 (
            .O(N__22438),
            .I(timer_30));
    LocalMux I__2898 (
            .O(N__22435),
            .I(timer_30));
    Odrv4 I__2897 (
            .O(N__22432),
            .I(timer_30));
    InMux I__2896 (
            .O(N__22425),
            .I(N__22419));
    InMux I__2895 (
            .O(N__22424),
            .I(N__22419));
    LocalMux I__2894 (
            .O(N__22419),
            .I(neo_pixel_transmitter_t0_30));
    InMux I__2893 (
            .O(N__22416),
            .I(N__22413));
    LocalMux I__2892 (
            .O(N__22413),
            .I(N__22410));
    Span4Mux_h I__2891 (
            .O(N__22410),
            .I(N__22407));
    Odrv4 I__2890 (
            .O(N__22407),
            .I(\nx.n1272 ));
    CascadeMux I__2889 (
            .O(N__22404),
            .I(N__22400));
    CascadeMux I__2888 (
            .O(N__22403),
            .I(N__22397));
    InMux I__2887 (
            .O(N__22400),
            .I(N__22393));
    InMux I__2886 (
            .O(N__22397),
            .I(N__22390));
    InMux I__2885 (
            .O(N__22396),
            .I(N__22387));
    LocalMux I__2884 (
            .O(N__22393),
            .I(\nx.n1205 ));
    LocalMux I__2883 (
            .O(N__22390),
            .I(\nx.n1205 ));
    LocalMux I__2882 (
            .O(N__22387),
            .I(\nx.n1205 ));
    CascadeMux I__2881 (
            .O(N__22380),
            .I(N__22374));
    CascadeMux I__2880 (
            .O(N__22379),
            .I(N__22371));
    CascadeMux I__2879 (
            .O(N__22378),
            .I(N__22368));
    InMux I__2878 (
            .O(N__22377),
            .I(N__22355));
    InMux I__2877 (
            .O(N__22374),
            .I(N__22355));
    InMux I__2876 (
            .O(N__22371),
            .I(N__22355));
    InMux I__2875 (
            .O(N__22368),
            .I(N__22355));
    InMux I__2874 (
            .O(N__22367),
            .I(N__22350));
    InMux I__2873 (
            .O(N__22366),
            .I(N__22350));
    InMux I__2872 (
            .O(N__22365),
            .I(N__22345));
    InMux I__2871 (
            .O(N__22364),
            .I(N__22345));
    LocalMux I__2870 (
            .O(N__22355),
            .I(N__22342));
    LocalMux I__2869 (
            .O(N__22350),
            .I(\nx.n1235 ));
    LocalMux I__2868 (
            .O(N__22345),
            .I(\nx.n1235 ));
    Odrv4 I__2867 (
            .O(N__22342),
            .I(\nx.n1235 ));
    InMux I__2866 (
            .O(N__22335),
            .I(N__22332));
    LocalMux I__2865 (
            .O(N__22332),
            .I(\nx.n1377 ));
    InMux I__2864 (
            .O(N__22329),
            .I(bfn_3_31_0_));
    InMux I__2863 (
            .O(N__22326),
            .I(\nx.n10582 ));
    InMux I__2862 (
            .O(N__22323),
            .I(\nx.n10583 ));
    InMux I__2861 (
            .O(N__22320),
            .I(\nx.n10584 ));
    InMux I__2860 (
            .O(N__22317),
            .I(\nx.n10585 ));
    InMux I__2859 (
            .O(N__22314),
            .I(\nx.n10586 ));
    InMux I__2858 (
            .O(N__22311),
            .I(\nx.n10587 ));
    InMux I__2857 (
            .O(N__22308),
            .I(N__22305));
    LocalMux I__2856 (
            .O(N__22305),
            .I(N__22302));
    Span4Mux_v I__2855 (
            .O(N__22302),
            .I(N__22299));
    Odrv4 I__2854 (
            .O(N__22299),
            .I(\nx.n3053 ));
    InMux I__2853 (
            .O(N__22296),
            .I(bfn_3_29_0_));
    InMux I__2852 (
            .O(N__22293),
            .I(N__22290));
    LocalMux I__2851 (
            .O(N__22290),
            .I(\nx.n3052 ));
    InMux I__2850 (
            .O(N__22287),
            .I(\nx.n10886 ));
    InMux I__2849 (
            .O(N__22284),
            .I(\nx.n10887 ));
    CascadeMux I__2848 (
            .O(N__22281),
            .I(N__22278));
    InMux I__2847 (
            .O(N__22278),
            .I(N__22274));
    InMux I__2846 (
            .O(N__22277),
            .I(N__22271));
    LocalMux I__2845 (
            .O(N__22274),
            .I(N__22268));
    LocalMux I__2844 (
            .O(N__22271),
            .I(N__22265));
    Span4Mux_s2_h I__2843 (
            .O(N__22268),
            .I(N__22262));
    Odrv4 I__2842 (
            .O(N__22265),
            .I(\nx.n3083 ));
    Odrv4 I__2841 (
            .O(N__22262),
            .I(\nx.n3083 ));
    InMux I__2840 (
            .O(N__22257),
            .I(N__22254));
    LocalMux I__2839 (
            .O(N__22254),
            .I(\nx.n45_adj_707 ));
    CascadeMux I__2838 (
            .O(N__22251),
            .I(\nx.n11_adj_628_cascade_ ));
    InMux I__2837 (
            .O(N__22248),
            .I(N__22245));
    LocalMux I__2836 (
            .O(N__22245),
            .I(\nx.n16_adj_627 ));
    InMux I__2835 (
            .O(N__22242),
            .I(N__22237));
    InMux I__2834 (
            .O(N__22241),
            .I(N__22234));
    InMux I__2833 (
            .O(N__22240),
            .I(N__22231));
    LocalMux I__2832 (
            .O(N__22237),
            .I(\nx.n1307 ));
    LocalMux I__2831 (
            .O(N__22234),
            .I(\nx.n1307 ));
    LocalMux I__2830 (
            .O(N__22231),
            .I(\nx.n1307 ));
    CascadeMux I__2829 (
            .O(N__22224),
            .I(\nx.n1334_cascade_ ));
    InMux I__2828 (
            .O(N__22221),
            .I(N__22218));
    LocalMux I__2827 (
            .O(N__22218),
            .I(\nx.n1374 ));
    InMux I__2826 (
            .O(N__22215),
            .I(N__22212));
    LocalMux I__2825 (
            .O(N__22212),
            .I(N__22209));
    Span4Mux_v I__2824 (
            .O(N__22209),
            .I(N__22206));
    Odrv4 I__2823 (
            .O(N__22206),
            .I(\nx.n1277 ));
    CascadeMux I__2822 (
            .O(N__22203),
            .I(N__22199));
    InMux I__2821 (
            .O(N__22202),
            .I(N__22196));
    InMux I__2820 (
            .O(N__22199),
            .I(N__22193));
    LocalMux I__2819 (
            .O(N__22196),
            .I(\nx.n1309 ));
    LocalMux I__2818 (
            .O(N__22193),
            .I(\nx.n1309 ));
    InMux I__2817 (
            .O(N__22188),
            .I(N__22185));
    LocalMux I__2816 (
            .O(N__22185),
            .I(\nx.n1376 ));
    CascadeMux I__2815 (
            .O(N__22182),
            .I(\nx.n1309_cascade_ ));
    InMux I__2814 (
            .O(N__22179),
            .I(bfn_3_28_0_));
    InMux I__2813 (
            .O(N__22176),
            .I(\nx.n10878 ));
    InMux I__2812 (
            .O(N__22173),
            .I(N__22170));
    LocalMux I__2811 (
            .O(N__22170),
            .I(\nx.n3059 ));
    InMux I__2810 (
            .O(N__22167),
            .I(\nx.n10879 ));
    InMux I__2809 (
            .O(N__22164),
            .I(\nx.n10880 ));
    InMux I__2808 (
            .O(N__22161),
            .I(\nx.n10881 ));
    InMux I__2807 (
            .O(N__22158),
            .I(\nx.n10882 ));
    InMux I__2806 (
            .O(N__22155),
            .I(N__22152));
    LocalMux I__2805 (
            .O(N__22152),
            .I(N__22149));
    Span4Mux_v I__2804 (
            .O(N__22149),
            .I(N__22146));
    Odrv4 I__2803 (
            .O(N__22146),
            .I(\nx.n3055 ));
    InMux I__2802 (
            .O(N__22143),
            .I(\nx.n10883 ));
    InMux I__2801 (
            .O(N__22140),
            .I(N__22137));
    LocalMux I__2800 (
            .O(N__22137),
            .I(N__22134));
    Span4Mux_v I__2799 (
            .O(N__22134),
            .I(N__22131));
    Odrv4 I__2798 (
            .O(N__22131),
            .I(\nx.n3054 ));
    InMux I__2797 (
            .O(N__22128),
            .I(\nx.n10884 ));
    CascadeMux I__2796 (
            .O(N__22125),
            .I(N__22122));
    InMux I__2795 (
            .O(N__22122),
            .I(N__22119));
    LocalMux I__2794 (
            .O(N__22119),
            .I(N__22116));
    Span4Mux_v I__2793 (
            .O(N__22116),
            .I(N__22113));
    Odrv4 I__2792 (
            .O(N__22113),
            .I(\nx.n3070 ));
    InMux I__2791 (
            .O(N__22110),
            .I(\nx.n10868 ));
    InMux I__2790 (
            .O(N__22107),
            .I(N__22104));
    LocalMux I__2789 (
            .O(N__22104),
            .I(N__22101));
    Span4Mux_s2_h I__2788 (
            .O(N__22101),
            .I(N__22098));
    Odrv4 I__2787 (
            .O(N__22098),
            .I(\nx.n3069 ));
    InMux I__2786 (
            .O(N__22095),
            .I(bfn_3_27_0_));
    CascadeMux I__2785 (
            .O(N__22092),
            .I(N__22089));
    InMux I__2784 (
            .O(N__22089),
            .I(N__22086));
    LocalMux I__2783 (
            .O(N__22086),
            .I(N__22081));
    InMux I__2782 (
            .O(N__22085),
            .I(N__22078));
    InMux I__2781 (
            .O(N__22084),
            .I(N__22075));
    Span4Mux_v I__2780 (
            .O(N__22081),
            .I(N__22072));
    LocalMux I__2779 (
            .O(N__22078),
            .I(\nx.n3001 ));
    LocalMux I__2778 (
            .O(N__22075),
            .I(\nx.n3001 ));
    Odrv4 I__2777 (
            .O(N__22072),
            .I(\nx.n3001 ));
    InMux I__2776 (
            .O(N__22065),
            .I(N__22062));
    LocalMux I__2775 (
            .O(N__22062),
            .I(N__22059));
    Span4Mux_s2_h I__2774 (
            .O(N__22059),
            .I(N__22056));
    Odrv4 I__2773 (
            .O(N__22056),
            .I(\nx.n3068 ));
    InMux I__2772 (
            .O(N__22053),
            .I(\nx.n10870 ));
    CascadeMux I__2771 (
            .O(N__22050),
            .I(N__22047));
    InMux I__2770 (
            .O(N__22047),
            .I(N__22044));
    LocalMux I__2769 (
            .O(N__22044),
            .I(\nx.n3067 ));
    InMux I__2768 (
            .O(N__22041),
            .I(\nx.n10871 ));
    CascadeMux I__2767 (
            .O(N__22038),
            .I(N__22035));
    InMux I__2766 (
            .O(N__22035),
            .I(N__22032));
    LocalMux I__2765 (
            .O(N__22032),
            .I(N__22027));
    InMux I__2764 (
            .O(N__22031),
            .I(N__22024));
    InMux I__2763 (
            .O(N__22030),
            .I(N__22021));
    Span4Mux_v I__2762 (
            .O(N__22027),
            .I(N__22018));
    LocalMux I__2761 (
            .O(N__22024),
            .I(\nx.n2999 ));
    LocalMux I__2760 (
            .O(N__22021),
            .I(\nx.n2999 ));
    Odrv4 I__2759 (
            .O(N__22018),
            .I(\nx.n2999 ));
    CascadeMux I__2758 (
            .O(N__22011),
            .I(N__22008));
    InMux I__2757 (
            .O(N__22008),
            .I(N__22005));
    LocalMux I__2756 (
            .O(N__22005),
            .I(N__22002));
    Odrv4 I__2755 (
            .O(N__22002),
            .I(\nx.n3066 ));
    InMux I__2754 (
            .O(N__21999),
            .I(\nx.n10872 ));
    CascadeMux I__2753 (
            .O(N__21996),
            .I(N__21993));
    InMux I__2752 (
            .O(N__21993),
            .I(N__21990));
    LocalMux I__2751 (
            .O(N__21990),
            .I(N__21987));
    Odrv4 I__2750 (
            .O(N__21987),
            .I(\nx.n3065 ));
    InMux I__2749 (
            .O(N__21984),
            .I(\nx.n10873 ));
    CascadeMux I__2748 (
            .O(N__21981),
            .I(N__21978));
    InMux I__2747 (
            .O(N__21978),
            .I(N__21975));
    LocalMux I__2746 (
            .O(N__21975),
            .I(N__21972));
    Span4Mux_s3_h I__2745 (
            .O(N__21972),
            .I(N__21969));
    Odrv4 I__2744 (
            .O(N__21969),
            .I(\nx.n3064 ));
    InMux I__2743 (
            .O(N__21966),
            .I(\nx.n10874 ));
    InMux I__2742 (
            .O(N__21963),
            .I(N__21960));
    LocalMux I__2741 (
            .O(N__21960),
            .I(N__21957));
    Span4Mux_s1_h I__2740 (
            .O(N__21957),
            .I(N__21954));
    Span4Mux_v I__2739 (
            .O(N__21954),
            .I(N__21951));
    Odrv4 I__2738 (
            .O(N__21951),
            .I(\nx.n3063 ));
    InMux I__2737 (
            .O(N__21948),
            .I(\nx.n10875 ));
    InMux I__2736 (
            .O(N__21945),
            .I(\nx.n10876 ));
    InMux I__2735 (
            .O(N__21942),
            .I(N__21936));
    InMux I__2734 (
            .O(N__21941),
            .I(N__21936));
    LocalMux I__2733 (
            .O(N__21936),
            .I(neo_pixel_transmitter_t0_27));
    InMux I__2732 (
            .O(N__21933),
            .I(N__21930));
    LocalMux I__2731 (
            .O(N__21930),
            .I(\nx.n6 ));
    InMux I__2730 (
            .O(N__21927),
            .I(N__21924));
    LocalMux I__2729 (
            .O(N__21924),
            .I(N__21921));
    Odrv4 I__2728 (
            .O(N__21921),
            .I(\nx.n3077 ));
    InMux I__2727 (
            .O(N__21918),
            .I(bfn_3_26_0_));
    InMux I__2726 (
            .O(N__21915),
            .I(N__21912));
    LocalMux I__2725 (
            .O(N__21912),
            .I(\nx.n3076 ));
    InMux I__2724 (
            .O(N__21909),
            .I(\nx.n10862 ));
    CascadeMux I__2723 (
            .O(N__21906),
            .I(N__21902));
    InMux I__2722 (
            .O(N__21905),
            .I(N__21899));
    InMux I__2721 (
            .O(N__21902),
            .I(N__21896));
    LocalMux I__2720 (
            .O(N__21899),
            .I(N__21891));
    LocalMux I__2719 (
            .O(N__21896),
            .I(N__21891));
    Odrv4 I__2718 (
            .O(N__21891),
            .I(\nx.n3008 ));
    CascadeMux I__2717 (
            .O(N__21888),
            .I(N__21885));
    InMux I__2716 (
            .O(N__21885),
            .I(N__21882));
    LocalMux I__2715 (
            .O(N__21882),
            .I(\nx.n3075 ));
    InMux I__2714 (
            .O(N__21879),
            .I(\nx.n10863 ));
    CascadeMux I__2713 (
            .O(N__21876),
            .I(N__21873));
    InMux I__2712 (
            .O(N__21873),
            .I(N__21870));
    LocalMux I__2711 (
            .O(N__21870),
            .I(N__21866));
    InMux I__2710 (
            .O(N__21869),
            .I(N__21863));
    Span4Mux_h I__2709 (
            .O(N__21866),
            .I(N__21860));
    LocalMux I__2708 (
            .O(N__21863),
            .I(\nx.n3007 ));
    Odrv4 I__2707 (
            .O(N__21860),
            .I(\nx.n3007 ));
    InMux I__2706 (
            .O(N__21855),
            .I(N__21852));
    LocalMux I__2705 (
            .O(N__21852),
            .I(N__21849));
    Span4Mux_s2_h I__2704 (
            .O(N__21849),
            .I(N__21846));
    Odrv4 I__2703 (
            .O(N__21846),
            .I(\nx.n3074 ));
    InMux I__2702 (
            .O(N__21843),
            .I(\nx.n10864 ));
    CascadeMux I__2701 (
            .O(N__21840),
            .I(N__21837));
    InMux I__2700 (
            .O(N__21837),
            .I(N__21834));
    LocalMux I__2699 (
            .O(N__21834),
            .I(N__21831));
    Span4Mux_s2_h I__2698 (
            .O(N__21831),
            .I(N__21828));
    Odrv4 I__2697 (
            .O(N__21828),
            .I(\nx.n3073 ));
    InMux I__2696 (
            .O(N__21825),
            .I(\nx.n10865 ));
    InMux I__2695 (
            .O(N__21822),
            .I(N__21819));
    LocalMux I__2694 (
            .O(N__21819),
            .I(\nx.n3072 ));
    InMux I__2693 (
            .O(N__21816),
            .I(\nx.n10866 ));
    InMux I__2692 (
            .O(N__21813),
            .I(N__21810));
    LocalMux I__2691 (
            .O(N__21810),
            .I(N__21807));
    Odrv4 I__2690 (
            .O(N__21807),
            .I(\nx.n3071 ));
    InMux I__2689 (
            .O(N__21804),
            .I(\nx.n10867 ));
    InMux I__2688 (
            .O(N__21801),
            .I(N__21798));
    LocalMux I__2687 (
            .O(N__21798),
            .I(\nx.n12973 ));
    InMux I__2686 (
            .O(N__21795),
            .I(bfn_3_25_0_));
    InMux I__2685 (
            .O(N__21792),
            .I(N__21789));
    LocalMux I__2684 (
            .O(N__21789),
            .I(\nx.n12975 ));
    InMux I__2683 (
            .O(N__21786),
            .I(\nx.n10449 ));
    InMux I__2682 (
            .O(N__21783),
            .I(N__21780));
    LocalMux I__2681 (
            .O(N__21780),
            .I(\nx.n12977 ));
    InMux I__2680 (
            .O(N__21777),
            .I(\nx.n10450 ));
    InMux I__2679 (
            .O(N__21774),
            .I(N__21771));
    LocalMux I__2678 (
            .O(N__21771),
            .I(\nx.n12979 ));
    InMux I__2677 (
            .O(N__21768),
            .I(\nx.n10451 ));
    InMux I__2676 (
            .O(N__21765),
            .I(N__21761));
    InMux I__2675 (
            .O(N__21764),
            .I(N__21758));
    LocalMux I__2674 (
            .O(N__21761),
            .I(N__21754));
    LocalMux I__2673 (
            .O(N__21758),
            .I(N__21751));
    InMux I__2672 (
            .O(N__21757),
            .I(N__21748));
    Span4Mux_v I__2671 (
            .O(N__21754),
            .I(N__21743));
    Span4Mux_v I__2670 (
            .O(N__21751),
            .I(N__21743));
    LocalMux I__2669 (
            .O(N__21748),
            .I(timer_31));
    Odrv4 I__2668 (
            .O(N__21743),
            .I(timer_31));
    InMux I__2667 (
            .O(N__21738),
            .I(N__21735));
    LocalMux I__2666 (
            .O(N__21735),
            .I(N__21732));
    Span4Mux_v I__2665 (
            .O(N__21732),
            .I(N__21729));
    Span4Mux_v I__2664 (
            .O(N__21729),
            .I(N__21726));
    Odrv4 I__2663 (
            .O(N__21726),
            .I(\nx.n2 ));
    CascadeMux I__2662 (
            .O(N__21723),
            .I(N__21720));
    InMux I__2661 (
            .O(N__21720),
            .I(N__21717));
    LocalMux I__2660 (
            .O(N__21717),
            .I(\nx.n12981 ));
    InMux I__2659 (
            .O(N__21714),
            .I(\nx.n10452 ));
    InMux I__2658 (
            .O(N__21711),
            .I(N__21706));
    InMux I__2657 (
            .O(N__21710),
            .I(N__21703));
    InMux I__2656 (
            .O(N__21709),
            .I(N__21700));
    LocalMux I__2655 (
            .O(N__21706),
            .I(N__21697));
    LocalMux I__2654 (
            .O(N__21703),
            .I(N__21692));
    LocalMux I__2653 (
            .O(N__21700),
            .I(N__21692));
    Span4Mux_s3_h I__2652 (
            .O(N__21697),
            .I(N__21689));
    Span4Mux_s3_h I__2651 (
            .O(N__21692),
            .I(N__21686));
    Span4Mux_v I__2650 (
            .O(N__21689),
            .I(N__21683));
    Span4Mux_v I__2649 (
            .O(N__21686),
            .I(N__21680));
    Odrv4 I__2648 (
            .O(N__21683),
            .I(\nx.n7181 ));
    Odrv4 I__2647 (
            .O(N__21680),
            .I(\nx.n7181 ));
    CascadeMux I__2646 (
            .O(N__21675),
            .I(N__21671));
    InMux I__2645 (
            .O(N__21674),
            .I(N__21667));
    InMux I__2644 (
            .O(N__21671),
            .I(N__21664));
    InMux I__2643 (
            .O(N__21670),
            .I(N__21661));
    LocalMux I__2642 (
            .O(N__21667),
            .I(N__21656));
    LocalMux I__2641 (
            .O(N__21664),
            .I(N__21656));
    LocalMux I__2640 (
            .O(N__21661),
            .I(timer_27));
    Odrv12 I__2639 (
            .O(N__21656),
            .I(timer_27));
    InMux I__2638 (
            .O(N__21651),
            .I(N__21648));
    LocalMux I__2637 (
            .O(N__21648),
            .I(\nx.n12961 ));
    InMux I__2636 (
            .O(N__21645),
            .I(bfn_3_24_0_));
    InMux I__2635 (
            .O(N__21642),
            .I(N__21639));
    LocalMux I__2634 (
            .O(N__21639),
            .I(\nx.n12963 ));
    InMux I__2633 (
            .O(N__21636),
            .I(\nx.n10443 ));
    InMux I__2632 (
            .O(N__21633),
            .I(N__21630));
    LocalMux I__2631 (
            .O(N__21630),
            .I(\nx.n12965 ));
    InMux I__2630 (
            .O(N__21627),
            .I(N__21624));
    LocalMux I__2629 (
            .O(N__21624),
            .I(N__21621));
    Span4Mux_v I__2628 (
            .O(N__21621),
            .I(N__21618));
    Span4Mux_v I__2627 (
            .O(N__21618),
            .I(N__21615));
    Odrv4 I__2626 (
            .O(N__21615),
            .I(\nx.n10 ));
    CascadeMux I__2625 (
            .O(N__21612),
            .I(N__21608));
    InMux I__2624 (
            .O(N__21611),
            .I(N__21605));
    InMux I__2623 (
            .O(N__21608),
            .I(N__21602));
    LocalMux I__2622 (
            .O(N__21605),
            .I(N__21599));
    LocalMux I__2621 (
            .O(N__21602),
            .I(N__21595));
    Span4Mux_s2_h I__2620 (
            .O(N__21599),
            .I(N__21592));
    InMux I__2619 (
            .O(N__21598),
            .I(N__21589));
    Span4Mux_v I__2618 (
            .O(N__21595),
            .I(N__21586));
    Odrv4 I__2617 (
            .O(N__21592),
            .I(timer_23));
    LocalMux I__2616 (
            .O(N__21589),
            .I(timer_23));
    Odrv4 I__2615 (
            .O(N__21586),
            .I(timer_23));
    InMux I__2614 (
            .O(N__21579),
            .I(\nx.n10444 ));
    InMux I__2613 (
            .O(N__21576),
            .I(N__21573));
    LocalMux I__2612 (
            .O(N__21573),
            .I(N__21570));
    Odrv4 I__2611 (
            .O(N__21570),
            .I(\nx.n12967 ));
    InMux I__2610 (
            .O(N__21567),
            .I(N__21564));
    LocalMux I__2609 (
            .O(N__21564),
            .I(N__21561));
    Span4Mux_v I__2608 (
            .O(N__21561),
            .I(N__21558));
    Odrv4 I__2607 (
            .O(N__21558),
            .I(\nx.n9 ));
    InMux I__2606 (
            .O(N__21555),
            .I(N__21551));
    CascadeMux I__2605 (
            .O(N__21554),
            .I(N__21548));
    LocalMux I__2604 (
            .O(N__21551),
            .I(N__21544));
    InMux I__2603 (
            .O(N__21548),
            .I(N__21541));
    InMux I__2602 (
            .O(N__21547),
            .I(N__21538));
    Sp12to4 I__2601 (
            .O(N__21544),
            .I(N__21533));
    LocalMux I__2600 (
            .O(N__21541),
            .I(N__21533));
    LocalMux I__2599 (
            .O(N__21538),
            .I(timer_24));
    Odrv12 I__2598 (
            .O(N__21533),
            .I(timer_24));
    InMux I__2597 (
            .O(N__21528),
            .I(\nx.n10445 ));
    InMux I__2596 (
            .O(N__21525),
            .I(N__21522));
    LocalMux I__2595 (
            .O(N__21522),
            .I(N__21519));
    Odrv4 I__2594 (
            .O(N__21519),
            .I(\nx.n12969 ));
    InMux I__2593 (
            .O(N__21516),
            .I(\nx.n10446 ));
    InMux I__2592 (
            .O(N__21513),
            .I(N__21510));
    LocalMux I__2591 (
            .O(N__21510),
            .I(\nx.n12971 ));
    InMux I__2590 (
            .O(N__21507),
            .I(N__21504));
    LocalMux I__2589 (
            .O(N__21504),
            .I(N__21501));
    Span4Mux_v I__2588 (
            .O(N__21501),
            .I(N__21498));
    Span4Mux_h I__2587 (
            .O(N__21498),
            .I(N__21495));
    Odrv4 I__2586 (
            .O(N__21495),
            .I(\nx.n7_adj_597 ));
    CascadeMux I__2585 (
            .O(N__21492),
            .I(N__21488));
    InMux I__2584 (
            .O(N__21491),
            .I(N__21485));
    InMux I__2583 (
            .O(N__21488),
            .I(N__21482));
    LocalMux I__2582 (
            .O(N__21485),
            .I(N__21476));
    LocalMux I__2581 (
            .O(N__21482),
            .I(N__21476));
    InMux I__2580 (
            .O(N__21481),
            .I(N__21473));
    Span4Mux_v I__2579 (
            .O(N__21476),
            .I(N__21470));
    LocalMux I__2578 (
            .O(N__21473),
            .I(timer_26));
    Odrv4 I__2577 (
            .O(N__21470),
            .I(timer_26));
    InMux I__2576 (
            .O(N__21465),
            .I(\nx.n10447 ));
    InMux I__2575 (
            .O(N__21462),
            .I(N__21459));
    LocalMux I__2574 (
            .O(N__21459),
            .I(\nx.n12947 ));
    InMux I__2573 (
            .O(N__21456),
            .I(N__21453));
    LocalMux I__2572 (
            .O(N__21453),
            .I(N__21450));
    Odrv4 I__2571 (
            .O(N__21450),
            .I(\nx.n19_adj_622 ));
    CascadeMux I__2570 (
            .O(N__21447),
            .I(N__21444));
    InMux I__2569 (
            .O(N__21444),
            .I(N__21441));
    LocalMux I__2568 (
            .O(N__21441),
            .I(N__21436));
    InMux I__2567 (
            .O(N__21440),
            .I(N__21433));
    InMux I__2566 (
            .O(N__21439),
            .I(N__21430));
    Span4Mux_v I__2565 (
            .O(N__21436),
            .I(N__21427));
    LocalMux I__2564 (
            .O(N__21433),
            .I(timer_14));
    LocalMux I__2563 (
            .O(N__21430),
            .I(timer_14));
    Odrv4 I__2562 (
            .O(N__21427),
            .I(timer_14));
    InMux I__2561 (
            .O(N__21420),
            .I(\nx.n10435 ));
    InMux I__2560 (
            .O(N__21417),
            .I(N__21414));
    LocalMux I__2559 (
            .O(N__21414),
            .I(\nx.n12949 ));
    InMux I__2558 (
            .O(N__21411),
            .I(N__21408));
    LocalMux I__2557 (
            .O(N__21408),
            .I(N__21405));
    Span4Mux_v I__2556 (
            .O(N__21405),
            .I(N__21402));
    Odrv4 I__2555 (
            .O(N__21402),
            .I(\nx.n18_adj_623 ));
    InMux I__2554 (
            .O(N__21399),
            .I(N__21395));
    CascadeMux I__2553 (
            .O(N__21398),
            .I(N__21392));
    LocalMux I__2552 (
            .O(N__21395),
            .I(N__21389));
    InMux I__2551 (
            .O(N__21392),
            .I(N__21385));
    Span4Mux_v I__2550 (
            .O(N__21389),
            .I(N__21382));
    InMux I__2549 (
            .O(N__21388),
            .I(N__21379));
    LocalMux I__2548 (
            .O(N__21385),
            .I(N__21376));
    Odrv4 I__2547 (
            .O(N__21382),
            .I(timer_15));
    LocalMux I__2546 (
            .O(N__21379),
            .I(timer_15));
    Odrv12 I__2545 (
            .O(N__21376),
            .I(timer_15));
    InMux I__2544 (
            .O(N__21369),
            .I(bfn_3_23_0_));
    InMux I__2543 (
            .O(N__21366),
            .I(N__21363));
    LocalMux I__2542 (
            .O(N__21363),
            .I(\nx.n12951 ));
    InMux I__2541 (
            .O(N__21360),
            .I(N__21357));
    LocalMux I__2540 (
            .O(N__21357),
            .I(\nx.n17 ));
    InMux I__2539 (
            .O(N__21354),
            .I(N__21351));
    LocalMux I__2538 (
            .O(N__21351),
            .I(N__21347));
    CascadeMux I__2537 (
            .O(N__21350),
            .I(N__21344));
    Span4Mux_v I__2536 (
            .O(N__21347),
            .I(N__21341));
    InMux I__2535 (
            .O(N__21344),
            .I(N__21338));
    Span4Mux_v I__2534 (
            .O(N__21341),
            .I(N__21332));
    LocalMux I__2533 (
            .O(N__21338),
            .I(N__21332));
    InMux I__2532 (
            .O(N__21337),
            .I(N__21329));
    Span4Mux_v I__2531 (
            .O(N__21332),
            .I(N__21326));
    LocalMux I__2530 (
            .O(N__21329),
            .I(timer_16));
    Odrv4 I__2529 (
            .O(N__21326),
            .I(timer_16));
    InMux I__2528 (
            .O(N__21321),
            .I(\nx.n10437 ));
    InMux I__2527 (
            .O(N__21318),
            .I(N__21315));
    LocalMux I__2526 (
            .O(N__21315),
            .I(\nx.n12953 ));
    InMux I__2525 (
            .O(N__21312),
            .I(\nx.n10438 ));
    InMux I__2524 (
            .O(N__21309),
            .I(N__21306));
    LocalMux I__2523 (
            .O(N__21306),
            .I(\nx.n12955 ));
    InMux I__2522 (
            .O(N__21303),
            .I(\nx.n10439 ));
    InMux I__2521 (
            .O(N__21300),
            .I(N__21297));
    LocalMux I__2520 (
            .O(N__21297),
            .I(\nx.n12957 ));
    InMux I__2519 (
            .O(N__21294),
            .I(\nx.n10440 ));
    InMux I__2518 (
            .O(N__21291),
            .I(N__21288));
    LocalMux I__2517 (
            .O(N__21288),
            .I(\nx.n12959 ));
    InMux I__2516 (
            .O(N__21285),
            .I(\nx.n10441 ));
    InMux I__2515 (
            .O(N__21282),
            .I(N__21278));
    InMux I__2514 (
            .O(N__21281),
            .I(N__21274));
    LocalMux I__2513 (
            .O(N__21278),
            .I(N__21271));
    InMux I__2512 (
            .O(N__21277),
            .I(N__21268));
    LocalMux I__2511 (
            .O(N__21274),
            .I(N__21265));
    Odrv4 I__2510 (
            .O(N__21271),
            .I(timer_6));
    LocalMux I__2509 (
            .O(N__21268),
            .I(timer_6));
    Odrv12 I__2508 (
            .O(N__21265),
            .I(timer_6));
    CascadeMux I__2507 (
            .O(N__21258),
            .I(N__21255));
    InMux I__2506 (
            .O(N__21255),
            .I(N__21252));
    LocalMux I__2505 (
            .O(N__21252),
            .I(N__21249));
    Odrv4 I__2504 (
            .O(N__21249),
            .I(\nx.n27 ));
    InMux I__2503 (
            .O(N__21246),
            .I(N__21240));
    InMux I__2502 (
            .O(N__21245),
            .I(N__21240));
    LocalMux I__2501 (
            .O(N__21240),
            .I(N__21237));
    Span4Mux_s2_h I__2500 (
            .O(N__21237),
            .I(N__21234));
    Odrv4 I__2499 (
            .O(N__21234),
            .I(\nx.one_wire_N_528_6 ));
    InMux I__2498 (
            .O(N__21231),
            .I(\nx.n10427 ));
    InMux I__2497 (
            .O(N__21228),
            .I(N__21224));
    InMux I__2496 (
            .O(N__21227),
            .I(N__21221));
    LocalMux I__2495 (
            .O(N__21224),
            .I(N__21218));
    LocalMux I__2494 (
            .O(N__21221),
            .I(N__21213));
    Span4Mux_s2_h I__2493 (
            .O(N__21218),
            .I(N__21213));
    Odrv4 I__2492 (
            .O(N__21213),
            .I(\nx.one_wire_N_528_7 ));
    InMux I__2491 (
            .O(N__21210),
            .I(\nx.n10428 ));
    InMux I__2490 (
            .O(N__21207),
            .I(N__21204));
    LocalMux I__2489 (
            .O(N__21204),
            .I(N__21201));
    Odrv4 I__2488 (
            .O(N__21201),
            .I(\nx.n25 ));
    InMux I__2487 (
            .O(N__21198),
            .I(N__21194));
    CascadeMux I__2486 (
            .O(N__21197),
            .I(N__21191));
    LocalMux I__2485 (
            .O(N__21194),
            .I(N__21188));
    InMux I__2484 (
            .O(N__21191),
            .I(N__21184));
    Span4Mux_v I__2483 (
            .O(N__21188),
            .I(N__21181));
    InMux I__2482 (
            .O(N__21187),
            .I(N__21178));
    LocalMux I__2481 (
            .O(N__21184),
            .I(N__21175));
    Odrv4 I__2480 (
            .O(N__21181),
            .I(timer_8));
    LocalMux I__2479 (
            .O(N__21178),
            .I(timer_8));
    Odrv12 I__2478 (
            .O(N__21175),
            .I(timer_8));
    InMux I__2477 (
            .O(N__21168),
            .I(N__21163));
    InMux I__2476 (
            .O(N__21167),
            .I(N__21160));
    InMux I__2475 (
            .O(N__21166),
            .I(N__21157));
    LocalMux I__2474 (
            .O(N__21163),
            .I(N__21152));
    LocalMux I__2473 (
            .O(N__21160),
            .I(N__21152));
    LocalMux I__2472 (
            .O(N__21157),
            .I(N__21149));
    Span4Mux_v I__2471 (
            .O(N__21152),
            .I(N__21146));
    Span4Mux_s3_h I__2470 (
            .O(N__21149),
            .I(N__21143));
    Odrv4 I__2469 (
            .O(N__21146),
            .I(\nx.one_wire_N_528_8 ));
    Odrv4 I__2468 (
            .O(N__21143),
            .I(\nx.one_wire_N_528_8 ));
    InMux I__2467 (
            .O(N__21138),
            .I(bfn_3_22_0_));
    CascadeMux I__2466 (
            .O(N__21135),
            .I(N__21131));
    CascadeMux I__2465 (
            .O(N__21134),
            .I(N__21127));
    InMux I__2464 (
            .O(N__21131),
            .I(N__21124));
    InMux I__2463 (
            .O(N__21130),
            .I(N__21121));
    InMux I__2462 (
            .O(N__21127),
            .I(N__21118));
    LocalMux I__2461 (
            .O(N__21124),
            .I(N__21115));
    LocalMux I__2460 (
            .O(N__21121),
            .I(N__21110));
    LocalMux I__2459 (
            .O(N__21118),
            .I(N__21110));
    Span4Mux_s2_h I__2458 (
            .O(N__21115),
            .I(N__21107));
    Span4Mux_s2_h I__2457 (
            .O(N__21110),
            .I(N__21104));
    Odrv4 I__2456 (
            .O(N__21107),
            .I(\nx.one_wire_N_528_9 ));
    Odrv4 I__2455 (
            .O(N__21104),
            .I(\nx.one_wire_N_528_9 ));
    InMux I__2454 (
            .O(N__21099),
            .I(\nx.n10430 ));
    InMux I__2453 (
            .O(N__21096),
            .I(N__21092));
    CascadeMux I__2452 (
            .O(N__21095),
            .I(N__21089));
    LocalMux I__2451 (
            .O(N__21092),
            .I(N__21086));
    InMux I__2450 (
            .O(N__21089),
            .I(N__21083));
    Span4Mux_v I__2449 (
            .O(N__21086),
            .I(N__21077));
    LocalMux I__2448 (
            .O(N__21083),
            .I(N__21077));
    InMux I__2447 (
            .O(N__21082),
            .I(N__21074));
    Span4Mux_v I__2446 (
            .O(N__21077),
            .I(N__21071));
    LocalMux I__2445 (
            .O(N__21074),
            .I(timer_10));
    Odrv4 I__2444 (
            .O(N__21071),
            .I(timer_10));
    InMux I__2443 (
            .O(N__21066),
            .I(N__21061));
    InMux I__2442 (
            .O(N__21065),
            .I(N__21058));
    InMux I__2441 (
            .O(N__21064),
            .I(N__21055));
    LocalMux I__2440 (
            .O(N__21061),
            .I(N__21052));
    LocalMux I__2439 (
            .O(N__21058),
            .I(N__21049));
    LocalMux I__2438 (
            .O(N__21055),
            .I(N__21046));
    Span12Mux_s2_h I__2437 (
            .O(N__21052),
            .I(N__21043));
    Span4Mux_v I__2436 (
            .O(N__21049),
            .I(N__21038));
    Span4Mux_s2_h I__2435 (
            .O(N__21046),
            .I(N__21038));
    Odrv12 I__2434 (
            .O(N__21043),
            .I(\nx.one_wire_N_528_10 ));
    Odrv4 I__2433 (
            .O(N__21038),
            .I(\nx.one_wire_N_528_10 ));
    InMux I__2432 (
            .O(N__21033),
            .I(\nx.n10431 ));
    InMux I__2431 (
            .O(N__21030),
            .I(\nx.n10432 ));
    InMux I__2430 (
            .O(N__21027),
            .I(N__21024));
    LocalMux I__2429 (
            .O(N__21024),
            .I(\nx.one_wire_N_528_11 ));
    InMux I__2428 (
            .O(N__21021),
            .I(N__21017));
    InMux I__2427 (
            .O(N__21020),
            .I(N__21013));
    LocalMux I__2426 (
            .O(N__21017),
            .I(N__21010));
    InMux I__2425 (
            .O(N__21016),
            .I(N__21007));
    LocalMux I__2424 (
            .O(N__21013),
            .I(N__21004));
    Odrv4 I__2423 (
            .O(N__21010),
            .I(timer_12));
    LocalMux I__2422 (
            .O(N__21007),
            .I(timer_12));
    Odrv12 I__2421 (
            .O(N__21004),
            .I(timer_12));
    CascadeMux I__2420 (
            .O(N__20997),
            .I(N__20994));
    InMux I__2419 (
            .O(N__20994),
            .I(N__20991));
    LocalMux I__2418 (
            .O(N__20991),
            .I(N__20988));
    Span4Mux_v I__2417 (
            .O(N__20988),
            .I(N__20985));
    Span4Mux_s2_h I__2416 (
            .O(N__20985),
            .I(N__20982));
    Odrv4 I__2415 (
            .O(N__20982),
            .I(\nx.n21_adj_620 ));
    InMux I__2414 (
            .O(N__20979),
            .I(\nx.n10433 ));
    InMux I__2413 (
            .O(N__20976),
            .I(N__20973));
    LocalMux I__2412 (
            .O(N__20973),
            .I(\nx.n12945 ));
    InMux I__2411 (
            .O(N__20970),
            .I(\nx.n10434 ));
    InMux I__2410 (
            .O(N__20967),
            .I(\nx.n10508 ));
    InMux I__2409 (
            .O(N__20964),
            .I(\nx.n10509 ));
    InMux I__2408 (
            .O(N__20961),
            .I(N__20958));
    LocalMux I__2407 (
            .O(N__20958),
            .I(N__20955));
    Odrv12 I__2406 (
            .O(N__20955),
            .I(\nx.n32_adj_651 ));
    CascadeMux I__2405 (
            .O(N__20952),
            .I(N__20948));
    InMux I__2404 (
            .O(N__20951),
            .I(N__20944));
    InMux I__2403 (
            .O(N__20948),
            .I(N__20941));
    InMux I__2402 (
            .O(N__20947),
            .I(N__20938));
    LocalMux I__2401 (
            .O(N__20944),
            .I(N__20933));
    LocalMux I__2400 (
            .O(N__20941),
            .I(N__20933));
    LocalMux I__2399 (
            .O(N__20938),
            .I(timer_1));
    Odrv12 I__2398 (
            .O(N__20933),
            .I(timer_1));
    InMux I__2397 (
            .O(N__20928),
            .I(N__20925));
    LocalMux I__2396 (
            .O(N__20925),
            .I(N__20921));
    InMux I__2395 (
            .O(N__20924),
            .I(N__20918));
    Span4Mux_s2_h I__2394 (
            .O(N__20921),
            .I(N__20915));
    LocalMux I__2393 (
            .O(N__20918),
            .I(\nx.n11533 ));
    Odrv4 I__2392 (
            .O(N__20915),
            .I(\nx.n11533 ));
    InMux I__2391 (
            .O(N__20910),
            .I(\nx.n10422 ));
    InMux I__2390 (
            .O(N__20907),
            .I(N__20902));
    InMux I__2389 (
            .O(N__20906),
            .I(N__20899));
    InMux I__2388 (
            .O(N__20905),
            .I(N__20896));
    LocalMux I__2387 (
            .O(N__20902),
            .I(N__20893));
    LocalMux I__2386 (
            .O(N__20899),
            .I(\nx.one_wire_N_528_2 ));
    LocalMux I__2385 (
            .O(N__20896),
            .I(\nx.one_wire_N_528_2 ));
    Odrv4 I__2384 (
            .O(N__20893),
            .I(\nx.one_wire_N_528_2 ));
    InMux I__2383 (
            .O(N__20886),
            .I(\nx.n10423 ));
    InMux I__2382 (
            .O(N__20883),
            .I(N__20880));
    LocalMux I__2381 (
            .O(N__20880),
            .I(\nx.n30_adj_598 ));
    CascadeMux I__2380 (
            .O(N__20877),
            .I(N__20873));
    InMux I__2379 (
            .O(N__20876),
            .I(N__20870));
    InMux I__2378 (
            .O(N__20873),
            .I(N__20866));
    LocalMux I__2377 (
            .O(N__20870),
            .I(N__20863));
    InMux I__2376 (
            .O(N__20869),
            .I(N__20860));
    LocalMux I__2375 (
            .O(N__20866),
            .I(N__20857));
    Odrv4 I__2374 (
            .O(N__20863),
            .I(timer_3));
    LocalMux I__2373 (
            .O(N__20860),
            .I(timer_3));
    Odrv12 I__2372 (
            .O(N__20857),
            .I(timer_3));
    InMux I__2371 (
            .O(N__20850),
            .I(N__20845));
    InMux I__2370 (
            .O(N__20849),
            .I(N__20842));
    InMux I__2369 (
            .O(N__20848),
            .I(N__20839));
    LocalMux I__2368 (
            .O(N__20845),
            .I(N__20836));
    LocalMux I__2367 (
            .O(N__20842),
            .I(\nx.one_wire_N_528_3 ));
    LocalMux I__2366 (
            .O(N__20839),
            .I(\nx.one_wire_N_528_3 ));
    Odrv4 I__2365 (
            .O(N__20836),
            .I(\nx.one_wire_N_528_3 ));
    InMux I__2364 (
            .O(N__20829),
            .I(\nx.n10424 ));
    InMux I__2363 (
            .O(N__20826),
            .I(N__20823));
    LocalMux I__2362 (
            .O(N__20823),
            .I(N__20820));
    Odrv12 I__2361 (
            .O(N__20820),
            .I(\nx.n29 ));
    InMux I__2360 (
            .O(N__20817),
            .I(N__20813));
    CascadeMux I__2359 (
            .O(N__20816),
            .I(N__20810));
    LocalMux I__2358 (
            .O(N__20813),
            .I(N__20807));
    InMux I__2357 (
            .O(N__20810),
            .I(N__20804));
    Span4Mux_v I__2356 (
            .O(N__20807),
            .I(N__20798));
    LocalMux I__2355 (
            .O(N__20804),
            .I(N__20798));
    InMux I__2354 (
            .O(N__20803),
            .I(N__20795));
    Span4Mux_v I__2353 (
            .O(N__20798),
            .I(N__20792));
    LocalMux I__2352 (
            .O(N__20795),
            .I(timer_4));
    Odrv4 I__2351 (
            .O(N__20792),
            .I(timer_4));
    InMux I__2350 (
            .O(N__20787),
            .I(N__20781));
    InMux I__2349 (
            .O(N__20786),
            .I(N__20781));
    LocalMux I__2348 (
            .O(N__20781),
            .I(N__20778));
    Odrv4 I__2347 (
            .O(N__20778),
            .I(\nx.one_wire_N_528_4 ));
    InMux I__2346 (
            .O(N__20775),
            .I(\nx.n10425 ));
    InMux I__2345 (
            .O(N__20772),
            .I(N__20768));
    InMux I__2344 (
            .O(N__20771),
            .I(N__20765));
    LocalMux I__2343 (
            .O(N__20768),
            .I(N__20762));
    LocalMux I__2342 (
            .O(N__20765),
            .I(N__20758));
    Span12Mux_s2_h I__2341 (
            .O(N__20762),
            .I(N__20755));
    InMux I__2340 (
            .O(N__20761),
            .I(N__20752));
    Span4Mux_v I__2339 (
            .O(N__20758),
            .I(N__20749));
    Odrv12 I__2338 (
            .O(N__20755),
            .I(timer_5));
    LocalMux I__2337 (
            .O(N__20752),
            .I(timer_5));
    Odrv4 I__2336 (
            .O(N__20749),
            .I(timer_5));
    CascadeMux I__2335 (
            .O(N__20742),
            .I(N__20739));
    InMux I__2334 (
            .O(N__20739),
            .I(N__20736));
    LocalMux I__2333 (
            .O(N__20736),
            .I(\nx.n28 ));
    InMux I__2332 (
            .O(N__20733),
            .I(N__20730));
    LocalMux I__2331 (
            .O(N__20730),
            .I(N__20726));
    InMux I__2330 (
            .O(N__20729),
            .I(N__20723));
    Span12Mux_v I__2329 (
            .O(N__20726),
            .I(N__20720));
    LocalMux I__2328 (
            .O(N__20723),
            .I(N__20717));
    Odrv12 I__2327 (
            .O(N__20720),
            .I(\nx.one_wire_N_528_5 ));
    Odrv4 I__2326 (
            .O(N__20717),
            .I(\nx.one_wire_N_528_5 ));
    InMux I__2325 (
            .O(N__20712),
            .I(\nx.n10426 ));
    InMux I__2324 (
            .O(N__20709),
            .I(\nx.n10499 ));
    InMux I__2323 (
            .O(N__20706),
            .I(\nx.n10500 ));
    InMux I__2322 (
            .O(N__20703),
            .I(\nx.n10501 ));
    InMux I__2321 (
            .O(N__20700),
            .I(bfn_3_20_0_));
    InMux I__2320 (
            .O(N__20697),
            .I(\nx.n10503 ));
    InMux I__2319 (
            .O(N__20694),
            .I(\nx.n10504 ));
    InMux I__2318 (
            .O(N__20691),
            .I(\nx.n10505 ));
    InMux I__2317 (
            .O(N__20688),
            .I(\nx.n10506 ));
    InMux I__2316 (
            .O(N__20685),
            .I(\nx.n10507 ));
    InMux I__2315 (
            .O(N__20682),
            .I(\nx.n10490 ));
    InMux I__2314 (
            .O(N__20679),
            .I(\nx.n10491 ));
    InMux I__2313 (
            .O(N__20676),
            .I(\nx.n10492 ));
    InMux I__2312 (
            .O(N__20673),
            .I(\nx.n10493 ));
    InMux I__2311 (
            .O(N__20670),
            .I(bfn_3_19_0_));
    InMux I__2310 (
            .O(N__20667),
            .I(\nx.n10495 ));
    InMux I__2309 (
            .O(N__20664),
            .I(\nx.n10496 ));
    InMux I__2308 (
            .O(N__20661),
            .I(\nx.n10497 ));
    InMux I__2307 (
            .O(N__20658),
            .I(\nx.n10498 ));
    InMux I__2306 (
            .O(N__20655),
            .I(\nx.n10480 ));
    InMux I__2305 (
            .O(N__20652),
            .I(\nx.n10481 ));
    InMux I__2304 (
            .O(N__20649),
            .I(\nx.n10482 ));
    InMux I__2303 (
            .O(N__20646),
            .I(\nx.n10483 ));
    InMux I__2302 (
            .O(N__20643),
            .I(\nx.n10484 ));
    InMux I__2301 (
            .O(N__20640),
            .I(\nx.n10485 ));
    InMux I__2300 (
            .O(N__20637),
            .I(bfn_3_18_0_));
    InMux I__2299 (
            .O(N__20634),
            .I(\nx.n10487 ));
    InMux I__2298 (
            .O(N__20631),
            .I(\nx.n10488 ));
    InMux I__2297 (
            .O(N__20628),
            .I(\nx.n10489 ));
    CascadeMux I__2296 (
            .O(N__20625),
            .I(N__20621));
    InMux I__2295 (
            .O(N__20624),
            .I(N__20616));
    InMux I__2294 (
            .O(N__20621),
            .I(N__20616));
    LocalMux I__2293 (
            .O(N__20616),
            .I(\nx.n1302 ));
    CascadeMux I__2292 (
            .O(N__20613),
            .I(N__20610));
    InMux I__2291 (
            .O(N__20610),
            .I(N__20607));
    LocalMux I__2290 (
            .O(N__20607),
            .I(\nx.n1369 ));
    InMux I__2289 (
            .O(N__20604),
            .I(N__20598));
    InMux I__2288 (
            .O(N__20603),
            .I(N__20598));
    LocalMux I__2287 (
            .O(N__20598),
            .I(neo_pixel_transmitter_t0_1));
    InMux I__2286 (
            .O(N__20595),
            .I(N__20591));
    InMux I__2285 (
            .O(N__20594),
            .I(N__20588));
    LocalMux I__2284 (
            .O(N__20591),
            .I(neo_pixel_transmitter_t0_31));
    LocalMux I__2283 (
            .O(N__20588),
            .I(neo_pixel_transmitter_t0_31));
    InMux I__2282 (
            .O(N__20583),
            .I(N__20579));
    InMux I__2281 (
            .O(N__20582),
            .I(N__20576));
    LocalMux I__2280 (
            .O(N__20579),
            .I(neo_pixel_transmitter_t0_4));
    LocalMux I__2279 (
            .O(N__20576),
            .I(neo_pixel_transmitter_t0_4));
    InMux I__2278 (
            .O(N__20571),
            .I(bfn_3_17_0_));
    InMux I__2277 (
            .O(N__20568),
            .I(\nx.n10479 ));
    InMux I__2276 (
            .O(N__20565),
            .I(\nx.n10573 ));
    InMux I__2275 (
            .O(N__20562),
            .I(\nx.n10574 ));
    InMux I__2274 (
            .O(N__20559),
            .I(\nx.n10575 ));
    InMux I__2273 (
            .O(N__20556),
            .I(\nx.n10576 ));
    InMux I__2272 (
            .O(N__20553),
            .I(\nx.n10577 ));
    InMux I__2271 (
            .O(N__20550),
            .I(\nx.n10578 ));
    InMux I__2270 (
            .O(N__20547),
            .I(\nx.n10579 ));
    InMux I__2269 (
            .O(N__20544),
            .I(bfn_2_32_0_));
    CascadeMux I__2268 (
            .O(N__20541),
            .I(N__20538));
    InMux I__2267 (
            .O(N__20538),
            .I(N__20534));
    InMux I__2266 (
            .O(N__20537),
            .I(N__20531));
    LocalMux I__2265 (
            .O(N__20534),
            .I(\nx.n1301 ));
    LocalMux I__2264 (
            .O(N__20531),
            .I(\nx.n1301 ));
    InMux I__2263 (
            .O(N__20526),
            .I(\nx.n10581 ));
    InMux I__2262 (
            .O(N__20523),
            .I(N__20520));
    LocalMux I__2261 (
            .O(N__20520),
            .I(\nx.n1172 ));
    CascadeMux I__2260 (
            .O(N__20517),
            .I(N__20514));
    InMux I__2259 (
            .O(N__20514),
            .I(N__20510));
    InMux I__2258 (
            .O(N__20513),
            .I(N__20507));
    LocalMux I__2257 (
            .O(N__20510),
            .I(\nx.n1204 ));
    LocalMux I__2256 (
            .O(N__20507),
            .I(\nx.n1204 ));
    InMux I__2255 (
            .O(N__20502),
            .I(N__20499));
    LocalMux I__2254 (
            .O(N__20499),
            .I(\nx.n1271 ));
    CascadeMux I__2253 (
            .O(N__20496),
            .I(\nx.n1204_cascade_ ));
    InMux I__2252 (
            .O(N__20493),
            .I(N__20490));
    LocalMux I__2251 (
            .O(N__20490),
            .I(\nx.n11_adj_624 ));
    CascadeMux I__2250 (
            .O(N__20487),
            .I(N__20484));
    InMux I__2249 (
            .O(N__20484),
            .I(N__20481));
    LocalMux I__2248 (
            .O(N__20481),
            .I(\nx.n13 ));
    InMux I__2247 (
            .O(N__20478),
            .I(N__20474));
    CascadeMux I__2246 (
            .O(N__20477),
            .I(N__20471));
    LocalMux I__2245 (
            .O(N__20474),
            .I(N__20468));
    InMux I__2244 (
            .O(N__20471),
            .I(N__20465));
    Span4Mux_h I__2243 (
            .O(N__20468),
            .I(N__20462));
    LocalMux I__2242 (
            .O(N__20465),
            .I(\nx.n1206 ));
    Odrv4 I__2241 (
            .O(N__20462),
            .I(\nx.n1206 ));
    InMux I__2240 (
            .O(N__20457),
            .I(N__20454));
    LocalMux I__2239 (
            .O(N__20454),
            .I(\nx.n1275 ));
    CascadeMux I__2238 (
            .O(N__20451),
            .I(\nx.n1235_cascade_ ));
    CascadeMux I__2237 (
            .O(N__20448),
            .I(N__20444));
    InMux I__2236 (
            .O(N__20447),
            .I(N__20441));
    InMux I__2235 (
            .O(N__20444),
            .I(N__20438));
    LocalMux I__2234 (
            .O(N__20441),
            .I(\nx.n1208 ));
    LocalMux I__2233 (
            .O(N__20438),
            .I(\nx.n1208 ));
    InMux I__2232 (
            .O(N__20433),
            .I(N__20430));
    LocalMux I__2231 (
            .O(N__20430),
            .I(\nx.n1175 ));
    InMux I__2230 (
            .O(N__20427),
            .I(N__20420));
    CascadeMux I__2229 (
            .O(N__20426),
            .I(N__20416));
    CascadeMux I__2228 (
            .O(N__20425),
            .I(N__20413));
    InMux I__2227 (
            .O(N__20424),
            .I(N__20407));
    InMux I__2226 (
            .O(N__20423),
            .I(N__20407));
    LocalMux I__2225 (
            .O(N__20420),
            .I(N__20404));
    InMux I__2224 (
            .O(N__20419),
            .I(N__20401));
    InMux I__2223 (
            .O(N__20416),
            .I(N__20394));
    InMux I__2222 (
            .O(N__20413),
            .I(N__20394));
    InMux I__2221 (
            .O(N__20412),
            .I(N__20394));
    LocalMux I__2220 (
            .O(N__20407),
            .I(\nx.n1136 ));
    Odrv4 I__2219 (
            .O(N__20404),
            .I(\nx.n1136 ));
    LocalMux I__2218 (
            .O(N__20401),
            .I(\nx.n1136 ));
    LocalMux I__2217 (
            .O(N__20394),
            .I(\nx.n1136 ));
    CascadeMux I__2216 (
            .O(N__20385),
            .I(N__20382));
    InMux I__2215 (
            .O(N__20382),
            .I(N__20378));
    InMux I__2214 (
            .O(N__20381),
            .I(N__20375));
    LocalMux I__2213 (
            .O(N__20378),
            .I(\nx.n1207 ));
    LocalMux I__2212 (
            .O(N__20375),
            .I(\nx.n1207 ));
    InMux I__2211 (
            .O(N__20370),
            .I(N__20367));
    LocalMux I__2210 (
            .O(N__20367),
            .I(\nx.n1274 ));
    CascadeMux I__2209 (
            .O(N__20364),
            .I(\nx.n1207_cascade_ ));
    CascadeMux I__2208 (
            .O(N__20361),
            .I(\nx.n1306_cascade_ ));
    InMux I__2207 (
            .O(N__20358),
            .I(N__20355));
    LocalMux I__2206 (
            .O(N__20355),
            .I(N__20352));
    Odrv4 I__2205 (
            .O(N__20352),
            .I(\nx.n10_adj_626 ));
    InMux I__2204 (
            .O(N__20349),
            .I(bfn_2_31_0_));
    InMux I__2203 (
            .O(N__20346),
            .I(N__20343));
    LocalMux I__2202 (
            .O(N__20343),
            .I(\nx.n1177 ));
    InMux I__2201 (
            .O(N__20340),
            .I(bfn_2_29_0_));
    CascadeMux I__2200 (
            .O(N__20337),
            .I(N__20332));
    InMux I__2199 (
            .O(N__20336),
            .I(N__20327));
    InMux I__2198 (
            .O(N__20335),
            .I(N__20327));
    InMux I__2197 (
            .O(N__20332),
            .I(N__20324));
    LocalMux I__2196 (
            .O(N__20327),
            .I(\nx.n1109 ));
    LocalMux I__2195 (
            .O(N__20324),
            .I(\nx.n1109 ));
    CascadeMux I__2194 (
            .O(N__20319),
            .I(N__20316));
    InMux I__2193 (
            .O(N__20316),
            .I(N__20313));
    LocalMux I__2192 (
            .O(N__20313),
            .I(N__20310));
    Odrv4 I__2191 (
            .O(N__20310),
            .I(\nx.n1176 ));
    InMux I__2190 (
            .O(N__20307),
            .I(\nx.n10461 ));
    InMux I__2189 (
            .O(N__20304),
            .I(\nx.n10462 ));
    InMux I__2188 (
            .O(N__20301),
            .I(N__20298));
    LocalMux I__2187 (
            .O(N__20298),
            .I(N__20295));
    Odrv4 I__2186 (
            .O(N__20295),
            .I(\nx.n1174 ));
    InMux I__2185 (
            .O(N__20292),
            .I(\nx.n10463 ));
    InMux I__2184 (
            .O(N__20289),
            .I(\nx.n10464 ));
    InMux I__2183 (
            .O(N__20286),
            .I(\nx.n10465 ));
    CascadeMux I__2182 (
            .O(N__20283),
            .I(N__20280));
    InMux I__2181 (
            .O(N__20280),
            .I(N__20277));
    LocalMux I__2180 (
            .O(N__20277),
            .I(\nx.n1171 ));
    InMux I__2179 (
            .O(N__20274),
            .I(\nx.n10466 ));
    InMux I__2178 (
            .O(N__20271),
            .I(\nx.n10467 ));
    InMux I__2177 (
            .O(N__20268),
            .I(N__20265));
    LocalMux I__2176 (
            .O(N__20265),
            .I(N__20262));
    Span4Mux_s1_v I__2175 (
            .O(N__20262),
            .I(N__20258));
    InMux I__2174 (
            .O(N__20261),
            .I(N__20255));
    Odrv4 I__2173 (
            .O(N__20258),
            .I(\nx.n1202 ));
    LocalMux I__2172 (
            .O(N__20255),
            .I(\nx.n1202 ));
    CascadeMux I__2171 (
            .O(N__20250),
            .I(N__20247));
    InMux I__2170 (
            .O(N__20247),
            .I(N__20244));
    LocalMux I__2169 (
            .O(N__20244),
            .I(\nx.n1173 ));
    InMux I__2168 (
            .O(N__20241),
            .I(N__20238));
    LocalMux I__2167 (
            .O(N__20238),
            .I(N__20235));
    Odrv4 I__2166 (
            .O(N__20235),
            .I(\nx.n3151 ));
    InMux I__2165 (
            .O(N__20232),
            .I(N__20229));
    LocalMux I__2164 (
            .O(N__20229),
            .I(N__20226));
    Odrv12 I__2163 (
            .O(N__20226),
            .I(\nx.n61 ));
    CascadeMux I__2162 (
            .O(N__20223),
            .I(N__20218));
    InMux I__2161 (
            .O(N__20222),
            .I(N__20215));
    InMux I__2160 (
            .O(N__20221),
            .I(N__20212));
    InMux I__2159 (
            .O(N__20218),
            .I(N__20209));
    LocalMux I__2158 (
            .O(N__20215),
            .I(N__20204));
    LocalMux I__2157 (
            .O(N__20212),
            .I(N__20204));
    LocalMux I__2156 (
            .O(N__20209),
            .I(\nx.n3099 ));
    Odrv4 I__2155 (
            .O(N__20204),
            .I(\nx.n3099 ));
    InMux I__2154 (
            .O(N__20199),
            .I(N__20196));
    LocalMux I__2153 (
            .O(N__20196),
            .I(N__20193));
    Span4Mux_v I__2152 (
            .O(N__20193),
            .I(N__20190));
    Odrv4 I__2151 (
            .O(N__20190),
            .I(neopxl_color_prev_7));
    InMux I__2150 (
            .O(N__20187),
            .I(N__20184));
    LocalMux I__2149 (
            .O(N__20184),
            .I(\nx.n54 ));
    CascadeMux I__2148 (
            .O(N__20181),
            .I(\nx.n43_adj_709_cascade_ ));
    InMux I__2147 (
            .O(N__20178),
            .I(N__20175));
    LocalMux I__2146 (
            .O(N__20175),
            .I(\nx.n49_adj_710 ));
    InMux I__2145 (
            .O(N__20172),
            .I(N__20168));
    InMux I__2144 (
            .O(N__20171),
            .I(N__20165));
    LocalMux I__2143 (
            .O(N__20168),
            .I(N__20158));
    LocalMux I__2142 (
            .O(N__20165),
            .I(N__20158));
    InMux I__2141 (
            .O(N__20164),
            .I(N__20153));
    InMux I__2140 (
            .O(N__20163),
            .I(N__20153));
    Span4Mux_v I__2139 (
            .O(N__20158),
            .I(N__20148));
    LocalMux I__2138 (
            .O(N__20153),
            .I(N__20148));
    Span4Mux_v I__2137 (
            .O(N__20148),
            .I(N__20145));
    Odrv4 I__2136 (
            .O(N__20145),
            .I(state_3_N_377_1));
    InMux I__2135 (
            .O(N__20142),
            .I(N__20139));
    LocalMux I__2134 (
            .O(N__20139),
            .I(N__20134));
    InMux I__2133 (
            .O(N__20138),
            .I(N__20131));
    InMux I__2132 (
            .O(N__20137),
            .I(N__20128));
    Span4Mux_s1_h I__2131 (
            .O(N__20134),
            .I(N__20125));
    LocalMux I__2130 (
            .O(N__20131),
            .I(\nx.n3084 ));
    LocalMux I__2129 (
            .O(N__20128),
            .I(\nx.n3084 ));
    Odrv4 I__2128 (
            .O(N__20125),
            .I(\nx.n3084 ));
    InMux I__2127 (
            .O(N__20118),
            .I(N__20115));
    LocalMux I__2126 (
            .O(N__20115),
            .I(\nx.n3174 ));
    InMux I__2125 (
            .O(N__20112),
            .I(N__20109));
    LocalMux I__2124 (
            .O(N__20109),
            .I(\nx.n23_adj_700 ));
    CascadeMux I__2123 (
            .O(N__20106),
            .I(N__20103));
    InMux I__2122 (
            .O(N__20103),
            .I(N__20098));
    InMux I__2121 (
            .O(N__20102),
            .I(N__20095));
    InMux I__2120 (
            .O(N__20101),
            .I(N__20092));
    LocalMux I__2119 (
            .O(N__20098),
            .I(\nx.n3107 ));
    LocalMux I__2118 (
            .O(N__20095),
            .I(\nx.n3107 ));
    LocalMux I__2117 (
            .O(N__20092),
            .I(\nx.n3107 ));
    InMux I__2116 (
            .O(N__20085),
            .I(N__20082));
    LocalMux I__2115 (
            .O(N__20082),
            .I(\nx.n3162 ));
    CascadeMux I__2114 (
            .O(N__20079),
            .I(\nx.n12327_cascade_ ));
    InMux I__2113 (
            .O(N__20076),
            .I(N__20072));
    CascadeMux I__2112 (
            .O(N__20075),
            .I(N__20069));
    LocalMux I__2111 (
            .O(N__20072),
            .I(N__20066));
    InMux I__2110 (
            .O(N__20069),
            .I(N__20063));
    Span4Mux_v I__2109 (
            .O(N__20066),
            .I(N__20059));
    LocalMux I__2108 (
            .O(N__20063),
            .I(N__20056));
    InMux I__2107 (
            .O(N__20062),
            .I(N__20053));
    Odrv4 I__2106 (
            .O(N__20059),
            .I(\nx.n3095 ));
    Odrv12 I__2105 (
            .O(N__20056),
            .I(\nx.n3095 ));
    LocalMux I__2104 (
            .O(N__20053),
            .I(\nx.n3095 ));
    CascadeMux I__2103 (
            .O(N__20046),
            .I(N__20043));
    InMux I__2102 (
            .O(N__20043),
            .I(N__20040));
    LocalMux I__2101 (
            .O(N__20040),
            .I(\nx.n3166 ));
    InMux I__2100 (
            .O(N__20037),
            .I(N__20034));
    LocalMux I__2099 (
            .O(N__20034),
            .I(\nx.n3177 ));
    InMux I__2098 (
            .O(N__20031),
            .I(N__20028));
    LocalMux I__2097 (
            .O(N__20028),
            .I(N__20024));
    InMux I__2096 (
            .O(N__20027),
            .I(N__20021));
    Odrv12 I__2095 (
            .O(N__20024),
            .I(\nx.n3209 ));
    LocalMux I__2094 (
            .O(N__20021),
            .I(\nx.n3209 ));
    InMux I__2093 (
            .O(N__20016),
            .I(N__20013));
    LocalMux I__2092 (
            .O(N__20013),
            .I(\nx.n3171 ));
    InMux I__2091 (
            .O(N__20010),
            .I(N__20007));
    LocalMux I__2090 (
            .O(N__20007),
            .I(\nx.n3175 ));
    InMux I__2089 (
            .O(N__20004),
            .I(N__19999));
    CascadeMux I__2088 (
            .O(N__20003),
            .I(N__19996));
    InMux I__2087 (
            .O(N__20002),
            .I(N__19993));
    LocalMux I__2086 (
            .O(N__19999),
            .I(N__19990));
    InMux I__2085 (
            .O(N__19996),
            .I(N__19987));
    LocalMux I__2084 (
            .O(N__19993),
            .I(\nx.n3108 ));
    Odrv4 I__2083 (
            .O(N__19990),
            .I(\nx.n3108 ));
    LocalMux I__2082 (
            .O(N__19987),
            .I(\nx.n3108 ));
    InMux I__2081 (
            .O(N__19980),
            .I(N__19977));
    LocalMux I__2080 (
            .O(N__19977),
            .I(\nx.n3165 ));
    InMux I__2079 (
            .O(N__19974),
            .I(N__19970));
    InMux I__2078 (
            .O(N__19973),
            .I(N__19967));
    LocalMux I__2077 (
            .O(N__19970),
            .I(N__19961));
    LocalMux I__2076 (
            .O(N__19967),
            .I(N__19961));
    InMux I__2075 (
            .O(N__19966),
            .I(N__19958));
    Odrv4 I__2074 (
            .O(N__19961),
            .I(\nx.n3098 ));
    LocalMux I__2073 (
            .O(N__19958),
            .I(\nx.n3098 ));
    CascadeMux I__2072 (
            .O(N__19953),
            .I(\nx.n13_adj_696_cascade_ ));
    InMux I__2071 (
            .O(N__19950),
            .I(N__19947));
    LocalMux I__2070 (
            .O(N__19947),
            .I(\nx.n31_adj_702 ));
    InMux I__2069 (
            .O(N__19944),
            .I(N__19941));
    LocalMux I__2068 (
            .O(N__19941),
            .I(\nx.n21_adj_701 ));
    CascadeMux I__2067 (
            .O(N__19938),
            .I(\nx.n12325_cascade_ ));
    InMux I__2066 (
            .O(N__19935),
            .I(N__19932));
    LocalMux I__2065 (
            .O(N__19932),
            .I(\nx.n12339 ));
    CascadeMux I__2064 (
            .O(N__19929),
            .I(N__19926));
    InMux I__2063 (
            .O(N__19926),
            .I(N__19923));
    LocalMux I__2062 (
            .O(N__19923),
            .I(\nx.n12347 ));
    CascadeMux I__2061 (
            .O(N__19920),
            .I(N__19917));
    InMux I__2060 (
            .O(N__19917),
            .I(N__19912));
    InMux I__2059 (
            .O(N__19916),
            .I(N__19907));
    InMux I__2058 (
            .O(N__19915),
            .I(N__19907));
    LocalMux I__2057 (
            .O(N__19912),
            .I(N__19904));
    LocalMux I__2056 (
            .O(N__19907),
            .I(\nx.n3103 ));
    Odrv4 I__2055 (
            .O(N__19904),
            .I(\nx.n3103 ));
    InMux I__2054 (
            .O(N__19899),
            .I(N__19895));
    InMux I__2053 (
            .O(N__19898),
            .I(N__19892));
    LocalMux I__2052 (
            .O(N__19895),
            .I(N__19889));
    LocalMux I__2051 (
            .O(N__19892),
            .I(N__19886));
    Odrv4 I__2050 (
            .O(N__19889),
            .I(\nx.n3097 ));
    Odrv4 I__2049 (
            .O(N__19886),
            .I(\nx.n3097 ));
    InMux I__2048 (
            .O(N__19881),
            .I(N__19878));
    LocalMux I__2047 (
            .O(N__19878),
            .I(N__19875));
    Odrv4 I__2046 (
            .O(N__19875),
            .I(\nx.n3164 ));
    CascadeMux I__2045 (
            .O(N__19872),
            .I(\nx.n3097_cascade_ ));
    InMux I__2044 (
            .O(N__19869),
            .I(N__19866));
    LocalMux I__2043 (
            .O(N__19866),
            .I(N__19863));
    Odrv4 I__2042 (
            .O(N__19863),
            .I(\nx.n3168 ));
    CascadeMux I__2041 (
            .O(N__19860),
            .I(\nx.n35_adj_699_cascade_ ));
    CascadeMux I__2040 (
            .O(N__19857),
            .I(N__19854));
    InMux I__2039 (
            .O(N__19854),
            .I(N__19851));
    LocalMux I__2038 (
            .O(N__19851),
            .I(N__19847));
    InMux I__2037 (
            .O(N__19850),
            .I(N__19843));
    Span4Mux_v I__2036 (
            .O(N__19847),
            .I(N__19840));
    InMux I__2035 (
            .O(N__19846),
            .I(N__19837));
    LocalMux I__2034 (
            .O(N__19843),
            .I(\nx.n3101 ));
    Odrv4 I__2033 (
            .O(N__19840),
            .I(\nx.n3101 ));
    LocalMux I__2032 (
            .O(N__19837),
            .I(\nx.n3101 ));
    InMux I__2031 (
            .O(N__19830),
            .I(N__19827));
    LocalMux I__2030 (
            .O(N__19827),
            .I(\nx.n12337 ));
    CascadeMux I__2029 (
            .O(N__19824),
            .I(N__19819));
    InMux I__2028 (
            .O(N__19823),
            .I(N__19816));
    InMux I__2027 (
            .O(N__19822),
            .I(N__19813));
    InMux I__2026 (
            .O(N__19819),
            .I(N__19810));
    LocalMux I__2025 (
            .O(N__19816),
            .I(\nx.n3109 ));
    LocalMux I__2024 (
            .O(N__19813),
            .I(\nx.n3109 ));
    LocalMux I__2023 (
            .O(N__19810),
            .I(\nx.n3109 ));
    InMux I__2022 (
            .O(N__19803),
            .I(N__19800));
    LocalMux I__2021 (
            .O(N__19800),
            .I(\nx.n12349 ));
    CascadeMux I__2020 (
            .O(N__19797),
            .I(N__19794));
    InMux I__2019 (
            .O(N__19794),
            .I(N__19790));
    InMux I__2018 (
            .O(N__19793),
            .I(N__19787));
    LocalMux I__2017 (
            .O(N__19790),
            .I(N__19784));
    LocalMux I__2016 (
            .O(N__19787),
            .I(N__19779));
    Span4Mux_v I__2015 (
            .O(N__19784),
            .I(N__19779));
    Odrv4 I__2014 (
            .O(N__19779),
            .I(\nx.n3096 ));
    CascadeMux I__2013 (
            .O(N__19776),
            .I(\nx.n3096_cascade_ ));
    InMux I__2012 (
            .O(N__19773),
            .I(N__19770));
    LocalMux I__2011 (
            .O(N__19770),
            .I(N__19767));
    Odrv4 I__2010 (
            .O(N__19767),
            .I(\nx.n47_adj_694 ));
    CascadeMux I__2009 (
            .O(N__19764),
            .I(N__19761));
    InMux I__2008 (
            .O(N__19761),
            .I(N__19758));
    LocalMux I__2007 (
            .O(N__19758),
            .I(\nx.n45 ));
    CascadeMux I__2006 (
            .O(N__19755),
            .I(\nx.n49_cascade_ ));
    CascadeMux I__2005 (
            .O(N__19752),
            .I(\nx.n3017_cascade_ ));
    InMux I__2004 (
            .O(N__19749),
            .I(N__19745));
    InMux I__2003 (
            .O(N__19748),
            .I(N__19742));
    LocalMux I__2002 (
            .O(N__19745),
            .I(N__19739));
    LocalMux I__2001 (
            .O(N__19742),
            .I(N__19736));
    Span4Mux_v I__2000 (
            .O(N__19739),
            .I(N__19733));
    Odrv4 I__1999 (
            .O(N__19736),
            .I(\nx.n3086 ));
    Odrv4 I__1998 (
            .O(N__19733),
            .I(\nx.n3086 ));
    InMux I__1997 (
            .O(N__19728),
            .I(N__19724));
    InMux I__1996 (
            .O(N__19727),
            .I(N__19721));
    LocalMux I__1995 (
            .O(N__19724),
            .I(N__19718));
    LocalMux I__1994 (
            .O(N__19721),
            .I(N__19714));
    Span4Mux_v I__1993 (
            .O(N__19718),
            .I(N__19711));
    InMux I__1992 (
            .O(N__19717),
            .I(N__19708));
    Odrv4 I__1991 (
            .O(N__19714),
            .I(\nx.n3087 ));
    Odrv4 I__1990 (
            .O(N__19711),
            .I(\nx.n3087 ));
    LocalMux I__1989 (
            .O(N__19708),
            .I(\nx.n3087 ));
    CascadeMux I__1988 (
            .O(N__19701),
            .I(\nx.n3086_cascade_ ));
    InMux I__1987 (
            .O(N__19698),
            .I(N__19695));
    LocalMux I__1986 (
            .O(N__19695),
            .I(N__19691));
    InMux I__1985 (
            .O(N__19694),
            .I(N__19687));
    Span4Mux_v I__1984 (
            .O(N__19691),
            .I(N__19684));
    InMux I__1983 (
            .O(N__19690),
            .I(N__19681));
    LocalMux I__1982 (
            .O(N__19687),
            .I(\nx.n3085 ));
    Odrv4 I__1981 (
            .O(N__19684),
            .I(\nx.n3085 ));
    LocalMux I__1980 (
            .O(N__19681),
            .I(\nx.n3085 ));
    InMux I__1979 (
            .O(N__19674),
            .I(N__19671));
    LocalMux I__1978 (
            .O(N__19671),
            .I(\nx.n42_adj_689 ));
    CascadeMux I__1977 (
            .O(N__19668),
            .I(N__19665));
    InMux I__1976 (
            .O(N__19665),
            .I(N__19662));
    LocalMux I__1975 (
            .O(N__19662),
            .I(\nx.color_bit_N_571_4 ));
    InMux I__1974 (
            .O(N__19659),
            .I(N__19656));
    LocalMux I__1973 (
            .O(N__19656),
            .I(\nx.n13158 ));
    InMux I__1972 (
            .O(N__19653),
            .I(N__19650));
    LocalMux I__1971 (
            .O(N__19650),
            .I(\nx.n59 ));
    CascadeMux I__1970 (
            .O(N__19647),
            .I(N__19644));
    InMux I__1969 (
            .O(N__19644),
            .I(N__19641));
    LocalMux I__1968 (
            .O(N__19641),
            .I(\nx.n12371 ));
    InMux I__1967 (
            .O(N__19638),
            .I(N__19635));
    LocalMux I__1966 (
            .O(N__19635),
            .I(N__19632));
    Span4Mux_v I__1965 (
            .O(N__19632),
            .I(N__19629));
    Odrv4 I__1964 (
            .O(N__19629),
            .I(\nx.n13042 ));
    InMux I__1963 (
            .O(N__19626),
            .I(N__19623));
    LocalMux I__1962 (
            .O(N__19623),
            .I(\nx.n10947 ));
    CascadeMux I__1961 (
            .O(N__19620),
            .I(\nx.n10947_cascade_ ));
    InMux I__1960 (
            .O(N__19617),
            .I(N__19611));
    InMux I__1959 (
            .O(N__19616),
            .I(N__19611));
    LocalMux I__1958 (
            .O(N__19611),
            .I(\nx.n10975 ));
    CascadeMux I__1957 (
            .O(N__19608),
            .I(\nx.n3008_cascade_ ));
    CascadeMux I__1956 (
            .O(N__19605),
            .I(N__19600));
    CascadeMux I__1955 (
            .O(N__19604),
            .I(N__19597));
    InMux I__1954 (
            .O(N__19603),
            .I(N__19587));
    InMux I__1953 (
            .O(N__19600),
            .I(N__19587));
    InMux I__1952 (
            .O(N__19597),
            .I(N__19587));
    CascadeMux I__1951 (
            .O(N__19596),
            .I(N__19583));
    InMux I__1950 (
            .O(N__19595),
            .I(N__19575));
    InMux I__1949 (
            .O(N__19594),
            .I(N__19575));
    LocalMux I__1948 (
            .O(N__19587),
            .I(N__19571));
    InMux I__1947 (
            .O(N__19586),
            .I(N__19566));
    InMux I__1946 (
            .O(N__19583),
            .I(N__19566));
    InMux I__1945 (
            .O(N__19582),
            .I(N__19561));
    InMux I__1944 (
            .O(N__19581),
            .I(N__19556));
    InMux I__1943 (
            .O(N__19580),
            .I(N__19556));
    LocalMux I__1942 (
            .O(N__19575),
            .I(N__19553));
    InMux I__1941 (
            .O(N__19574),
            .I(N__19550));
    Span4Mux_v I__1940 (
            .O(N__19571),
            .I(N__19545));
    LocalMux I__1939 (
            .O(N__19566),
            .I(N__19545));
    InMux I__1938 (
            .O(N__19565),
            .I(N__19540));
    InMux I__1937 (
            .O(N__19564),
            .I(N__19540));
    LocalMux I__1936 (
            .O(N__19561),
            .I(state_0_adj_727));
    LocalMux I__1935 (
            .O(N__19556),
            .I(state_0_adj_727));
    Odrv4 I__1934 (
            .O(N__19553),
            .I(state_0_adj_727));
    LocalMux I__1933 (
            .O(N__19550),
            .I(state_0_adj_727));
    Odrv4 I__1932 (
            .O(N__19545),
            .I(state_0_adj_727));
    LocalMux I__1931 (
            .O(N__19540),
            .I(state_0_adj_727));
    InMux I__1930 (
            .O(N__19527),
            .I(N__19524));
    LocalMux I__1929 (
            .O(N__19524),
            .I(N__19520));
    InMux I__1928 (
            .O(N__19523),
            .I(N__19517));
    Span4Mux_v I__1927 (
            .O(N__19520),
            .I(N__19505));
    LocalMux I__1926 (
            .O(N__19517),
            .I(N__19505));
    CascadeMux I__1925 (
            .O(N__19516),
            .I(N__19501));
    CascadeMux I__1924 (
            .O(N__19515),
            .I(N__19497));
    InMux I__1923 (
            .O(N__19514),
            .I(N__19492));
    InMux I__1922 (
            .O(N__19513),
            .I(N__19489));
    InMux I__1921 (
            .O(N__19512),
            .I(N__19484));
    InMux I__1920 (
            .O(N__19511),
            .I(N__19484));
    InMux I__1919 (
            .O(N__19510),
            .I(N__19481));
    Span4Mux_v I__1918 (
            .O(N__19505),
            .I(N__19476));
    InMux I__1917 (
            .O(N__19504),
            .I(N__19473));
    InMux I__1916 (
            .O(N__19501),
            .I(N__19470));
    InMux I__1915 (
            .O(N__19500),
            .I(N__19461));
    InMux I__1914 (
            .O(N__19497),
            .I(N__19461));
    InMux I__1913 (
            .O(N__19496),
            .I(N__19461));
    InMux I__1912 (
            .O(N__19495),
            .I(N__19461));
    LocalMux I__1911 (
            .O(N__19492),
            .I(N__19452));
    LocalMux I__1910 (
            .O(N__19489),
            .I(N__19452));
    LocalMux I__1909 (
            .O(N__19484),
            .I(N__19452));
    LocalMux I__1908 (
            .O(N__19481),
            .I(N__19452));
    InMux I__1907 (
            .O(N__19480),
            .I(N__19449));
    InMux I__1906 (
            .O(N__19479),
            .I(N__19446));
    Odrv4 I__1905 (
            .O(N__19476),
            .I(state_1_adj_726));
    LocalMux I__1904 (
            .O(N__19473),
            .I(state_1_adj_726));
    LocalMux I__1903 (
            .O(N__19470),
            .I(state_1_adj_726));
    LocalMux I__1902 (
            .O(N__19461),
            .I(state_1_adj_726));
    Odrv4 I__1901 (
            .O(N__19452),
            .I(state_1_adj_726));
    LocalMux I__1900 (
            .O(N__19449),
            .I(state_1_adj_726));
    LocalMux I__1899 (
            .O(N__19446),
            .I(state_1_adj_726));
    CEMux I__1898 (
            .O(N__19431),
            .I(N__19427));
    InMux I__1897 (
            .O(N__19430),
            .I(N__19424));
    LocalMux I__1896 (
            .O(N__19427),
            .I(n7239));
    LocalMux I__1895 (
            .O(N__19424),
            .I(n7239));
    SRMux I__1894 (
            .O(N__19419),
            .I(N__19416));
    LocalMux I__1893 (
            .O(N__19416),
            .I(N__19413));
    Odrv4 I__1892 (
            .O(N__19413),
            .I(\nx.n7392 ));
    InMux I__1891 (
            .O(N__19410),
            .I(N__19407));
    LocalMux I__1890 (
            .O(N__19407),
            .I(\nx.n13155 ));
    CascadeMux I__1889 (
            .O(N__19404),
            .I(\nx.n13456_cascade_ ));
    InMux I__1888 (
            .O(N__19401),
            .I(N__19398));
    LocalMux I__1887 (
            .O(N__19398),
            .I(\nx.n13156 ));
    InMux I__1886 (
            .O(N__19395),
            .I(N__19392));
    LocalMux I__1885 (
            .O(N__19392),
            .I(\nx.n13459 ));
    InMux I__1884 (
            .O(N__19389),
            .I(N__19382));
    InMux I__1883 (
            .O(N__19388),
            .I(N__19382));
    InMux I__1882 (
            .O(N__19387),
            .I(N__19379));
    LocalMux I__1881 (
            .O(N__19382),
            .I(N__19374));
    LocalMux I__1880 (
            .O(N__19379),
            .I(N__19371));
    InMux I__1879 (
            .O(N__19378),
            .I(N__19366));
    InMux I__1878 (
            .O(N__19377),
            .I(N__19366));
    Span4Mux_v I__1877 (
            .O(N__19374),
            .I(N__19363));
    Span4Mux_s1_h I__1876 (
            .O(N__19371),
            .I(N__19358));
    LocalMux I__1875 (
            .O(N__19366),
            .I(N__19358));
    Odrv4 I__1874 (
            .O(N__19363),
            .I(\nx.n4_adj_642 ));
    Odrv4 I__1873 (
            .O(N__19358),
            .I(\nx.n4_adj_642 ));
    InMux I__1872 (
            .O(N__19353),
            .I(N__19349));
    InMux I__1871 (
            .O(N__19352),
            .I(N__19346));
    LocalMux I__1870 (
            .O(N__19349),
            .I(neo_pixel_transmitter_t0_26));
    LocalMux I__1869 (
            .O(N__19346),
            .I(neo_pixel_transmitter_t0_26));
    InMux I__1868 (
            .O(N__19341),
            .I(N__19337));
    InMux I__1867 (
            .O(N__19340),
            .I(N__19334));
    LocalMux I__1866 (
            .O(N__19337),
            .I(neo_pixel_transmitter_t0_16));
    LocalMux I__1865 (
            .O(N__19334),
            .I(neo_pixel_transmitter_t0_16));
    InMux I__1864 (
            .O(N__19329),
            .I(N__19326));
    LocalMux I__1863 (
            .O(N__19326),
            .I(neopxl_color_prev_5));
    InMux I__1862 (
            .O(N__19323),
            .I(N__19320));
    LocalMux I__1861 (
            .O(N__19320),
            .I(N__19317));
    Odrv4 I__1860 (
            .O(N__19317),
            .I(n10_adj_776));
    InMux I__1859 (
            .O(N__19314),
            .I(N__19308));
    InMux I__1858 (
            .O(N__19313),
            .I(N__19308));
    LocalMux I__1857 (
            .O(N__19308),
            .I(neo_pixel_transmitter_t0_3));
    InMux I__1856 (
            .O(N__19305),
            .I(N__19302));
    LocalMux I__1855 (
            .O(N__19302),
            .I(n12_adj_774));
    InMux I__1854 (
            .O(N__19299),
            .I(N__19295));
    InMux I__1853 (
            .O(N__19298),
            .I(N__19292));
    LocalMux I__1852 (
            .O(N__19295),
            .I(neo_pixel_transmitter_t0_12));
    LocalMux I__1851 (
            .O(N__19292),
            .I(neo_pixel_transmitter_t0_12));
    CascadeMux I__1850 (
            .O(N__19287),
            .I(N__19283));
    InMux I__1849 (
            .O(N__19286),
            .I(N__19278));
    InMux I__1848 (
            .O(N__19283),
            .I(N__19273));
    InMux I__1847 (
            .O(N__19282),
            .I(N__19273));
    InMux I__1846 (
            .O(N__19281),
            .I(N__19268));
    LocalMux I__1845 (
            .O(N__19278),
            .I(N__19257));
    LocalMux I__1844 (
            .O(N__19273),
            .I(N__19257));
    InMux I__1843 (
            .O(N__19272),
            .I(N__19254));
    InMux I__1842 (
            .O(N__19271),
            .I(N__19251));
    LocalMux I__1841 (
            .O(N__19268),
            .I(N__19248));
    InMux I__1840 (
            .O(N__19267),
            .I(N__19243));
    InMux I__1839 (
            .O(N__19266),
            .I(N__19243));
    InMux I__1838 (
            .O(N__19265),
            .I(N__19240));
    InMux I__1837 (
            .O(N__19264),
            .I(N__19237));
    InMux I__1836 (
            .O(N__19263),
            .I(N__19232));
    InMux I__1835 (
            .O(N__19262),
            .I(N__19232));
    Sp12to4 I__1834 (
            .O(N__19257),
            .I(N__19227));
    LocalMux I__1833 (
            .O(N__19254),
            .I(N__19227));
    LocalMux I__1832 (
            .O(N__19251),
            .I(\nx.neo_pixel_transmitter_done ));
    Odrv4 I__1831 (
            .O(N__19248),
            .I(\nx.neo_pixel_transmitter_done ));
    LocalMux I__1830 (
            .O(N__19243),
            .I(\nx.neo_pixel_transmitter_done ));
    LocalMux I__1829 (
            .O(N__19240),
            .I(\nx.neo_pixel_transmitter_done ));
    LocalMux I__1828 (
            .O(N__19237),
            .I(\nx.neo_pixel_transmitter_done ));
    LocalMux I__1827 (
            .O(N__19232),
            .I(\nx.neo_pixel_transmitter_done ));
    Odrv12 I__1826 (
            .O(N__19227),
            .I(\nx.neo_pixel_transmitter_done ));
    CascadeMux I__1825 (
            .O(N__19212),
            .I(\nx.n11487_cascade_ ));
    InMux I__1824 (
            .O(N__19209),
            .I(N__19206));
    LocalMux I__1823 (
            .O(N__19206),
            .I(\nx.n103 ));
    CascadeMux I__1822 (
            .O(N__19203),
            .I(N__19200));
    InMux I__1821 (
            .O(N__19200),
            .I(N__19197));
    LocalMux I__1820 (
            .O(N__19197),
            .I(N__19194));
    Span4Mux_v I__1819 (
            .O(N__19194),
            .I(N__19191));
    Odrv4 I__1818 (
            .O(N__19191),
            .I(n9_adj_777));
    InMux I__1817 (
            .O(N__19188),
            .I(N__19185));
    LocalMux I__1816 (
            .O(N__19185),
            .I(neopxl_color_prev_4));
    InMux I__1815 (
            .O(N__19182),
            .I(N__19178));
    CascadeMux I__1814 (
            .O(N__19181),
            .I(N__19175));
    LocalMux I__1813 (
            .O(N__19178),
            .I(N__19170));
    InMux I__1812 (
            .O(N__19175),
            .I(N__19165));
    InMux I__1811 (
            .O(N__19174),
            .I(N__19165));
    InMux I__1810 (
            .O(N__19173),
            .I(N__19162));
    Odrv4 I__1809 (
            .O(N__19170),
            .I(\nx.n10918 ));
    LocalMux I__1808 (
            .O(N__19165),
            .I(\nx.n10918 ));
    LocalMux I__1807 (
            .O(N__19162),
            .I(\nx.n10918 ));
    InMux I__1806 (
            .O(N__19155),
            .I(N__19151));
    InMux I__1805 (
            .O(N__19154),
            .I(N__19146));
    LocalMux I__1804 (
            .O(N__19151),
            .I(N__19139));
    InMux I__1803 (
            .O(N__19150),
            .I(N__19134));
    InMux I__1802 (
            .O(N__19149),
            .I(N__19134));
    LocalMux I__1801 (
            .O(N__19146),
            .I(N__19131));
    InMux I__1800 (
            .O(N__19145),
            .I(N__19126));
    InMux I__1799 (
            .O(N__19144),
            .I(N__19126));
    InMux I__1798 (
            .O(N__19143),
            .I(N__19123));
    InMux I__1797 (
            .O(N__19142),
            .I(N__19119));
    Span4Mux_h I__1796 (
            .O(N__19139),
            .I(N__19108));
    LocalMux I__1795 (
            .O(N__19134),
            .I(N__19108));
    Span4Mux_v I__1794 (
            .O(N__19131),
            .I(N__19108));
    LocalMux I__1793 (
            .O(N__19126),
            .I(N__19108));
    LocalMux I__1792 (
            .O(N__19123),
            .I(N__19108));
    InMux I__1791 (
            .O(N__19122),
            .I(N__19105));
    LocalMux I__1790 (
            .O(N__19119),
            .I(N__19102));
    Span4Mux_v I__1789 (
            .O(N__19108),
            .I(N__19099));
    LocalMux I__1788 (
            .O(N__19105),
            .I(\nx.start ));
    Odrv12 I__1787 (
            .O(N__19102),
            .I(\nx.start ));
    Odrv4 I__1786 (
            .O(N__19099),
            .I(\nx.start ));
    CascadeMux I__1785 (
            .O(N__19092),
            .I(\nx.n18_adj_711_cascade_ ));
    InMux I__1784 (
            .O(N__19089),
            .I(N__19086));
    LocalMux I__1783 (
            .O(N__19086),
            .I(\nx.n20_adj_712 ));
    InMux I__1782 (
            .O(N__19083),
            .I(N__19077));
    InMux I__1781 (
            .O(N__19082),
            .I(N__19077));
    LocalMux I__1780 (
            .O(N__19077),
            .I(neo_pixel_transmitter_t0_6));
    InMux I__1779 (
            .O(N__19074),
            .I(N__19068));
    InMux I__1778 (
            .O(N__19073),
            .I(N__19068));
    LocalMux I__1777 (
            .O(N__19068),
            .I(neo_pixel_transmitter_t0_14));
    InMux I__1776 (
            .O(N__19065),
            .I(N__19061));
    InMux I__1775 (
            .O(N__19064),
            .I(N__19058));
    LocalMux I__1774 (
            .O(N__19061),
            .I(N__19055));
    LocalMux I__1773 (
            .O(N__19058),
            .I(neo_pixel_transmitter_t0_5));
    Odrv4 I__1772 (
            .O(N__19055),
            .I(neo_pixel_transmitter_t0_5));
    InMux I__1771 (
            .O(N__19050),
            .I(N__19044));
    InMux I__1770 (
            .O(N__19049),
            .I(N__19044));
    LocalMux I__1769 (
            .O(N__19044),
            .I(neo_pixel_transmitter_t0_23));
    CascadeMux I__1768 (
            .O(N__19041),
            .I(N__19038));
    InMux I__1767 (
            .O(N__19038),
            .I(N__19032));
    InMux I__1766 (
            .O(N__19037),
            .I(N__19032));
    LocalMux I__1765 (
            .O(N__19032),
            .I(neo_pixel_transmitter_t0_24));
    CascadeMux I__1764 (
            .O(N__19029),
            .I(\nx.n7_adj_713_cascade_ ));
    CEMux I__1763 (
            .O(N__19026),
            .I(N__19023));
    LocalMux I__1762 (
            .O(N__19023),
            .I(\nx.n13491 ));
    CascadeMux I__1761 (
            .O(N__19020),
            .I(\nx.n12933_cascade_ ));
    InMux I__1760 (
            .O(N__19017),
            .I(N__19014));
    LocalMux I__1759 (
            .O(N__19014),
            .I(\nx.n12939 ));
    InMux I__1758 (
            .O(N__19011),
            .I(\nx.n10459 ));
    InMux I__1757 (
            .O(N__19008),
            .I(bfn_1_32_0_));
    InMux I__1756 (
            .O(N__19005),
            .I(N__19001));
    CascadeMux I__1755 (
            .O(N__19004),
            .I(N__18998));
    LocalMux I__1754 (
            .O(N__19001),
            .I(N__18995));
    InMux I__1753 (
            .O(N__18998),
            .I(N__18992));
    Odrv4 I__1752 (
            .O(N__18995),
            .I(\nx.n1203 ));
    LocalMux I__1751 (
            .O(N__18992),
            .I(\nx.n1203 ));
    InMux I__1750 (
            .O(N__18987),
            .I(N__18984));
    LocalMux I__1749 (
            .O(N__18984),
            .I(\nx.n1270 ));
    CascadeMux I__1748 (
            .O(N__18981),
            .I(\nx.n1302_cascade_ ));
    InMux I__1747 (
            .O(N__18978),
            .I(N__18975));
    LocalMux I__1746 (
            .O(N__18975),
            .I(\nx.n1276 ));
    InMux I__1745 (
            .O(N__18972),
            .I(N__18968));
    CascadeMux I__1744 (
            .O(N__18971),
            .I(N__18964));
    LocalMux I__1743 (
            .O(N__18968),
            .I(N__18961));
    InMux I__1742 (
            .O(N__18967),
            .I(N__18958));
    InMux I__1741 (
            .O(N__18964),
            .I(N__18955));
    Odrv4 I__1740 (
            .O(N__18961),
            .I(\nx.n1209 ));
    LocalMux I__1739 (
            .O(N__18958),
            .I(\nx.n1209 ));
    LocalMux I__1738 (
            .O(N__18955),
            .I(\nx.n1209 ));
    CascadeMux I__1737 (
            .O(N__18948),
            .I(\nx.n1206_cascade_ ));
    InMux I__1736 (
            .O(N__18945),
            .I(N__18942));
    LocalMux I__1735 (
            .O(N__18942),
            .I(\nx.n1273 ));
    CEMux I__1734 (
            .O(N__18939),
            .I(N__18936));
    LocalMux I__1733 (
            .O(N__18936),
            .I(N__18933));
    Span4Mux_v I__1732 (
            .O(N__18933),
            .I(N__18930));
    Span4Mux_s1_h I__1731 (
            .O(N__18930),
            .I(N__18927));
    Odrv4 I__1730 (
            .O(N__18927),
            .I(\nx.n7 ));
    CascadeMux I__1729 (
            .O(N__18924),
            .I(\nx.n1203_cascade_ ));
    CascadeMux I__1728 (
            .O(N__18921),
            .I(\nx.n1208_cascade_ ));
    InMux I__1727 (
            .O(N__18918),
            .I(bfn_1_31_0_));
    InMux I__1726 (
            .O(N__18915),
            .I(\nx.n10453 ));
    InMux I__1725 (
            .O(N__18912),
            .I(\nx.n10454 ));
    InMux I__1724 (
            .O(N__18909),
            .I(\nx.n10455 ));
    InMux I__1723 (
            .O(N__18906),
            .I(\nx.n10456 ));
    InMux I__1722 (
            .O(N__18903),
            .I(\nx.n10457 ));
    InMux I__1721 (
            .O(N__18900),
            .I(\nx.n10458 ));
    InMux I__1720 (
            .O(N__18897),
            .I(N__18894));
    LocalMux I__1719 (
            .O(N__18894),
            .I(N__18891));
    Odrv12 I__1718 (
            .O(N__18891),
            .I(\nx.n3152 ));
    InMux I__1717 (
            .O(N__18888),
            .I(\nx.n10912 ));
    InMux I__1716 (
            .O(N__18885),
            .I(\nx.n10913 ));
    InMux I__1715 (
            .O(N__18882),
            .I(\nx.n10914 ));
    CascadeMux I__1714 (
            .O(N__18879),
            .I(\nx.n10_adj_619_cascade_ ));
    CascadeMux I__1713 (
            .O(N__18876),
            .I(\nx.n12_adj_621_cascade_ ));
    CascadeMux I__1712 (
            .O(N__18873),
            .I(\nx.n1136_cascade_ ));
    InMux I__1711 (
            .O(N__18870),
            .I(bfn_1_28_0_));
    InMux I__1710 (
            .O(N__18867),
            .I(\nx.n10904 ));
    InMux I__1709 (
            .O(N__18864),
            .I(\nx.n10905 ));
    InMux I__1708 (
            .O(N__18861),
            .I(\nx.n10906 ));
    InMux I__1707 (
            .O(N__18858),
            .I(\nx.n10907 ));
    InMux I__1706 (
            .O(N__18855),
            .I(\nx.n10908 ));
    InMux I__1705 (
            .O(N__18852),
            .I(\nx.n10909 ));
    CascadeMux I__1704 (
            .O(N__18849),
            .I(N__18846));
    InMux I__1703 (
            .O(N__18846),
            .I(N__18843));
    LocalMux I__1702 (
            .O(N__18843),
            .I(N__18840));
    Span4Mux_v I__1701 (
            .O(N__18840),
            .I(N__18837));
    Odrv4 I__1700 (
            .O(N__18837),
            .I(\nx.n3154 ));
    InMux I__1699 (
            .O(N__18834),
            .I(\nx.n10910 ));
    InMux I__1698 (
            .O(N__18831),
            .I(N__18828));
    LocalMux I__1697 (
            .O(N__18828),
            .I(N__18825));
    Span4Mux_v I__1696 (
            .O(N__18825),
            .I(N__18822));
    Odrv4 I__1695 (
            .O(N__18822),
            .I(\nx.n3153 ));
    InMux I__1694 (
            .O(N__18819),
            .I(bfn_1_29_0_));
    CascadeMux I__1693 (
            .O(N__18816),
            .I(N__18812));
    InMux I__1692 (
            .O(N__18815),
            .I(N__18808));
    InMux I__1691 (
            .O(N__18812),
            .I(N__18805));
    InMux I__1690 (
            .O(N__18811),
            .I(N__18802));
    LocalMux I__1689 (
            .O(N__18808),
            .I(N__18797));
    LocalMux I__1688 (
            .O(N__18805),
            .I(N__18797));
    LocalMux I__1687 (
            .O(N__18802),
            .I(\nx.n3102 ));
    Odrv4 I__1686 (
            .O(N__18797),
            .I(\nx.n3102 ));
    InMux I__1685 (
            .O(N__18792),
            .I(N__18789));
    LocalMux I__1684 (
            .O(N__18789),
            .I(N__18786));
    Odrv4 I__1683 (
            .O(N__18786),
            .I(\nx.n3169 ));
    InMux I__1682 (
            .O(N__18783),
            .I(bfn_1_27_0_));
    InMux I__1681 (
            .O(N__18780),
            .I(\nx.n10896 ));
    CascadeMux I__1680 (
            .O(N__18777),
            .I(N__18774));
    InMux I__1679 (
            .O(N__18774),
            .I(N__18771));
    LocalMux I__1678 (
            .O(N__18771),
            .I(N__18767));
    InMux I__1677 (
            .O(N__18770),
            .I(N__18764));
    Odrv4 I__1676 (
            .O(N__18767),
            .I(\nx.n3100 ));
    LocalMux I__1675 (
            .O(N__18764),
            .I(\nx.n3100 ));
    InMux I__1674 (
            .O(N__18759),
            .I(N__18756));
    LocalMux I__1673 (
            .O(N__18756),
            .I(N__18753));
    Odrv4 I__1672 (
            .O(N__18753),
            .I(\nx.n3167 ));
    InMux I__1671 (
            .O(N__18750),
            .I(\nx.n10897 ));
    InMux I__1670 (
            .O(N__18747),
            .I(\nx.n10898 ));
    InMux I__1669 (
            .O(N__18744),
            .I(\nx.n10899 ));
    InMux I__1668 (
            .O(N__18741),
            .I(\nx.n10900 ));
    CascadeMux I__1667 (
            .O(N__18738),
            .I(N__18735));
    InMux I__1666 (
            .O(N__18735),
            .I(N__18732));
    LocalMux I__1665 (
            .O(N__18732),
            .I(N__18729));
    Odrv4 I__1664 (
            .O(N__18729),
            .I(\nx.n3163 ));
    InMux I__1663 (
            .O(N__18726),
            .I(\nx.n10901 ));
    InMux I__1662 (
            .O(N__18723),
            .I(\nx.n10902 ));
    CascadeMux I__1661 (
            .O(N__18720),
            .I(\nx.n3116_cascade_ ));
    InMux I__1660 (
            .O(N__18717),
            .I(bfn_1_26_0_));
    InMux I__1659 (
            .O(N__18714),
            .I(N__18711));
    LocalMux I__1658 (
            .O(N__18711),
            .I(N__18708));
    Span4Mux_h I__1657 (
            .O(N__18708),
            .I(N__18705));
    Odrv4 I__1656 (
            .O(N__18705),
            .I(\nx.n3176 ));
    InMux I__1655 (
            .O(N__18702),
            .I(\nx.n10888 ));
    InMux I__1654 (
            .O(N__18699),
            .I(\nx.n10889 ));
    InMux I__1653 (
            .O(N__18696),
            .I(\nx.n10890 ));
    InMux I__1652 (
            .O(N__18693),
            .I(N__18689));
    InMux I__1651 (
            .O(N__18692),
            .I(N__18686));
    LocalMux I__1650 (
            .O(N__18689),
            .I(N__18681));
    LocalMux I__1649 (
            .O(N__18686),
            .I(N__18681));
    Odrv4 I__1648 (
            .O(N__18681),
            .I(\nx.n3106 ));
    InMux I__1647 (
            .O(N__18678),
            .I(N__18675));
    LocalMux I__1646 (
            .O(N__18675),
            .I(N__18672));
    Odrv12 I__1645 (
            .O(N__18672),
            .I(\nx.n3173 ));
    InMux I__1644 (
            .O(N__18669),
            .I(\nx.n10891 ));
    CascadeMux I__1643 (
            .O(N__18666),
            .I(N__18662));
    CascadeMux I__1642 (
            .O(N__18665),
            .I(N__18659));
    InMux I__1641 (
            .O(N__18662),
            .I(N__18656));
    InMux I__1640 (
            .O(N__18659),
            .I(N__18653));
    LocalMux I__1639 (
            .O(N__18656),
            .I(N__18650));
    LocalMux I__1638 (
            .O(N__18653),
            .I(\nx.n3105 ));
    Odrv4 I__1637 (
            .O(N__18650),
            .I(\nx.n3105 ));
    InMux I__1636 (
            .O(N__18645),
            .I(N__18642));
    LocalMux I__1635 (
            .O(N__18642),
            .I(N__18639));
    Odrv4 I__1634 (
            .O(N__18639),
            .I(\nx.n3172 ));
    InMux I__1633 (
            .O(N__18636),
            .I(\nx.n10892 ));
    InMux I__1632 (
            .O(N__18633),
            .I(\nx.n10893 ));
    InMux I__1631 (
            .O(N__18630),
            .I(N__18627));
    LocalMux I__1630 (
            .O(N__18627),
            .I(\nx.n3170 ));
    InMux I__1629 (
            .O(N__18624),
            .I(\nx.n10894 ));
    CascadeMux I__1628 (
            .O(N__18621),
            .I(\nx.n3100_cascade_ ));
    CascadeMux I__1627 (
            .O(N__18618),
            .I(\nx.n29_adj_697_cascade_ ));
    CascadeMux I__1626 (
            .O(N__18615),
            .I(\nx.n12331_cascade_ ));
    InMux I__1625 (
            .O(N__18612),
            .I(N__18609));
    LocalMux I__1624 (
            .O(N__18609),
            .I(\nx.n12335 ));
    CascadeMux I__1623 (
            .O(N__18606),
            .I(\nx.n37_adj_695_cascade_ ));
    InMux I__1622 (
            .O(N__18603),
            .I(N__18600));
    LocalMux I__1621 (
            .O(N__18600),
            .I(\nx.n12333 ));
    CascadeMux I__1620 (
            .O(N__18597),
            .I(\nx.n31_adj_691_cascade_ ));
    CascadeMux I__1619 (
            .O(N__18594),
            .I(\nx.n49_adj_693_cascade_ ));
    InMux I__1618 (
            .O(N__18591),
            .I(N__18588));
    LocalMux I__1617 (
            .O(N__18588),
            .I(\nx.n48_adj_692 ));
    CascadeMux I__1616 (
            .O(N__18585),
            .I(\nx.n2908_cascade_ ));
    CascadeMux I__1615 (
            .O(N__18582),
            .I(\nx.n3007_cascade_ ));
    CascadeMux I__1614 (
            .O(N__18579),
            .I(\nx.n3106_cascade_ ));
    InMux I__1613 (
            .O(N__18576),
            .I(N__18573));
    LocalMux I__1612 (
            .O(N__18573),
            .I(\nx.n19_adj_698 ));
    CascadeMux I__1611 (
            .O(N__18570),
            .I(\nx.n3105_cascade_ ));
    InMux I__1610 (
            .O(N__18567),
            .I(N__18564));
    LocalMux I__1609 (
            .O(N__18564),
            .I(\nx.n13271 ));
    CascadeMux I__1608 (
            .O(N__18561),
            .I(\nx.n12369_cascade_ ));
    InMux I__1607 (
            .O(N__18558),
            .I(N__18552));
    InMux I__1606 (
            .O(N__18557),
            .I(N__18552));
    LocalMux I__1605 (
            .O(N__18552),
            .I(neo_pixel_transmitter_t0_15));
    InMux I__1604 (
            .O(N__18549),
            .I(N__18543));
    InMux I__1603 (
            .O(N__18548),
            .I(N__18543));
    LocalMux I__1602 (
            .O(N__18543),
            .I(neo_pixel_transmitter_t0_8));
    CascadeMux I__1601 (
            .O(N__18540),
            .I(\nx.n9700_cascade_ ));
    InMux I__1600 (
            .O(N__18537),
            .I(N__18534));
    LocalMux I__1599 (
            .O(N__18534),
            .I(N__18531));
    Odrv4 I__1598 (
            .O(N__18531),
            .I(\nx.n7131 ));
    CascadeMux I__1597 (
            .O(N__18528),
            .I(\nx.n12117_cascade_ ));
    CascadeMux I__1596 (
            .O(N__18525),
            .I(n7239_cascade_));
    InMux I__1595 (
            .O(N__18522),
            .I(N__18515));
    InMux I__1594 (
            .O(N__18521),
            .I(N__18515));
    InMux I__1593 (
            .O(N__18520),
            .I(N__18512));
    LocalMux I__1592 (
            .O(N__18515),
            .I(N__18509));
    LocalMux I__1591 (
            .O(N__18512),
            .I(\nx.n9700 ));
    Odrv4 I__1590 (
            .O(N__18509),
            .I(\nx.n9700 ));
    InMux I__1589 (
            .O(N__18504),
            .I(N__18498));
    InMux I__1588 (
            .O(N__18503),
            .I(N__18498));
    LocalMux I__1587 (
            .O(N__18498),
            .I(\nx.n9702 ));
    InMux I__1586 (
            .O(N__18495),
            .I(N__18492));
    LocalMux I__1585 (
            .O(N__18492),
            .I(\nx.n11606 ));
    CascadeMux I__1584 (
            .O(N__18489),
            .I(N__18485));
    InMux I__1583 (
            .O(N__18488),
            .I(N__18482));
    InMux I__1582 (
            .O(N__18485),
            .I(N__18479));
    LocalMux I__1581 (
            .O(N__18482),
            .I(N__18474));
    LocalMux I__1580 (
            .O(N__18479),
            .I(N__18474));
    Odrv12 I__1579 (
            .O(N__18474),
            .I(update_color));
    InMux I__1578 (
            .O(N__18471),
            .I(N__18468));
    LocalMux I__1577 (
            .O(N__18468),
            .I(N__18465));
    Odrv4 I__1576 (
            .O(N__18465),
            .I(\nx.n10_adj_653 ));
    CascadeMux I__1575 (
            .O(N__18462),
            .I(\nx.n7131_cascade_ ));
    CascadeMux I__1574 (
            .O(N__18459),
            .I(\nx.n13263_cascade_ ));
    CascadeMux I__1573 (
            .O(N__18456),
            .I(\nx.n7120_cascade_ ));
    CascadeMux I__1572 (
            .O(N__18453),
            .I(\nx.n13262_cascade_ ));
    InMux I__1571 (
            .O(N__18450),
            .I(N__18447));
    LocalMux I__1570 (
            .O(N__18447),
            .I(\nx.n3739 ));
    CascadeMux I__1569 (
            .O(N__18444),
            .I(\nx.n3739_cascade_ ));
    InMux I__1568 (
            .O(N__18441),
            .I(N__18435));
    InMux I__1567 (
            .O(N__18440),
            .I(N__18435));
    LocalMux I__1566 (
            .O(N__18435),
            .I(N__18429));
    InMux I__1565 (
            .O(N__18434),
            .I(N__18424));
    InMux I__1564 (
            .O(N__18433),
            .I(N__18424));
    InMux I__1563 (
            .O(N__18432),
            .I(N__18421));
    Odrv4 I__1562 (
            .O(N__18429),
            .I(\nx.n7120 ));
    LocalMux I__1561 (
            .O(N__18424),
            .I(\nx.n7120 ));
    LocalMux I__1560 (
            .O(N__18421),
            .I(\nx.n7120 ));
    IoInMux I__1559 (
            .O(N__18414),
            .I(N__18411));
    LocalMux I__1558 (
            .O(N__18411),
            .I(NEOPXL_c));
    CascadeMux I__1557 (
            .O(N__18408),
            .I(\nx.n13325_cascade_ ));
    CascadeMux I__1556 (
            .O(N__18405),
            .I(\nx.n11535_cascade_ ));
    CascadeMux I__1555 (
            .O(N__18402),
            .I(\nx.n11672_cascade_ ));
    InMux I__1554 (
            .O(N__18399),
            .I(N__18396));
    LocalMux I__1553 (
            .O(N__18396),
            .I(\nx.n13326 ));
    CEMux I__1552 (
            .O(N__18393),
            .I(N__18390));
    LocalMux I__1551 (
            .O(N__18390),
            .I(N__18387));
    Odrv12 I__1550 (
            .O(N__18387),
            .I(\nx.n11692 ));
    SRMux I__1549 (
            .O(N__18384),
            .I(N__18381));
    LocalMux I__1548 (
            .O(N__18381),
            .I(N__18378));
    Span4Mux_s1_h I__1547 (
            .O(N__18378),
            .I(N__18375));
    Odrv4 I__1546 (
            .O(N__18375),
            .I(\nx.n12204 ));
    CascadeMux I__1545 (
            .O(N__18372),
            .I(\nx.n11696_cascade_ ));
    IoInMux I__1544 (
            .O(N__18369),
            .I(N__18366));
    LocalMux I__1543 (
            .O(N__18366),
            .I(N__18363));
    IoSpan4Mux I__1542 (
            .O(N__18363),
            .I(N__18360));
    IoSpan4Mux I__1541 (
            .O(N__18360),
            .I(N__18357));
    IoSpan4Mux I__1540 (
            .O(N__18357),
            .I(N__18354));
    Odrv4 I__1539 (
            .O(N__18354),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_3_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_21_0_));
    defparam IN_MUX_bfv_3_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_22_0_ (
            .carryinitin(\nx.n10429 ),
            .carryinitout(bfn_3_22_0_));
    defparam IN_MUX_bfv_3_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_23_0_ (
            .carryinitin(\nx.n10436_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_3_23_0_));
    defparam IN_MUX_bfv_3_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_24_0_ (
            .carryinitin(\nx.n10442_THRU_CRY_1_THRU_CO ),
            .carryinitout(bfn_3_24_0_));
    defparam IN_MUX_bfv_3_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_25_0_ (
            .carryinitin(\nx.n10448_THRU_CRY_1_THRU_CO ),
            .carryinitout(bfn_3_25_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(\nx.n10486 ),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(\nx.n10494 ),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\nx.n10502 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_2_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_31_0_));
    defparam IN_MUX_bfv_2_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_32_0_ (
            .carryinitin(\nx.n10580 ),
            .carryinitout(bfn_2_32_0_));
    defparam IN_MUX_bfv_1_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_31_0_));
    defparam IN_MUX_bfv_1_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_32_0_ (
            .carryinitin(\nx.n10460 ),
            .carryinitout(bfn_1_32_0_));
    defparam IN_MUX_bfv_2_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_29_0_));
    defparam IN_MUX_bfv_5_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_26_0_));
    defparam IN_MUX_bfv_6_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_28_0_));
    defparam IN_MUX_bfv_1_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_26_0_));
    defparam IN_MUX_bfv_1_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_27_0_ (
            .carryinitin(\nx.n10895 ),
            .carryinitout(bfn_1_27_0_));
    defparam IN_MUX_bfv_1_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_28_0_ (
            .carryinitin(\nx.n10903 ),
            .carryinitout(bfn_1_28_0_));
    defparam IN_MUX_bfv_1_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_29_0_ (
            .carryinitin(\nx.n10911 ),
            .carryinitout(bfn_1_29_0_));
    defparam IN_MUX_bfv_3_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_26_0_));
    defparam IN_MUX_bfv_3_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_27_0_ (
            .carryinitin(\nx.n10869 ),
            .carryinitout(bfn_3_27_0_));
    defparam IN_MUX_bfv_3_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_28_0_ (
            .carryinitin(\nx.n10877 ),
            .carryinitout(bfn_3_28_0_));
    defparam IN_MUX_bfv_3_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_29_0_ (
            .carryinitin(\nx.n10885 ),
            .carryinitout(bfn_3_29_0_));
    defparam IN_MUX_bfv_5_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_22_0_));
    defparam IN_MUX_bfv_5_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_23_0_ (
            .carryinitin(\nx.n10844 ),
            .carryinitout(bfn_5_23_0_));
    defparam IN_MUX_bfv_5_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_24_0_ (
            .carryinitin(\nx.n10852 ),
            .carryinitout(bfn_5_24_0_));
    defparam IN_MUX_bfv_5_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_25_0_ (
            .carryinitin(\nx.n10860 ),
            .carryinitout(bfn_5_25_0_));
    defparam IN_MUX_bfv_6_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_21_0_));
    defparam IN_MUX_bfv_6_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_22_0_ (
            .carryinitin(\nx.n10820 ),
            .carryinitout(bfn_6_22_0_));
    defparam IN_MUX_bfv_6_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_23_0_ (
            .carryinitin(\nx.n10828 ),
            .carryinitout(bfn_6_23_0_));
    defparam IN_MUX_bfv_6_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_24_0_ (
            .carryinitin(\nx.n10836 ),
            .carryinitout(bfn_6_24_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\nx.n10797 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(\nx.n10805 ),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\nx.n10775 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\nx.n10783 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(\nx.n10754 ),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(\nx.n10762 ),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\nx.n10734 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(\nx.n10742 ),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\nx.n10715 ),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(\nx.n10723 ),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(\nx.n10697 ),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\nx.n10705 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(\nx.n10680 ),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_11_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_25_0_ (
            .carryinitin(\nx.n10688 ),
            .carryinitout(bfn_11_25_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\nx.n10664 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(\nx.n10672 ),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_7_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_25_0_));
    defparam IN_MUX_bfv_7_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_26_0_ (
            .carryinitin(\nx.n10649 ),
            .carryinitout(bfn_7_26_0_));
    defparam IN_MUX_bfv_10_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_28_0_));
    defparam IN_MUX_bfv_10_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_29_0_ (
            .carryinitin(\nx.n10622 ),
            .carryinitout(bfn_10_29_0_));
    defparam IN_MUX_bfv_7_30_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_30_0_));
    defparam IN_MUX_bfv_7_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_31_0_ (
            .carryinitin(\nx.n10610 ),
            .carryinitout(bfn_7_31_0_));
    defparam IN_MUX_bfv_6_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_31_0_));
    defparam IN_MUX_bfv_6_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_32_0_ (
            .carryinitin(\nx.n10599 ),
            .carryinitout(bfn_6_32_0_));
    defparam IN_MUX_bfv_3_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_31_0_));
    defparam IN_MUX_bfv_3_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_32_0_ (
            .carryinitin(\nx.n10589 ),
            .carryinitout(bfn_3_32_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\nx.n10635 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_4_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_27_0_));
    defparam IN_MUX_bfv_4_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_28_0_ (
            .carryinitin(\nx.n10398 ),
            .carryinitout(bfn_4_28_0_));
    defparam IN_MUX_bfv_4_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_29_0_ (
            .carryinitin(\nx.n10406 ),
            .carryinitout(bfn_4_29_0_));
    defparam IN_MUX_bfv_4_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_30_0_ (
            .carryinitin(\nx.n10414 ),
            .carryinitout(bfn_4_30_0_));
    defparam IN_MUX_bfv_12_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_26_0_));
    defparam IN_MUX_bfv_12_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_27_0_ (
            .carryinitin(n10524),
            .carryinitout(bfn_12_27_0_));
    defparam IN_MUX_bfv_12_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_28_0_ (
            .carryinitin(n10532),
            .carryinitout(bfn_12_28_0_));
    defparam IN_MUX_bfv_12_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_29_0_ (
            .carryinitin(n10540),
            .carryinitout(bfn_12_29_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_15_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_27_0_ (
            .carryinitin(n10555),
            .carryinitout(bfn_15_27_0_));
    defparam IN_MUX_bfv_15_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_28_0_ (
            .carryinitin(n10563),
            .carryinitout(bfn_15_28_0_));
    defparam IN_MUX_bfv_15_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_29_0_ (
            .carryinitin(n10571),
            .carryinitout(bfn_15_29_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_17_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18369),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \nx.one_wire_108_LC_1_16_0 .C_ON=1'b0;
    defparam \nx.one_wire_108_LC_1_16_0 .SEQ_MODE=4'b1000;
    defparam \nx.one_wire_108_LC_1_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.one_wire_108_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19281),
            .lcout(NEOPXL_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48384),
            .ce(N__18393),
            .sr(N__18384));
    defparam \nx.i9488_4_lut_LC_1_17_0 .C_ON=1'b0;
    defparam \nx.i9488_4_lut_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.i9488_4_lut_LC_1_17_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \nx.i9488_4_lut_LC_1_17_0  (
            .in0(N__19265),
            .in1(N__19388),
            .in2(N__19604),
            .in3(N__19182),
            .lcout(),
            .ltout(\nx.n13325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9478_3_lut_4_lut_LC_1_17_1 .C_ON=1'b0;
    defparam \nx.i9478_3_lut_4_lut_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9478_3_lut_4_lut_LC_1_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9478_3_lut_4_lut_LC_1_17_1  (
            .in0(N__19149),
            .in1(N__18440),
            .in2(N__18408),
            .in3(N__19511),
            .lcout(\nx.n13326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7775_2_lut_LC_1_17_2 .C_ON=1'b0;
    defparam \nx.i7775_2_lut_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \nx.i7775_2_lut_LC_1_17_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \nx.i7775_2_lut_LC_1_17_2  (
            .in0(N__18441),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19150),
            .lcout(),
            .ltout(\nx.n11535_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i53_4_lut_LC_1_17_3 .C_ON=1'b0;
    defparam \nx.i53_4_lut_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.i53_4_lut_LC_1_17_3 .LUT_INIT=16'b1111111000110010;
    LogicCell40 \nx.i53_4_lut_LC_1_17_3  (
            .in0(N__19389),
            .in1(N__19512),
            .in2(N__18405),
            .in3(N__18521),
            .lcout(),
            .ltout(\nx.n11672_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i52_4_lut_LC_1_17_4 .C_ON=1'b0;
    defparam \nx.i52_4_lut_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \nx.i52_4_lut_LC_1_17_4 .LUT_INIT=16'b0000000111101111;
    LogicCell40 \nx.i52_4_lut_LC_1_17_4  (
            .in0(N__19603),
            .in1(N__19267),
            .in2(N__18402),
            .in3(N__18399),
            .lcout(\nx.n11692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_4_lut_4_lut_LC_1_17_6 .C_ON=1'b0;
    defparam \nx.i3_4_lut_4_lut_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.i3_4_lut_4_lut_LC_1_17_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \nx.i3_4_lut_4_lut_LC_1_17_6  (
            .in0(N__18522),
            .in1(N__19514),
            .in2(N__19605),
            .in3(N__19266),
            .lcout(\nx.n12204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i22_4_lut_adj_157_LC_1_18_1 .C_ON=1'b0;
    defparam \nx.i22_4_lut_adj_157_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.i22_4_lut_adj_157_LC_1_18_1 .LUT_INIT=16'b1011100011100010;
    LogicCell40 \nx.i22_4_lut_adj_157_LC_1_18_1  (
            .in0(N__19387),
            .in1(N__19263),
            .in2(N__19181),
            .in3(N__19595),
            .lcout(),
            .ltout(\nx.n11696_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7914_4_lut_LC_1_18_2 .C_ON=1'b0;
    defparam \nx.i7914_4_lut_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.i7914_4_lut_LC_1_18_2 .LUT_INIT=16'b1010101010101011;
    LogicCell40 \nx.i7914_4_lut_LC_1_18_2  (
            .in0(N__19513),
            .in1(N__18434),
            .in2(N__18372),
            .in3(N__19145),
            .lcout(n11683),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.equal_607_i8_2_lut_LC_1_18_5 .C_ON=1'b0;
    defparam \nx.equal_607_i8_2_lut_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.equal_607_i8_2_lut_LC_1_18_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \nx.equal_607_i8_2_lut_LC_1_18_5  (
            .in0(N__19144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19262),
            .lcout(\nx.n7131 ),
            .ltout(\nx.n7131_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9439_3_lut_LC_1_18_6 .C_ON=1'b0;
    defparam \nx.i9439_3_lut_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9439_3_lut_LC_1_18_6 .LUT_INIT=16'b1111000011110011;
    LogicCell40 \nx.i9439_3_lut_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__18433),
            .in2(N__18462),
            .in3(N__19174),
            .lcout(),
            .ltout(\nx.n13263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9551_4_lut_4_lut_LC_1_18_7 .C_ON=1'b0;
    defparam \nx.i9551_4_lut_4_lut_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.i9551_4_lut_4_lut_LC_1_18_7 .LUT_INIT=16'b0000000111001101;
    LogicCell40 \nx.i9551_4_lut_4_lut_LC_1_18_7  (
            .in0(N__19510),
            .in1(N__19594),
            .in2(N__18459),
            .in3(N__18450),
            .lcout(\nx.n7230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_153_LC_1_19_1 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_153_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_153_LC_1_19_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_153_LC_1_19_1  (
            .in0(N__21064),
            .in1(N__19017),
            .in2(N__21134),
            .in3(N__21709),
            .lcout(\nx.n7120 ),
            .ltout(\nx.n7120_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9469_3_lut_4_lut_LC_1_19_2 .C_ON=1'b0;
    defparam \nx.i9469_3_lut_4_lut_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9469_3_lut_4_lut_LC_1_19_2 .LUT_INIT=16'b1011101110111111;
    LogicCell40 \nx.i9469_3_lut_4_lut_LC_1_19_2  (
            .in0(N__19143),
            .in1(N__19264),
            .in2(N__18456),
            .in3(N__19378),
            .lcout(),
            .ltout(\nx.n13262_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1393_4_lut_LC_1_19_3 .C_ON=1'b0;
    defparam \nx.i1393_4_lut_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1393_4_lut_LC_1_19_3 .LUT_INIT=16'b0111011111110000;
    LogicCell40 \nx.i1393_4_lut_LC_1_19_3  (
            .in0(N__20171),
            .in1(N__18488),
            .in2(N__18453),
            .in3(N__19480),
            .lcout(\nx.n3739 ),
            .ltout(\nx.n3739_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_3_lut_adj_144_LC_1_19_4 .C_ON=1'b0;
    defparam \nx.i5_3_lut_adj_144_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.i5_3_lut_adj_144_LC_1_19_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \nx.i5_3_lut_adj_144_LC_1_19_4  (
            .in0(N__19586),
            .in1(_gnd_net_),
            .in2(N__18444),
            .in3(N__18471),
            .lcout(\nx.n7411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam update_color_195_LC_1_19_5.C_ON=1'b0;
    defparam update_color_195_LC_1_19_5.SEQ_MODE=4'b1001;
    defparam update_color_195_LC_1_19_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 update_color_195_LC_1_19_5 (
            .in0(N__25014),
            .in1(N__19323),
            .in2(N__19203),
            .in3(N__19305),
            .lcout(update_color),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48386),
            .ce(),
            .sr(N__47115));
    defparam \nx.i7796_4_lut_LC_1_19_6 .C_ON=1'b0;
    defparam \nx.i7796_4_lut_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.i7796_4_lut_LC_1_19_6 .LUT_INIT=16'b1111111111001010;
    LogicCell40 \nx.i7796_4_lut_LC_1_19_6  (
            .in0(N__19173),
            .in1(N__19377),
            .in2(N__19596),
            .in3(N__18432),
            .lcout(\nx.n9702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6476_4_lut_LC_1_20_0 .C_ON=1'b0;
    defparam \nx.i6476_4_lut_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.i6476_4_lut_LC_1_20_0 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \nx.i6476_4_lut_LC_1_20_0  (
            .in0(N__21066),
            .in1(N__21167),
            .in2(N__21135),
            .in3(N__21711),
            .lcout(\nx.n9700 ),
            .ltout(\nx.n9700_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_3_lut_4_lut_LC_1_20_1 .C_ON=1'b0;
    defparam \nx.i1_3_lut_4_lut_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_3_lut_4_lut_LC_1_20_1 .LUT_INIT=16'b1101110011111111;
    LogicCell40 \nx.i1_3_lut_4_lut_LC_1_20_1  (
            .in0(N__19282),
            .in1(N__19580),
            .in2(N__18540),
            .in3(N__19495),
            .lcout(),
            .ltout(\nx.n12117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_131_LC_1_20_2 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_131_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_131_LC_1_20_2 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \nx.i1_4_lut_adj_131_LC_1_20_2  (
            .in0(N__19496),
            .in1(N__18537),
            .in2(N__18528),
            .in3(N__18503),
            .lcout(n7239),
            .ltout(n7239_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.state_i1_LC_1_20_3 .C_ON=1'b0;
    defparam \nx.state_i1_LC_1_20_3 .SEQ_MODE=4'b1000;
    defparam \nx.state_i1_LC_1_20_3 .LUT_INIT=16'b1011111111110000;
    LogicCell40 \nx.state_i1_LC_1_20_3  (
            .in0(N__20172),
            .in1(N__19581),
            .in2(N__18525),
            .in3(N__19500),
            .lcout(state_1_adj_726),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48389),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_145_LC_1_20_4 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_145_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_145_LC_1_20_4 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \nx.i15_4_lut_adj_145_LC_1_20_4  (
            .in0(N__18567),
            .in1(N__18520),
            .in2(N__19515),
            .in3(N__18495),
            .lcout(\nx.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i5_LC_1_20_5.C_ON=1'b0;
    defparam neopxl_color_prev_i5_LC_1_20_5.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i5_LC_1_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 neopxl_color_prev_i5_LC_1_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39795),
            .lcout(neopxl_color_prev_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48389),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7843_3_lut_LC_1_20_7 .C_ON=1'b0;
    defparam \nx.i7843_3_lut_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.i7843_3_lut_LC_1_20_7 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \nx.i7843_3_lut_LC_1_20_7  (
            .in0(N__18504),
            .in1(_gnd_net_),
            .in2(N__19287),
            .in3(N__19154),
            .lcout(\nx.n11606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.state_i0_LC_1_21_0 .C_ON=1'b0;
    defparam \nx.state_i0_LC_1_21_0 .SEQ_MODE=4'b1001;
    defparam \nx.state_i0_LC_1_21_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \nx.state_i0_LC_1_21_0  (
            .in0(N__23913),
            .in1(N__20164),
            .in2(N__19668),
            .in3(N__19395),
            .lcout(state_0_adj_727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48395),
            .ce(N__19431),
            .sr(N__19419));
    defparam \nx.i4_4_lut_4_lut_LC_1_21_2 .C_ON=1'b0;
    defparam \nx.i4_4_lut_4_lut_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i4_4_lut_4_lut_LC_1_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \nx.i4_4_lut_4_lut_LC_1_21_2  (
            .in0(N__19479),
            .in1(N__19564),
            .in2(N__18489),
            .in3(N__20163),
            .lcout(\nx.n10_adj_653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9438_2_lut_LC_1_21_3 .C_ON=1'b0;
    defparam \nx.i9438_2_lut_LC_1_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9438_2_lut_LC_1_21_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \nx.i9438_2_lut_LC_1_21_3  (
            .in0(N__19565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19286),
            .lcout(\nx.n13271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_128_LC_1_22_0 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_128_LC_1_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_128_LC_1_22_0 .LUT_INIT=16'b1111111111100100;
    LogicCell40 \nx.i1_4_lut_adj_128_LC_1_22_0  (
            .in0(N__24213),
            .in1(N__19727),
            .in2(N__18849),
            .in3(N__24072),
            .lcout(),
            .ltout(\nx.n12369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_129_LC_1_22_1 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_129_LC_1_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_129_LC_1_22_1 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \nx.i1_4_lut_adj_129_LC_1_22_1  (
            .in0(N__19748),
            .in1(N__18831),
            .in2(N__18561),
            .in3(N__24214),
            .lcout(\nx.n12371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i9_1_lut_LC_1_22_2 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i9_1_lut_LC_1_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i9_1_lut_LC_1_22_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \nx.sub_14_inv_0_i9_1_lut_LC_1_22_2  (
            .in0(N__18548),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\nx.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9309_3_lut_LC_1_22_3 .C_ON=1'b0;
    defparam \nx.i9309_3_lut_LC_1_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9309_3_lut_LC_1_22_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.i9309_3_lut_LC_1_22_3  (
            .in0(N__40756),
            .in1(N__37434),
            .in2(_gnd_net_),
            .in3(N__23990),
            .lcout(\nx.n13156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i15_LC_1_22_4 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i15_LC_1_22_4 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i15_LC_1_22_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i15_LC_1_22_4  (
            .in0(N__18558),
            .in1(N__21399),
            .in2(_gnd_net_),
            .in3(N__28864),
            .lcout(neo_pixel_transmitter_t0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i16_1_lut_LC_1_22_5 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i16_1_lut_LC_1_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i16_1_lut_LC_1_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i16_1_lut_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18557),
            .lcout(\nx.n18_adj_623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i8_LC_1_22_6 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i8_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i8_LC_1_22_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i8_LC_1_22_6  (
            .in0(N__18549),
            .in1(N__28863),
            .in2(_gnd_net_),
            .in3(N__21198),
            .lcout(neo_pixel_transmitter_t0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i5_LC_1_22_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i5_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i5_LC_1_22_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i5_LC_1_22_7  (
            .in0(N__28862),
            .in1(N__20772),
            .in2(_gnd_net_),
            .in3(N__19064),
            .lcout(neo_pixel_transmitter_t0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48401),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2090_3_lut_LC_1_23_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2090_3_lut_LC_1_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2090_3_lut_LC_1_23_0 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i2090_3_lut_LC_1_23_0  (
            .in0(_gnd_net_),
            .in1(N__27400),
            .in2(N__23354),
            .in3(N__21963),
            .lcout(\nx.n3095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1967_3_lut_LC_1_23_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1967_3_lut_LC_1_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1967_3_lut_LC_1_23_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1967_3_lut_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(N__30257),
            .in2(N__27027),
            .in3(N__27003),
            .lcout(\nx.n2908 ),
            .ltout(\nx.n2908_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2034_3_lut_LC_1_23_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2034_3_lut_LC_1_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2034_3_lut_LC_1_23_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2034_3_lut_LC_1_23_3  (
            .in0(_gnd_net_),
            .in1(N__25398),
            .in2(N__18585),
            .in3(N__31874),
            .lcout(\nx.n3007 ),
            .ltout(\nx.n3007_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2101_3_lut_LC_1_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2101_3_lut_LC_1_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2101_3_lut_LC_1_23_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i2101_3_lut_LC_1_23_4  (
            .in0(N__21855),
            .in1(_gnd_net_),
            .in2(N__18582),
            .in3(N__27401),
            .lcout(\nx.n3106 ),
            .ltout(\nx.n3106_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_112_LC_1_23_5 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_112_LC_1_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_112_LC_1_23_5 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \nx.i1_4_lut_adj_112_LC_1_23_5  (
            .in0(N__18678),
            .in1(N__18576),
            .in2(N__18579),
            .in3(N__24209),
            .lcout(\nx.n12335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2147_3_lut_LC_1_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2147_3_lut_LC_1_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2147_3_lut_LC_1_23_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2147_3_lut_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(N__18897),
            .in2(N__24235),
            .in3(N__19694),
            .lcout(\nx.n59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2167_3_lut_LC_1_24_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2167_3_lut_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2167_3_lut_LC_1_24_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2167_3_lut_LC_1_24_0  (
            .in0(_gnd_net_),
            .in1(N__18645),
            .in2(N__18665),
            .in3(N__24167),
            .lcout(\nx.n19_adj_698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2100_3_lut_LC_1_24_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2100_3_lut_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2100_3_lut_LC_1_24_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2100_3_lut_LC_1_24_1  (
            .in0(_gnd_net_),
            .in1(N__23192),
            .in2(N__21840),
            .in3(N__27387),
            .lcout(\nx.n3105 ),
            .ltout(\nx.n3105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_102_LC_1_24_2 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_102_LC_1_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_102_LC_1_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_102_LC_1_24_2  (
            .in0(N__18770),
            .in1(N__20101),
            .in2(N__18570),
            .in3(N__20062),
            .lcout(\nx.n46_adj_688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2097_3_lut_LC_1_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2097_3_lut_LC_1_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2097_3_lut_LC_1_24_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2097_3_lut_LC_1_24_3  (
            .in0(_gnd_net_),
            .in1(N__31733),
            .in2(N__22125),
            .in3(N__27388),
            .lcout(\nx.n3102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2095_3_lut_LC_1_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2095_3_lut_LC_1_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2095_3_lut_LC_1_24_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i2095_3_lut_LC_1_24_4  (
            .in0(N__22085),
            .in1(_gnd_net_),
            .in2(N__27436),
            .in3(N__22065),
            .lcout(\nx.n3100 ),
            .ltout(\nx.n3100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2162_3_lut_LC_1_24_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2162_3_lut_LC_1_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2162_3_lut_LC_1_24_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i2162_3_lut_LC_1_24_5  (
            .in0(N__24168),
            .in1(_gnd_net_),
            .in2(N__18621),
            .in3(N__18759),
            .lcout(),
            .ltout(\nx.n29_adj_697_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_114_LC_1_24_6 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_114_LC_1_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_114_LC_1_24_6 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \nx.i1_4_lut_adj_114_LC_1_24_6  (
            .in0(N__19823),
            .in1(N__18714),
            .in2(N__18618),
            .in3(N__24169),
            .lcout(),
            .ltout(\nx.n12331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_119_LC_1_24_7 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_119_LC_1_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_119_LC_1_24_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_119_LC_1_24_7  (
            .in0(N__19830),
            .in1(N__18603),
            .in2(N__18615),
            .in3(N__18612),
            .lcout(\nx.n12349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i21_4_lut_adj_107_LC_1_25_0 .C_ON=1'b0;
    defparam \nx.i21_4_lut_adj_107_LC_1_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.i21_4_lut_adj_107_LC_1_25_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i21_4_lut_adj_107_LC_1_25_0  (
            .in0(N__20221),
            .in1(N__20142),
            .in2(N__22281),
            .in3(N__19674),
            .lcout(\nx.n48_adj_692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2158_3_lut_LC_1_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2158_3_lut_LC_1_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2158_3_lut_LC_1_25_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i2158_3_lut_LC_1_25_1  (
            .in0(N__19793),
            .in1(_gnd_net_),
            .in2(N__18738),
            .in3(N__24170),
            .lcout(),
            .ltout(\nx.n37_adj_695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_111_LC_1_25_2 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_111_LC_1_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_111_LC_1_25_2 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \nx.i1_4_lut_adj_111_LC_1_25_2  (
            .in0(N__24171),
            .in1(N__18815),
            .in2(N__18606),
            .in3(N__18792),
            .lcout(\nx.n12333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_3_lut_adj_105_LC_1_25_3 .C_ON=1'b0;
    defparam \nx.i4_3_lut_adj_105_LC_1_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.i4_3_lut_adj_105_LC_1_25_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \nx.i4_3_lut_adj_105_LC_1_25_3  (
            .in0(N__24375),
            .in1(N__18811),
            .in2(_gnd_net_),
            .in3(N__19822),
            .lcout(),
            .ltout(\nx.n31_adj_691_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i22_4_lut_adj_108_LC_1_25_4 .C_ON=1'b0;
    defparam \nx.i22_4_lut_adj_108_LC_1_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.i22_4_lut_adj_108_LC_1_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i22_4_lut_adj_108_LC_1_25_4  (
            .in0(N__18693),
            .in1(N__19915),
            .in2(N__18597),
            .in3(N__23748),
            .lcout(),
            .ltout(\nx.n49_adj_693_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i26_4_lut_LC_1_25_5 .C_ON=1'b0;
    defparam \nx.i26_4_lut_LC_1_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.i26_4_lut_LC_1_25_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i26_4_lut_LC_1_25_5  (
            .in0(N__19773),
            .in1(N__25749),
            .in2(N__18594),
            .in3(N__18591),
            .lcout(\nx.n3116 ),
            .ltout(\nx.n3116_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2165_3_lut_LC_1_25_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2165_3_lut_LC_1_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2165_3_lut_LC_1_25_6 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \nx.mod_5_i2165_3_lut_LC_1_25_6  (
            .in0(N__18630),
            .in1(N__19916),
            .in2(N__18720),
            .in3(_gnd_net_),
            .lcout(\nx.n23_adj_700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_2_lut_LC_1_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_2_lut_LC_1_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_2_lut_LC_1_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_2_lut_LC_1_26_0  (
            .in0(_gnd_net_),
            .in1(N__24369),
            .in2(_gnd_net_),
            .in3(N__18717),
            .lcout(\nx.n3177 ),
            .ltout(),
            .carryin(bfn_1_26_0_),
            .carryout(\nx.n10888 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_3_lut_LC_1_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_3_lut_LC_1_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_3_lut_LC_1_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_3_lut_LC_1_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19824),
            .in3(N__18702),
            .lcout(\nx.n3176 ),
            .ltout(),
            .carryin(\nx.n10888 ),
            .carryout(\nx.n10889 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_4_lut_LC_1_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_4_lut_LC_1_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_4_lut_LC_1_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_4_lut_LC_1_26_2  (
            .in0(_gnd_net_),
            .in1(N__44706),
            .in2(N__20003),
            .in3(N__18699),
            .lcout(\nx.n3175 ),
            .ltout(),
            .carryin(\nx.n10889 ),
            .carryout(\nx.n10890 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_5_lut_LC_1_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_5_lut_LC_1_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_5_lut_LC_1_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_5_lut_LC_1_26_3  (
            .in0(_gnd_net_),
            .in1(N__20102),
            .in2(N__45093),
            .in3(N__18696),
            .lcout(\nx.n3174 ),
            .ltout(),
            .carryin(\nx.n10890 ),
            .carryout(\nx.n10891 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_6_lut_LC_1_26_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_6_lut_LC_1_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_6_lut_LC_1_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_6_lut_LC_1_26_4  (
            .in0(_gnd_net_),
            .in1(N__18692),
            .in2(N__45094),
            .in3(N__18669),
            .lcout(\nx.n3173 ),
            .ltout(),
            .carryin(\nx.n10891 ),
            .carryout(\nx.n10892 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_7_lut_LC_1_26_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_7_lut_LC_1_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_7_lut_LC_1_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_7_lut_LC_1_26_5  (
            .in0(_gnd_net_),
            .in1(N__44714),
            .in2(N__18666),
            .in3(N__18636),
            .lcout(\nx.n3172 ),
            .ltout(),
            .carryin(\nx.n10892 ),
            .carryout(\nx.n10893 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_8_lut_LC_1_26_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_8_lut_LC_1_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_8_lut_LC_1_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_8_lut_LC_1_26_6  (
            .in0(_gnd_net_),
            .in1(N__44710),
            .in2(N__23777),
            .in3(N__18633),
            .lcout(\nx.n3171 ),
            .ltout(),
            .carryin(\nx.n10893 ),
            .carryout(\nx.n10894 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_9_lut_LC_1_26_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_9_lut_LC_1_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_9_lut_LC_1_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_9_lut_LC_1_26_7  (
            .in0(_gnd_net_),
            .in1(N__44715),
            .in2(N__19920),
            .in3(N__18624),
            .lcout(\nx.n3170 ),
            .ltout(),
            .carryin(\nx.n10894 ),
            .carryout(\nx.n10895 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_10_lut_LC_1_27_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_10_lut_LC_1_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_10_lut_LC_1_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_10_lut_LC_1_27_0  (
            .in0(_gnd_net_),
            .in1(N__44665),
            .in2(N__18816),
            .in3(N__18783),
            .lcout(\nx.n3169 ),
            .ltout(),
            .carryin(bfn_1_27_0_),
            .carryout(\nx.n10896 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_11_lut_LC_1_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_11_lut_LC_1_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_11_lut_LC_1_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_11_lut_LC_1_27_1  (
            .in0(_gnd_net_),
            .in1(N__45671),
            .in2(N__19857),
            .in3(N__18780),
            .lcout(\nx.n3168 ),
            .ltout(),
            .carryin(\nx.n10896 ),
            .carryout(\nx.n10897 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_12_lut_LC_1_27_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_12_lut_LC_1_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_12_lut_LC_1_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_12_lut_LC_1_27_2  (
            .in0(_gnd_net_),
            .in1(N__44666),
            .in2(N__18777),
            .in3(N__18750),
            .lcout(\nx.n3167 ),
            .ltout(),
            .carryin(\nx.n10897 ),
            .carryout(\nx.n10898 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_13_lut_LC_1_27_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_13_lut_LC_1_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_13_lut_LC_1_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_13_lut_LC_1_27_3  (
            .in0(_gnd_net_),
            .in1(N__45672),
            .in2(N__20223),
            .in3(N__18747),
            .lcout(\nx.n3166 ),
            .ltout(),
            .carryin(\nx.n10898 ),
            .carryout(\nx.n10899 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_14_lut_LC_1_27_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_14_lut_LC_1_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_14_lut_LC_1_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_14_lut_LC_1_27_4  (
            .in0(_gnd_net_),
            .in1(N__19973),
            .in2(N__45755),
            .in3(N__18744),
            .lcout(\nx.n3165 ),
            .ltout(),
            .carryin(\nx.n10899 ),
            .carryout(\nx.n10900 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_15_lut_LC_1_27_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_15_lut_LC_1_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_15_lut_LC_1_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_15_lut_LC_1_27_5  (
            .in0(_gnd_net_),
            .in1(N__19899),
            .in2(N__45029),
            .in3(N__18741),
            .lcout(\nx.n3164 ),
            .ltout(),
            .carryin(\nx.n10900 ),
            .carryout(\nx.n10901 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_16_lut_LC_1_27_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_16_lut_LC_1_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_16_lut_LC_1_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_16_lut_LC_1_27_6  (
            .in0(_gnd_net_),
            .in1(N__44670),
            .in2(N__19797),
            .in3(N__18726),
            .lcout(\nx.n3163 ),
            .ltout(),
            .carryin(\nx.n10901 ),
            .carryout(\nx.n10902 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_17_lut_LC_1_27_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_17_lut_LC_1_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_17_lut_LC_1_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_17_lut_LC_1_27_7  (
            .in0(_gnd_net_),
            .in1(N__45676),
            .in2(N__20075),
            .in3(N__18723),
            .lcout(\nx.n3162 ),
            .ltout(),
            .carryin(\nx.n10902 ),
            .carryout(\nx.n10903 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_18_lut_LC_1_28_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_18_lut_LC_1_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_18_lut_LC_1_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_18_lut_LC_1_28_0  (
            .in0(_gnd_net_),
            .in1(N__27312),
            .in2(N__45758),
            .in3(N__18870),
            .lcout(\nx.n3161 ),
            .ltout(),
            .carryin(bfn_1_28_0_),
            .carryout(\nx.n10904 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_19_lut_LC_1_28_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_19_lut_LC_1_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_19_lut_LC_1_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_19_lut_LC_1_28_1  (
            .in0(_gnd_net_),
            .in1(N__25737),
            .in2(N__45761),
            .in3(N__18867),
            .lcout(\nx.n3160 ),
            .ltout(),
            .carryin(\nx.n10904 ),
            .carryout(\nx.n10905 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_20_lut_LC_1_28_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_20_lut_LC_1_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_20_lut_LC_1_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_20_lut_LC_1_28_2  (
            .in0(_gnd_net_),
            .in1(N__25812),
            .in2(N__45759),
            .in3(N__18864),
            .lcout(\nx.n3159 ),
            .ltout(),
            .carryin(\nx.n10905 ),
            .carryout(\nx.n10906 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_21_lut_LC_1_28_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_21_lut_LC_1_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_21_lut_LC_1_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_21_lut_LC_1_28_3  (
            .in0(_gnd_net_),
            .in1(N__25783),
            .in2(N__45762),
            .in3(N__18861),
            .lcout(\nx.n3158 ),
            .ltout(),
            .carryin(\nx.n10906 ),
            .carryout(\nx.n10907 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_22_lut_LC_1_28_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_22_lut_LC_1_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_22_lut_LC_1_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_22_lut_LC_1_28_4  (
            .in0(_gnd_net_),
            .in1(N__45720),
            .in2(N__24288),
            .in3(N__18858),
            .lcout(\nx.n3157 ),
            .ltout(),
            .carryin(\nx.n10907 ),
            .carryout(\nx.n10908 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_23_lut_LC_1_28_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_23_lut_LC_1_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_23_lut_LC_1_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_23_lut_LC_1_28_5  (
            .in0(_gnd_net_),
            .in1(N__24015),
            .in2(N__45763),
            .in3(N__18855),
            .lcout(\nx.n3156 ),
            .ltout(),
            .carryin(\nx.n10908 ),
            .carryout(\nx.n10909 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_24_lut_LC_1_28_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_24_lut_LC_1_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_24_lut_LC_1_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_24_lut_LC_1_28_6  (
            .in0(_gnd_net_),
            .in1(N__24105),
            .in2(N__45760),
            .in3(N__18852),
            .lcout(\nx.n3155 ),
            .ltout(),
            .carryin(\nx.n10909 ),
            .carryout(\nx.n10910 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_25_lut_LC_1_28_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_25_lut_LC_1_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_25_lut_LC_1_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_25_lut_LC_1_28_7  (
            .in0(_gnd_net_),
            .in1(N__19728),
            .in2(N__45764),
            .in3(N__18834),
            .lcout(\nx.n3154 ),
            .ltout(),
            .carryin(\nx.n10910 ),
            .carryout(\nx.n10911 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_26_lut_LC_1_29_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_26_lut_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_26_lut_LC_1_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_26_lut_LC_1_29_0  (
            .in0(_gnd_net_),
            .in1(N__19749),
            .in2(N__45625),
            .in3(N__18819),
            .lcout(\nx.n3153 ),
            .ltout(),
            .carryin(bfn_1_29_0_),
            .carryout(\nx.n10912 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_27_lut_LC_1_29_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_27_lut_LC_1_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_27_lut_LC_1_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_27_lut_LC_1_29_1  (
            .in0(_gnd_net_),
            .in1(N__19698),
            .in2(N__45627),
            .in3(N__18888),
            .lcout(\nx.n3152 ),
            .ltout(),
            .carryin(\nx.n10912 ),
            .carryout(\nx.n10913 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_28_lut_LC_1_29_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_28_lut_LC_1_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_28_lut_LC_1_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_28_lut_LC_1_29_2  (
            .in0(_gnd_net_),
            .in1(N__20137),
            .in2(N__45626),
            .in3(N__18885),
            .lcout(\nx.n3151 ),
            .ltout(),
            .carryin(\nx.n10913 ),
            .carryout(\nx.n10914 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_29_lut_LC_1_29_3 .C_ON=1'b0;
    defparam \nx.mod_5_add_2143_29_lut_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_29_lut_LC_1_29_3 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_2143_29_lut_LC_1_29_3  (
            .in0(N__22277),
            .in1(N__45292),
            .in2(N__24246),
            .in3(N__18882),
            .lcout(\nx.n13042 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i744_3_lut_LC_1_29_7 .C_ON=1'b0;
    defparam \nx.mod_5_i744_3_lut_LC_1_29_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i744_3_lut_LC_1_29_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i744_3_lut_LC_1_29_7  (
            .in0(N__25707),
            .in1(N__26231),
            .in2(_gnd_net_),
            .in3(N__26052),
            .lcout(\nx.n1109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_2_lut_adj_30_LC_1_30_0 .C_ON=1'b0;
    defparam \nx.i3_2_lut_adj_30_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \nx.i3_2_lut_adj_30_LC_1_30_0 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i3_2_lut_adj_30_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26351),
            .in3(N__26284),
            .lcout(),
            .ltout(\nx.n10_adj_619_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_4_lut_LC_1_30_1 .C_ON=1'b0;
    defparam \nx.i5_4_lut_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \nx.i5_4_lut_LC_1_30_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \nx.i5_4_lut_LC_1_30_1  (
            .in0(N__20335),
            .in1(N__24460),
            .in2(N__18879),
            .in3(N__26011),
            .lcout(),
            .ltout(\nx.n12_adj_621_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_4_lut_LC_1_30_2 .C_ON=1'b0;
    defparam \nx.i6_4_lut_LC_1_30_2 .SEQ_MODE=4'b0000;
    defparam \nx.i6_4_lut_LC_1_30_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i6_4_lut_LC_1_30_2  (
            .in0(N__25894),
            .in1(N__25976),
            .in2(N__18876),
            .in3(N__25931),
            .lcout(\nx.n1136 ),
            .ltout(\nx.n1136_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i812_3_lut_LC_1_30_3 .C_ON=1'b0;
    defparam \nx.mod_5_i812_3_lut_LC_1_30_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i812_3_lut_LC_1_30_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i812_3_lut_LC_1_30_3  (
            .in0(_gnd_net_),
            .in1(N__20346),
            .in2(N__18873),
            .in3(N__24461),
            .lcout(\nx.n1209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i806_3_lut_LC_1_30_4 .C_ON=1'b0;
    defparam \nx.mod_5_i806_3_lut_LC_1_30_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i806_3_lut_LC_1_30_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i806_3_lut_LC_1_30_4  (
            .in0(_gnd_net_),
            .in1(N__26012),
            .in2(N__20283),
            .in3(N__20424),
            .lcout(\nx.n1203 ),
            .ltout(\nx.n1203_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_4_lut_adj_31_LC_1_30_5 .C_ON=1'b0;
    defparam \nx.i5_4_lut_adj_31_LC_1_30_5 .SEQ_MODE=4'b0000;
    defparam \nx.i5_4_lut_adj_31_LC_1_30_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i5_4_lut_adj_31_LC_1_30_5  (
            .in0(N__20513),
            .in1(N__22396),
            .in2(N__18924),
            .in3(N__20261),
            .lcout(\nx.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i811_3_lut_LC_1_30_6 .C_ON=1'b0;
    defparam \nx.mod_5_i811_3_lut_LC_1_30_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i811_3_lut_LC_1_30_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i811_3_lut_LC_1_30_6  (
            .in0(_gnd_net_),
            .in1(N__20336),
            .in2(N__20319),
            .in3(N__20423),
            .lcout(\nx.n1208 ),
            .ltout(\nx.n1208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_3_lut_LC_1_30_7 .C_ON=1'b0;
    defparam \nx.i3_3_lut_LC_1_30_7 .SEQ_MODE=4'b0000;
    defparam \nx.i3_3_lut_LC_1_30_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i3_3_lut_LC_1_30_7  (
            .in0(_gnd_net_),
            .in1(N__24542),
            .in2(N__18921),
            .in3(N__18967),
            .lcout(\nx.n11_adj_624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_2_lut_LC_1_31_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_2_lut_LC_1_31_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_2_lut_LC_1_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_2_lut_LC_1_31_0  (
            .in0(_gnd_net_),
            .in1(N__24543),
            .in2(_gnd_net_),
            .in3(N__18918),
            .lcout(\nx.n1277 ),
            .ltout(),
            .carryin(bfn_1_31_0_),
            .carryout(\nx.n10453 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_3_lut_LC_1_31_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_3_lut_LC_1_31_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_3_lut_LC_1_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_3_lut_LC_1_31_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18971),
            .in3(N__18915),
            .lcout(\nx.n1276 ),
            .ltout(),
            .carryin(\nx.n10453 ),
            .carryout(\nx.n10454 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_4_lut_LC_1_31_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_4_lut_LC_1_31_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_4_lut_LC_1_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_4_lut_LC_1_31_2  (
            .in0(_gnd_net_),
            .in1(N__45308),
            .in2(N__20448),
            .in3(N__18912),
            .lcout(\nx.n1275 ),
            .ltout(),
            .carryin(\nx.n10454 ),
            .carryout(\nx.n10455 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_5_lut_LC_1_31_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_5_lut_LC_1_31_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_5_lut_LC_1_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_5_lut_LC_1_31_3  (
            .in0(_gnd_net_),
            .in1(N__45311),
            .in2(N__20385),
            .in3(N__18909),
            .lcout(\nx.n1274 ),
            .ltout(),
            .carryin(\nx.n10455 ),
            .carryout(\nx.n10456 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_6_lut_LC_1_31_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_6_lut_LC_1_31_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_6_lut_LC_1_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_6_lut_LC_1_31_4  (
            .in0(_gnd_net_),
            .in1(N__45309),
            .in2(N__20477),
            .in3(N__18906),
            .lcout(\nx.n1273 ),
            .ltout(),
            .carryin(\nx.n10456 ),
            .carryout(\nx.n10457 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_7_lut_LC_1_31_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_7_lut_LC_1_31_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_7_lut_LC_1_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_7_lut_LC_1_31_5  (
            .in0(_gnd_net_),
            .in1(N__45312),
            .in2(N__22403),
            .in3(N__18903),
            .lcout(\nx.n1272 ),
            .ltout(),
            .carryin(\nx.n10457 ),
            .carryout(\nx.n10458 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_8_lut_LC_1_31_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_8_lut_LC_1_31_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_8_lut_LC_1_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_8_lut_LC_1_31_6  (
            .in0(_gnd_net_),
            .in1(N__45310),
            .in2(N__20517),
            .in3(N__18900),
            .lcout(\nx.n1271 ),
            .ltout(),
            .carryin(\nx.n10458 ),
            .carryout(\nx.n10459 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_9_lut_LC_1_31_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_9_lut_LC_1_31_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_9_lut_LC_1_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_9_lut_LC_1_31_7  (
            .in0(_gnd_net_),
            .in1(N__45313),
            .in2(N__19004),
            .in3(N__19011),
            .lcout(\nx.n1270 ),
            .ltout(),
            .carryin(\nx.n10459 ),
            .carryout(\nx.n10460 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_10_lut_LC_1_32_0 .C_ON=1'b0;
    defparam \nx.mod_5_add_870_10_lut_LC_1_32_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_10_lut_LC_1_32_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_870_10_lut_LC_1_32_0  (
            .in0(N__44385),
            .in1(N__20268),
            .in2(N__22378),
            .in3(N__19008),
            .lcout(\nx.n1301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i873_3_lut_LC_1_32_2 .C_ON=1'b0;
    defparam \nx.mod_5_i873_3_lut_LC_1_32_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i873_3_lut_LC_1_32_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i873_3_lut_LC_1_32_2  (
            .in0(_gnd_net_),
            .in1(N__19005),
            .in2(N__22379),
            .in3(N__18987),
            .lcout(\nx.n1302 ),
            .ltout(\nx.n1302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_34_LC_1_32_3 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_34_LC_1_32_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_34_LC_1_32_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i1_2_lut_adj_34_LC_1_32_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18981),
            .in3(N__20537),
            .lcout(\nx.n10_adj_626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i879_3_lut_LC_1_32_4 .C_ON=1'b0;
    defparam \nx.mod_5_i879_3_lut_LC_1_32_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i879_3_lut_LC_1_32_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i879_3_lut_LC_1_32_4  (
            .in0(_gnd_net_),
            .in1(N__18978),
            .in2(N__22380),
            .in3(N__18972),
            .lcout(\nx.n1308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i809_3_lut_LC_1_32_5 .C_ON=1'b0;
    defparam \nx.mod_5_i809_3_lut_LC_1_32_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i809_3_lut_LC_1_32_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i809_3_lut_LC_1_32_5  (
            .in0(_gnd_net_),
            .in1(N__20301),
            .in2(N__25935),
            .in3(N__20427),
            .lcout(\nx.n1206 ),
            .ltout(\nx.n1206_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i876_3_lut_LC_1_32_6 .C_ON=1'b0;
    defparam \nx.mod_5_i876_3_lut_LC_1_32_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i876_3_lut_LC_1_32_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i876_3_lut_LC_1_32_6  (
            .in0(N__22377),
            .in1(_gnd_net_),
            .in2(N__18948),
            .in3(N__18945),
            .lcout(\nx.n1305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.start_103_LC_2_15_0 .C_ON=1'b0;
    defparam \nx.start_103_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \nx.start_103_LC_2_15_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \nx.start_103_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__19122),
            .in2(_gnd_net_),
            .in3(N__19527),
            .lcout(\nx.start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48390),
            .ce(N__18939),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i32_1_lut_LC_2_16_2 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i32_1_lut_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i32_1_lut_LC_2_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i32_1_lut_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20594),
            .lcout(\nx.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i24_1_lut_LC_2_17_1 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i24_1_lut_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i24_1_lut_LC_2_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i24_1_lut_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19049),
            .lcout(\nx.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_2 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_2 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_2  (
            .in0(N__19050),
            .in1(N__21611),
            .in2(_gnd_net_),
            .in3(N__28777),
            .lcout(neo_pixel_transmitter_t0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i24_LC_2_17_5 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i24_LC_2_17_5 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i24_LC_2_17_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i24_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__28774),
            .in2(N__19041),
            .in3(N__21555),
            .lcout(neo_pixel_transmitter_t0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48383),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i25_1_lut_LC_2_17_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i25_1_lut_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i25_1_lut_LC_2_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i25_1_lut_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19037),
            .lcout(\nx.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_done_104_LC_2_18_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_done_104_LC_2_18_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_done_104_LC_2_18_0 .LUT_INIT=16'b1100110000010001;
    LogicCell40 \nx.neo_pixel_transmitter_done_104_LC_2_18_0  (
            .in0(N__19142),
            .in1(N__19523),
            .in2(_gnd_net_),
            .in3(N__19271),
            .lcout(\nx.neo_pixel_transmitter_done ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48387),
            .ce(N__19026),
            .sr(_gnd_net_));
    defparam \nx.i2_2_lut_adj_149_LC_2_18_1 .C_ON=1'b0;
    defparam \nx.i2_2_lut_adj_149_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.i2_2_lut_adj_149_LC_2_18_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \nx.i2_2_lut_adj_149_LC_2_18_1  (
            .in0(N__21065),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21246),
            .lcout(),
            .ltout(\nx.n7_adj_713_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_4_lut_adj_150_LC_2_18_2 .C_ON=1'b0;
    defparam \nx.i4_4_lut_adj_150_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.i4_4_lut_adj_150_LC_2_18_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \nx.i4_4_lut_adj_150_LC_2_18_2  (
            .in0(N__20787),
            .in1(N__20733),
            .in2(N__19029),
            .in3(N__19089),
            .lcout(\nx.n13491 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_151_LC_2_18_3 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_151_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_151_LC_2_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \nx.i1_2_lut_adj_151_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__20786),
            .in2(_gnd_net_),
            .in3(N__20729),
            .lcout(),
            .ltout(\nx.n12933_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_152_LC_2_18_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_152_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_152_LC_2_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_152_LC_2_18_4  (
            .in0(N__21245),
            .in1(N__21228),
            .in2(N__19020),
            .in3(N__21166),
            .lcout(\nx.n12939 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i13_1_lut_LC_2_19_0 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i13_1_lut_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i13_1_lut_LC_2_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i13_1_lut_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19298),
            .lcout(\nx.n21_adj_620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2_2_lut_adj_154_LC_2_19_1 .C_ON=1'b0;
    defparam \nx.i2_2_lut_adj_154_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.i2_2_lut_adj_154_LC_2_19_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \nx.i2_2_lut_adj_154_LC_2_19_1  (
            .in0(N__20907),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20928),
            .lcout(\nx.n10918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i14_LC_2_19_2 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i14_LC_2_19_2 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i14_LC_2_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i14_LC_2_19_2  (
            .in0(N__19074),
            .in1(N__21440),
            .in2(_gnd_net_),
            .in3(N__28776),
            .lcout(neo_pixel_transmitter_t0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i7_1_lut_LC_2_19_3 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i7_1_lut_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i7_1_lut_LC_2_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i7_1_lut_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19082),
            .lcout(\nx.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_4_lut_adj_147_LC_2_19_4 .C_ON=1'b0;
    defparam \nx.i7_4_lut_adj_147_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.i7_4_lut_adj_147_LC_2_19_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \nx.i7_4_lut_adj_147_LC_2_19_4  (
            .in0(N__21130),
            .in1(N__19209),
            .in2(N__19516),
            .in3(N__21168),
            .lcout(),
            .ltout(\nx.n18_adj_711_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_148_LC_2_19_5 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_148_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_148_LC_2_19_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \nx.i9_4_lut_adj_148_LC_2_19_5  (
            .in0(N__19155),
            .in1(N__21227),
            .in2(N__19092),
            .in3(N__21710),
            .lcout(\nx.n20_adj_712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_19_6 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_19_6 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_19_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_19_6  (
            .in0(N__19083),
            .in1(N__28775),
            .in2(_gnd_net_),
            .in3(N__21282),
            .lcout(neo_pixel_transmitter_t0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48391),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i15_1_lut_LC_2_19_7 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i15_1_lut_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i15_1_lut_LC_2_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i15_1_lut_LC_2_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19073),
            .lcout(\nx.n19_adj_622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i6_1_lut_LC_2_20_0 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i6_1_lut_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i6_1_lut_LC_2_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i6_1_lut_LC_2_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19065),
            .lcout(\nx.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_221_LC_2_20_1.C_ON=1'b0;
    defparam i2_4_lut_adj_221_LC_2_20_1.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_221_LC_2_20_1.LUT_INIT=16'b0110111111110110;
    LogicCell40 i2_4_lut_adj_221_LC_2_20_1 (
            .in0(N__19329),
            .in1(N__39794),
            .in2(N__25005),
            .in3(N__28917),
            .lcout(n10_adj_776),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i4_1_lut_LC_2_20_2 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i4_1_lut_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i4_1_lut_LC_2_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i4_1_lut_LC_2_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19313),
            .lcout(\nx.n30_adj_598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i3_LC_2_20_3 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i3_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i3_LC_2_20_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i3_LC_2_20_3  (
            .in0(N__19314),
            .in1(N__28838),
            .in2(_gnd_net_),
            .in3(N__20876),
            .lcout(neo_pixel_transmitter_t0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48396),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_2_20_4.C_ON=1'b0;
    defparam i4_4_lut_LC_2_20_4.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_2_20_4.LUT_INIT=16'b0110111111110110;
    LogicCell40 i4_4_lut_LC_2_20_4 (
            .in0(N__38453),
            .in1(N__38427),
            .in2(N__43125),
            .in3(N__43167),
            .lcout(n12_adj_774),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i12_LC_2_20_5 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i12_LC_2_20_5 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i12_LC_2_20_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i12_LC_2_20_5  (
            .in0(N__21021),
            .in1(N__19299),
            .in2(_gnd_net_),
            .in3(N__28839),
            .lcout(neo_pixel_transmitter_t0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48396),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9545_2_lut_LC_2_20_6 .C_ON=1'b0;
    defparam \nx.i9545_2_lut_LC_2_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9545_2_lut_LC_2_20_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \nx.i9545_2_lut_LC_2_20_6  (
            .in0(N__19574),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19272),
            .lcout(),
            .ltout(\nx.n11487_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_146_LC_2_20_7 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_146_LC_2_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_146_LC_2_20_7 .LUT_INIT=16'b0111000001110101;
    LogicCell40 \nx.i1_4_lut_adj_146_LC_2_20_7  (
            .in0(N__20906),
            .in1(N__20924),
            .in2(N__19212),
            .in3(N__20849),
            .lcout(\nx.n103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_222_LC_2_21_0.C_ON=1'b0;
    defparam i1_4_lut_adj_222_LC_2_21_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_222_LC_2_21_0.LUT_INIT=16'b0110111111110110;
    LogicCell40 i1_4_lut_adj_222_LC_2_21_0 (
            .in0(N__40889),
            .in1(N__19188),
            .in2(N__37430),
            .in3(N__20199),
            .lcout(n9_adj_777),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i4_LC_2_21_1.C_ON=1'b0;
    defparam neopxl_color_prev_i4_LC_2_21_1.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i4_LC_2_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 neopxl_color_prev_i4_LC_2_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40890),
            .lcout(neopxl_color_prev_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48402),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4155_3_lut_LC_2_21_2 .C_ON=1'b0;
    defparam \nx.i4155_3_lut_LC_2_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i4155_3_lut_LC_2_21_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \nx.i4155_3_lut_LC_2_21_2  (
            .in0(N__19582),
            .in1(N__19504),
            .in2(_gnd_net_),
            .in3(N__19430),
            .lcout(\nx.n7392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i26_LC_2_21_3 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i26_LC_2_21_3 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i26_LC_2_21_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i26_LC_2_21_3  (
            .in0(N__28836),
            .in1(N__21491),
            .in2(_gnd_net_),
            .in3(N__19353),
            .lcout(neo_pixel_transmitter_t0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48402),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i16_LC_2_21_4 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i16_LC_2_21_4 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i16_LC_2_21_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i16_LC_2_21_4  (
            .in0(N__21354),
            .in1(N__19341),
            .in2(_gnd_net_),
            .in3(N__28837),
            .lcout(neo_pixel_transmitter_t0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48402),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9308_3_lut_LC_2_21_5 .C_ON=1'b0;
    defparam \nx.i9308_3_lut_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9308_3_lut_LC_2_21_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.i9308_3_lut_LC_2_21_5  (
            .in0(N__23991),
            .in1(N__40888),
            .in2(_gnd_net_),
            .in3(N__39793),
            .lcout(\nx.n13155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.bit_ctr_1__bdd_4_lut_LC_2_21_6 .C_ON=1'b0;
    defparam \nx.bit_ctr_1__bdd_4_lut_LC_2_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.bit_ctr_1__bdd_4_lut_LC_2_21_6 .LUT_INIT=16'b1100101011110000;
    LogicCell40 \nx.bit_ctr_1__bdd_4_lut_LC_2_21_6  (
            .in0(N__19659),
            .in1(N__22851),
            .in2(N__23940),
            .in3(N__19616),
            .lcout(),
            .ltout(\nx.n13456_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.n13456_bdd_4_lut_LC_2_21_7 .C_ON=1'b0;
    defparam \nx.n13456_bdd_4_lut_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.n13456_bdd_4_lut_LC_2_21_7 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \nx.n13456_bdd_4_lut_LC_2_21_7  (
            .in0(N__19617),
            .in1(N__19410),
            .in2(N__19404),
            .in3(N__19401),
            .lcout(\nx.n13459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_156_LC_2_22_0 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_156_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_156_LC_2_22_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \nx.i1_2_lut_adj_156_LC_2_22_0  (
            .in0(_gnd_net_),
            .in1(N__20905),
            .in2(_gnd_net_),
            .in3(N__20848),
            .lcout(\nx.n4_adj_642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i27_1_lut_LC_2_22_1 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i27_1_lut_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i27_1_lut_LC_2_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i27_1_lut_LC_2_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19352),
            .lcout(\nx.n7_adj_597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i17_1_lut_LC_2_22_2 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i17_1_lut_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i17_1_lut_LC_2_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i17_1_lut_LC_2_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19340),
            .lcout(\nx.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9470_3_lut_LC_2_22_3 .C_ON=1'b0;
    defparam \nx.i9470_3_lut_LC_2_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9470_3_lut_LC_2_22_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \nx.i9470_3_lut_LC_2_22_3  (
            .in0(N__20031),
            .in1(N__23889),
            .in2(_gnd_net_),
            .in3(N__19626),
            .lcout(\nx.color_bit_N_571_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9311_3_lut_LC_2_22_4 .C_ON=1'b0;
    defparam \nx.i9311_3_lut_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.i9311_3_lut_LC_2_22_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \nx.i9311_3_lut_LC_2_22_4  (
            .in0(N__28916),
            .in1(N__23989),
            .in2(_gnd_net_),
            .in3(N__38445),
            .lcout(\nx.n13158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i12_LC_2_22_5.C_ON=1'b0;
    defparam neopxl_color_i12_LC_2_22_5.SEQ_MODE=4'b1000;
    defparam neopxl_color_i12_LC_2_22_5.LUT_INIT=16'b1010101100101010;
    LogicCell40 neopxl_color_i12_LC_2_22_5 (
            .in0(N__38446),
            .in1(N__50079),
            .in2(N__49851),
            .in3(N__49589),
            .lcout(neopxl_color_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48407),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_130_LC_2_22_6 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_130_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_130_LC_2_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_130_LC_2_22_6  (
            .in0(N__19653),
            .in1(N__20232),
            .in2(N__19647),
            .in3(N__19638),
            .lcout(\nx.n10947 ),
            .ltout(\nx.n10947_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_58_LC_2_22_7 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_58_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_58_LC_2_22_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \nx.i1_2_lut_adj_58_LC_2_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19620),
            .in3(N__23888),
            .lcout(\nx.n10975 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2028_3_lut_LC_2_23_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2028_3_lut_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2028_3_lut_LC_2_23_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2028_3_lut_LC_2_23_0  (
            .in0(_gnd_net_),
            .in1(N__30411),
            .in2(N__25287),
            .in3(N__31852),
            .lcout(\nx.n3001 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2080_3_lut_LC_2_23_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2080_3_lut_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2080_3_lut_LC_2_23_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i2080_3_lut_LC_2_23_1  (
            .in0(_gnd_net_),
            .in1(N__27421),
            .in2(N__23460),
            .in3(N__22308),
            .lcout(\nx.n3085 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2035_3_lut_LC_2_23_2 .C_ON=1'b0;
    defparam \nx.mod_5_i2035_3_lut_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2035_3_lut_LC_2_23_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2035_3_lut_LC_2_23_2  (
            .in0(_gnd_net_),
            .in1(N__29776),
            .in2(N__25197),
            .in3(N__31851),
            .lcout(\nx.n3008 ),
            .ltout(\nx.n3008_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_96_LC_2_23_3 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_96_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_96_LC_2_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_96_LC_2_23_3  (
            .in0(N__23347),
            .in1(N__22030),
            .in2(N__19608),
            .in3(N__22084),
            .lcout(\nx.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2026_3_lut_LC_2_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2026_3_lut_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2026_3_lut_LC_2_23_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2026_3_lut_LC_2_23_4  (
            .in0(_gnd_net_),
            .in1(N__29715),
            .in2(N__25578),
            .in3(N__31853),
            .lcout(\nx.n2999 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2091_3_lut_LC_2_23_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2091_3_lut_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2091_3_lut_LC_2_23_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2091_3_lut_LC_2_23_5  (
            .in0(_gnd_net_),
            .in1(N__23319),
            .in2(N__21981),
            .in3(N__27422),
            .lcout(\nx.n3096 ),
            .ltout(\nx.n3096_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_adj_109_LC_2_23_6 .C_ON=1'b0;
    defparam \nx.i20_4_lut_adj_109_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_adj_109_LC_2_23_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i20_4_lut_adj_109_LC_2_23_6  (
            .in0(N__19966),
            .in1(N__19898),
            .in2(N__19776),
            .in3(N__20004),
            .lcout(\nx.n47_adj_694 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2096_3_lut_LC_2_24_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2096_3_lut_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2096_3_lut_LC_2_24_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2096_3_lut_LC_2_24_0  (
            .in0(_gnd_net_),
            .in1(N__22107),
            .in2(N__23534),
            .in3(N__27415),
            .lcout(\nx.n3101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i23_4_lut_adj_101_LC_2_24_1 .C_ON=1'b0;
    defparam \nx.i23_4_lut_adj_101_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.i23_4_lut_adj_101_LC_2_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i23_4_lut_adj_101_LC_2_24_1  (
            .in0(N__21869),
            .in1(N__23599),
            .in2(N__19764),
            .in3(N__23427),
            .lcout(),
            .ltout(\nx.n49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i25_4_lut_LC_2_24_2 .C_ON=1'b0;
    defparam \nx.i25_4_lut_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.i25_4_lut_LC_2_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i25_4_lut_LC_2_24_2  (
            .in0(N__23502),
            .in1(N__23547),
            .in2(N__19755),
            .in3(N__22986),
            .lcout(\nx.n3017 ),
            .ltout(\nx.n3017_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2082_3_lut_LC_2_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2082_3_lut_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2082_3_lut_LC_2_24_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2082_3_lut_LC_2_24_3  (
            .in0(_gnd_net_),
            .in1(N__23576),
            .in2(N__19752),
            .in3(N__22155),
            .lcout(\nx.n3087 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2081_3_lut_LC_2_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2081_3_lut_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2081_3_lut_LC_2_24_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i2081_3_lut_LC_2_24_4  (
            .in0(_gnd_net_),
            .in1(N__27420),
            .in2(N__23283),
            .in3(N__22140),
            .lcout(\nx.n3086 ),
            .ltout(\nx.n3086_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_103_LC_2_24_5 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_103_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_103_LC_2_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_103_LC_2_24_5  (
            .in0(N__19846),
            .in1(N__19717),
            .in2(N__19701),
            .in3(N__19690),
            .lcout(\nx.n42_adj_689 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2093_3_lut_LC_2_24_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2093_3_lut_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2093_3_lut_LC_2_24_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2093_3_lut_LC_2_24_6  (
            .in0(_gnd_net_),
            .in1(N__22031),
            .in2(N__22011),
            .in3(N__27419),
            .lcout(\nx.n3098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2098_3_lut_LC_2_24_7 .C_ON=1'b0;
    defparam \nx.mod_5_i2098_3_lut_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2098_3_lut_LC_2_24_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2098_3_lut_LC_2_24_7  (
            .in0(_gnd_net_),
            .in1(N__23600),
            .in2(N__27451),
            .in3(N__21813),
            .lcout(\nx.n3103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2092_3_lut_LC_2_25_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2092_3_lut_LC_2_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2092_3_lut_LC_2_25_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2092_3_lut_LC_2_25_0  (
            .in0(_gnd_net_),
            .in1(N__23159),
            .in2(N__21996),
            .in3(N__27399),
            .lcout(\nx.n3097 ),
            .ltout(\nx.n3097_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2159_3_lut_LC_2_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2159_3_lut_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2159_3_lut_LC_2_25_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2159_3_lut_LC_2_25_1  (
            .in0(_gnd_net_),
            .in1(N__19881),
            .in2(N__19872),
            .in3(N__24172),
            .lcout(),
            .ltout(\nx.n35_adj_699_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_113_LC_2_25_2 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_113_LC_2_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_113_LC_2_25_2 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \nx.i1_4_lut_adj_113_LC_2_25_2  (
            .in0(N__24173),
            .in1(N__19869),
            .in2(N__19860),
            .in3(N__19850),
            .lcout(\nx.n12337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2104_3_lut_LC_2_25_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2104_3_lut_LC_2_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2104_3_lut_LC_2_25_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i2104_3_lut_LC_2_25_3  (
            .in0(N__21927),
            .in1(_gnd_net_),
            .in2(N__27438),
            .in3(N__26175),
            .lcout(\nx.n3109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_120_LC_2_25_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_120_LC_2_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_120_LC_2_25_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \nx.i1_4_lut_adj_120_LC_2_25_4  (
            .in0(N__20027),
            .in1(N__23878),
            .in2(N__19929),
            .in3(N__19803),
            .lcout(\nx.n12353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2099_3_lut_LC_2_25_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2099_3_lut_LC_2_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2099_3_lut_LC_2_25_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2099_3_lut_LC_2_25_5  (
            .in0(_gnd_net_),
            .in1(N__23246),
            .in2(N__27437),
            .in3(N__21822),
            .lcout(\nx.n3104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2102_3_lut_LC_2_25_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2102_3_lut_LC_2_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2102_3_lut_LC_2_25_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2102_3_lut_LC_2_25_6  (
            .in0(_gnd_net_),
            .in1(N__21905),
            .in2(N__21888),
            .in3(N__27389),
            .lcout(\nx.n3107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2103_3_lut_LC_2_25_7 .C_ON=1'b0;
    defparam \nx.mod_5_i2103_3_lut_LC_2_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2103_3_lut_LC_2_25_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i2103_3_lut_LC_2_25_7  (
            .in0(N__23493),
            .in1(_gnd_net_),
            .in2(N__27439),
            .in3(N__21915),
            .lcout(\nx.n3108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_115_LC_2_26_0 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_115_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_115_LC_2_26_0 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \nx.i1_4_lut_adj_115_LC_2_26_0  (
            .in0(N__20118),
            .in1(N__20112),
            .in2(N__20106),
            .in3(N__24174),
            .lcout(),
            .ltout(\nx.n12327_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_117_LC_2_26_1 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_117_LC_2_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_117_LC_2_26_1 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \nx.i1_4_lut_adj_117_LC_2_26_1  (
            .in0(N__24176),
            .in1(N__20085),
            .in2(N__20079),
            .in3(N__20076),
            .lcout(\nx.n12339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2161_3_lut_LC_2_26_2 .C_ON=1'b0;
    defparam \nx.mod_5_i2161_3_lut_LC_2_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2161_3_lut_LC_2_26_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2161_3_lut_LC_2_26_2  (
            .in0(_gnd_net_),
            .in1(N__20222),
            .in2(N__20046),
            .in3(N__24177),
            .lcout(\nx.n31_adj_702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2172_3_lut_LC_2_26_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2172_3_lut_LC_2_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2172_3_lut_LC_2_26_3 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \nx.mod_5_i2172_3_lut_LC_2_26_3  (
            .in0(N__24370),
            .in1(N__20037),
            .in2(N__24208),
            .in3(_gnd_net_),
            .lcout(\nx.n3209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2166_3_lut_LC_2_26_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2166_3_lut_LC_2_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2166_3_lut_LC_2_26_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2166_3_lut_LC_2_26_4  (
            .in0(_gnd_net_),
            .in1(N__20016),
            .in2(N__23778),
            .in3(N__24175),
            .lcout(\nx.n21_adj_701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2170_3_lut_LC_2_26_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2170_3_lut_LC_2_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2170_3_lut_LC_2_26_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2170_3_lut_LC_2_26_5  (
            .in0(_gnd_net_),
            .in1(N__20010),
            .in2(N__24207),
            .in3(N__20002),
            .lcout(),
            .ltout(\nx.n13_adj_696_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_116_LC_2_26_6 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_116_LC_2_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_116_LC_2_26_6 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \nx.i1_4_lut_adj_116_LC_2_26_6  (
            .in0(N__19980),
            .in1(N__19974),
            .in2(N__19953),
            .in3(N__24181),
            .lcout(),
            .ltout(\nx.n12325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_118_LC_2_26_7 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_118_LC_2_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_118_LC_2_26_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_118_LC_2_26_7  (
            .in0(N__19950),
            .in1(N__19944),
            .in2(N__19938),
            .in3(N__19935),
            .lcout(\nx.n12347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2086_3_lut_LC_2_27_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2086_3_lut_LC_2_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2086_3_lut_LC_2_27_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2086_3_lut_LC_2_27_0  (
            .in0(_gnd_net_),
            .in1(N__22173),
            .in2(N__23847),
            .in3(N__27440),
            .lcout(\nx.n3091 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2146_3_lut_LC_2_27_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2146_3_lut_LC_2_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2146_3_lut_LC_2_27_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i2146_3_lut_LC_2_27_3  (
            .in0(N__20138),
            .in1(N__20241),
            .in2(_gnd_net_),
            .in3(N__24234),
            .lcout(\nx.n61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2094_3_lut_LC_2_27_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2094_3_lut_LC_2_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2094_3_lut_LC_2_27_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2094_3_lut_LC_2_27_6  (
            .in0(_gnd_net_),
            .in1(N__23390),
            .in2(N__22050),
            .in3(N__27441),
            .lcout(\nx.n3099 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i7_LC_2_27_7.C_ON=1'b0;
    defparam neopxl_color_prev_i7_LC_2_27_7.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i7_LC_2_27_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 neopxl_color_prev_i7_LC_2_27_7 (
            .in0(_gnd_net_),
            .in1(N__37423),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(neopxl_color_prev_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48419),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i26_4_lut_adj_141_LC_2_28_0 .C_ON=1'b0;
    defparam \nx.i26_4_lut_adj_141_LC_2_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.i26_4_lut_adj_141_LC_2_28_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i26_4_lut_adj_141_LC_2_28_0  (
            .in0(N__25953),
            .in1(N__24501),
            .in2(N__26406),
            .in3(N__22257),
            .lcout(\nx.n54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i21_4_lut_adj_142_LC_2_28_2 .C_ON=1'b0;
    defparam \nx.i21_4_lut_adj_142_LC_2_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.i21_4_lut_adj_142_LC_2_28_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i21_4_lut_adj_142_LC_2_28_2  (
            .in0(N__34977),
            .in1(N__28069),
            .in2(N__24462),
            .in3(N__28533),
            .lcout(\nx.n49_adj_710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_140_LC_2_28_3 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_140_LC_2_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_140_LC_2_28_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \nx.i15_4_lut_adj_140_LC_2_28_3  (
            .in0(N__23887),
            .in1(N__24374),
            .in2(N__39846),
            .in3(N__32682),
            .lcout(),
            .ltout(\nx.n43_adj_709_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i27_4_lut_LC_2_28_4 .C_ON=1'b0;
    defparam \nx.i27_4_lut_LC_2_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.i27_4_lut_LC_2_28_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i27_4_lut_LC_2_28_4  (
            .in0(N__20187),
            .in1(N__26091),
            .in2(N__20181),
            .in3(N__20178),
            .lcout(state_3_N_377_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2079_3_lut_LC_2_28_7 .C_ON=1'b0;
    defparam \nx.mod_5_i2079_3_lut_LC_2_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2079_3_lut_LC_2_28_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2079_3_lut_LC_2_28_7  (
            .in0(_gnd_net_),
            .in1(N__22293),
            .in2(N__23127),
            .in3(N__27459),
            .lcout(\nx.n3084 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_2_lut_LC_2_29_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_2_lut_LC_2_29_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_2_lut_LC_2_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_2_lut_LC_2_29_0  (
            .in0(_gnd_net_),
            .in1(N__24456),
            .in2(_gnd_net_),
            .in3(N__20340),
            .lcout(\nx.n1177 ),
            .ltout(),
            .carryin(bfn_2_29_0_),
            .carryout(\nx.n10461 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_3_lut_LC_2_29_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_3_lut_LC_2_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_3_lut_LC_2_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_3_lut_LC_2_29_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20337),
            .in3(N__20307),
            .lcout(\nx.n1176 ),
            .ltout(),
            .carryin(\nx.n10461 ),
            .carryout(\nx.n10462 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_4_lut_LC_2_29_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_4_lut_LC_2_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_4_lut_LC_2_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_4_lut_LC_2_29_2  (
            .in0(_gnd_net_),
            .in1(N__45280),
            .in2(N__26352),
            .in3(N__20304),
            .lcout(\nx.n1175 ),
            .ltout(),
            .carryin(\nx.n10462 ),
            .carryout(\nx.n10463 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_5_lut_LC_2_29_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_5_lut_LC_2_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_5_lut_LC_2_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_5_lut_LC_2_29_3  (
            .in0(_gnd_net_),
            .in1(N__45284),
            .in2(N__25930),
            .in3(N__20292),
            .lcout(\nx.n1174 ),
            .ltout(),
            .carryin(\nx.n10463 ),
            .carryout(\nx.n10464 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_6_lut_LC_2_29_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_6_lut_LC_2_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_6_lut_LC_2_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_6_lut_LC_2_29_4  (
            .in0(_gnd_net_),
            .in1(N__45281),
            .in2(N__26292),
            .in3(N__20289),
            .lcout(\nx.n1173 ),
            .ltout(),
            .carryin(\nx.n10464 ),
            .carryout(\nx.n10465 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_7_lut_LC_2_29_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_7_lut_LC_2_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_7_lut_LC_2_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_7_lut_LC_2_29_5  (
            .in0(_gnd_net_),
            .in1(N__45285),
            .in2(N__25896),
            .in3(N__20286),
            .lcout(\nx.n1172 ),
            .ltout(),
            .carryin(\nx.n10465 ),
            .carryout(\nx.n10466 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_8_lut_LC_2_29_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_8_lut_LC_2_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_8_lut_LC_2_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_8_lut_LC_2_29_6  (
            .in0(_gnd_net_),
            .in1(N__45282),
            .in2(N__26016),
            .in3(N__20274),
            .lcout(\nx.n1171 ),
            .ltout(),
            .carryin(\nx.n10466 ),
            .carryout(\nx.n10467 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_9_lut_LC_2_29_7 .C_ON=1'b0;
    defparam \nx.mod_5_add_803_9_lut_LC_2_29_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_9_lut_LC_2_29_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_803_9_lut_LC_2_29_7  (
            .in0(N__45283),
            .in1(N__20419),
            .in2(N__25977),
            .in3(N__20271),
            .lcout(\nx.n1202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i808_3_lut_LC_2_30_0 .C_ON=1'b0;
    defparam \nx.mod_5_i808_3_lut_LC_2_30_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i808_3_lut_LC_2_30_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i808_3_lut_LC_2_30_0  (
            .in0(_gnd_net_),
            .in1(N__26291),
            .in2(N__20250),
            .in3(N__20412),
            .lcout(\nx.n1205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i807_3_lut_LC_2_30_1 .C_ON=1'b0;
    defparam \nx.mod_5_i807_3_lut_LC_2_30_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i807_3_lut_LC_2_30_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i807_3_lut_LC_2_30_1  (
            .in0(_gnd_net_),
            .in1(N__25895),
            .in2(N__20425),
            .in3(N__20523),
            .lcout(\nx.n1204 ),
            .ltout(\nx.n1204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i874_3_lut_LC_2_30_2 .C_ON=1'b0;
    defparam \nx.mod_5_i874_3_lut_LC_2_30_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i874_3_lut_LC_2_30_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i874_3_lut_LC_2_30_2  (
            .in0(_gnd_net_),
            .in1(N__20502),
            .in2(N__20496),
            .in3(N__22367),
            .lcout(\nx.n1303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_4_lut_adj_32_LC_2_30_3 .C_ON=1'b0;
    defparam \nx.i7_4_lut_adj_32_LC_2_30_3 .SEQ_MODE=4'b0000;
    defparam \nx.i7_4_lut_adj_32_LC_2_30_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i7_4_lut_adj_32_LC_2_30_3  (
            .in0(N__20381),
            .in1(N__20493),
            .in2(N__20487),
            .in3(N__20478),
            .lcout(\nx.n1235 ),
            .ltout(\nx.n1235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i878_3_lut_LC_2_30_4 .C_ON=1'b0;
    defparam \nx.mod_5_i878_3_lut_LC_2_30_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i878_3_lut_LC_2_30_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i878_3_lut_LC_2_30_4  (
            .in0(_gnd_net_),
            .in1(N__20457),
            .in2(N__20451),
            .in3(N__20447),
            .lcout(\nx.n1307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i810_3_lut_LC_2_30_5 .C_ON=1'b0;
    defparam \nx.mod_5_i810_3_lut_LC_2_30_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i810_3_lut_LC_2_30_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i810_3_lut_LC_2_30_5  (
            .in0(_gnd_net_),
            .in1(N__20433),
            .in2(N__20426),
            .in3(N__26347),
            .lcout(\nx.n1207 ),
            .ltout(\nx.n1207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i877_3_lut_LC_2_30_6 .C_ON=1'b0;
    defparam \nx.mod_5_i877_3_lut_LC_2_30_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i877_3_lut_LC_2_30_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i877_3_lut_LC_2_30_6  (
            .in0(N__20370),
            .in1(_gnd_net_),
            .in2(N__20364),
            .in3(N__22366),
            .lcout(\nx.n1306 ),
            .ltout(\nx.n1306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_4_lut_adj_35_LC_2_30_7 .C_ON=1'b0;
    defparam \nx.i7_4_lut_adj_35_LC_2_30_7 .SEQ_MODE=4'b0000;
    defparam \nx.i7_4_lut_adj_35_LC_2_30_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i7_4_lut_adj_35_LC_2_30_7  (
            .in0(N__22240),
            .in1(N__24733),
            .in2(N__20361),
            .in3(N__20358),
            .lcout(\nx.n16_adj_627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_2_lut_LC_2_31_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_2_lut_LC_2_31_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_2_lut_LC_2_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_2_lut_LC_2_31_0  (
            .in0(_gnd_net_),
            .in1(N__32717),
            .in2(_gnd_net_),
            .in3(N__20349),
            .lcout(\nx.n1377 ),
            .ltout(),
            .carryin(bfn_2_31_0_),
            .carryout(\nx.n10573 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_3_lut_LC_2_31_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_3_lut_LC_2_31_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_3_lut_LC_2_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_3_lut_LC_2_31_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22203),
            .in3(N__20565),
            .lcout(\nx.n1376 ),
            .ltout(),
            .carryin(\nx.n10573 ),
            .carryout(\nx.n10574 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_4_lut_LC_2_31_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_4_lut_LC_2_31_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_4_lut_LC_2_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_4_lut_LC_2_31_2  (
            .in0(_gnd_net_),
            .in1(N__45298),
            .in2(N__24734),
            .in3(N__20562),
            .lcout(\nx.n1375 ),
            .ltout(),
            .carryin(\nx.n10574 ),
            .carryout(\nx.n10575 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_5_lut_LC_2_31_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_5_lut_LC_2_31_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_5_lut_LC_2_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_5_lut_LC_2_31_3  (
            .in0(_gnd_net_),
            .in1(N__22241),
            .in2(N__45628),
            .in3(N__20559),
            .lcout(\nx.n1374 ),
            .ltout(),
            .carryin(\nx.n10575 ),
            .carryout(\nx.n10576 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_6_lut_LC_2_31_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_6_lut_LC_2_31_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_6_lut_LC_2_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_6_lut_LC_2_31_4  (
            .in0(_gnd_net_),
            .in1(N__45302),
            .in2(N__24683),
            .in3(N__20556),
            .lcout(\nx.n1373 ),
            .ltout(),
            .carryin(\nx.n10576 ),
            .carryout(\nx.n10577 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_7_lut_LC_2_31_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_7_lut_LC_2_31_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_7_lut_LC_2_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_7_lut_LC_2_31_5  (
            .in0(_gnd_net_),
            .in1(N__45303),
            .in2(N__24631),
            .in3(N__20553),
            .lcout(\nx.n1372 ),
            .ltout(),
            .carryin(\nx.n10577 ),
            .carryout(\nx.n10578 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_8_lut_LC_2_31_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_8_lut_LC_2_31_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_8_lut_LC_2_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_8_lut_LC_2_31_6  (
            .in0(_gnd_net_),
            .in1(N__24652),
            .in2(N__45629),
            .in3(N__20550),
            .lcout(\nx.n1371 ),
            .ltout(),
            .carryin(\nx.n10578 ),
            .carryout(\nx.n10579 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_9_lut_LC_2_31_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_9_lut_LC_2_31_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_9_lut_LC_2_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_9_lut_LC_2_31_7  (
            .in0(_gnd_net_),
            .in1(N__45307),
            .in2(N__22517),
            .in3(N__20547),
            .lcout(\nx.n1370 ),
            .ltout(),
            .carryin(\nx.n10579 ),
            .carryout(\nx.n10580 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_10_lut_LC_2_32_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_10_lut_LC_2_32_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_10_lut_LC_2_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_10_lut_LC_2_32_0  (
            .in0(_gnd_net_),
            .in1(N__44833),
            .in2(N__20625),
            .in3(N__20544),
            .lcout(\nx.n1369 ),
            .ltout(),
            .carryin(bfn_2_32_0_),
            .carryout(\nx.n10581 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_11_lut_LC_2_32_1 .C_ON=1'b0;
    defparam \nx.mod_5_add_937_11_lut_LC_2_32_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_11_lut_LC_2_32_1 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_937_11_lut_LC_2_32_1  (
            .in0(N__44834),
            .in1(N__24589),
            .in2(N__20541),
            .in3(N__20526),
            .lcout(\nx.n1400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i940_3_lut_LC_2_32_5 .C_ON=1'b0;
    defparam \nx.mod_5_i940_3_lut_LC_2_32_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i940_3_lut_LC_2_32_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i940_3_lut_LC_2_32_5  (
            .in0(_gnd_net_),
            .in1(N__20624),
            .in2(N__20613),
            .in3(N__24588),
            .lcout(\nx.n1401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i4_LC_3_15_1 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i4_LC_3_15_1 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i4_LC_3_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i4_LC_3_15_1  (
            .in0(N__20583),
            .in1(N__20817),
            .in2(_gnd_net_),
            .in3(N__28858),
            .lcout(neo_pixel_transmitter_t0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48397),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i1_LC_3_15_2 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i1_LC_3_15_2 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i1_LC_3_15_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i1_LC_3_15_2  (
            .in0(N__28857),
            .in1(N__20951),
            .in2(_gnd_net_),
            .in3(N__20604),
            .lcout(neo_pixel_transmitter_t0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48397),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i2_1_lut_LC_3_15_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i2_1_lut_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i2_1_lut_LC_3_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i2_1_lut_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20603),
            .lcout(\nx.n32_adj_651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i31_LC_3_16_1 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i31_LC_3_16_1 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i31_LC_3_16_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i31_LC_3_16_1  (
            .in0(N__28841),
            .in1(N__21765),
            .in2(_gnd_net_),
            .in3(N__20595),
            .lcout(neo_pixel_transmitter_t0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48392),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i10_LC_3_16_3 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i10_LC_3_16_3 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i10_LC_3_16_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i10_LC_3_16_3  (
            .in0(N__28840),
            .in1(N__21096),
            .in2(_gnd_net_),
            .in3(N__22610),
            .lcout(neo_pixel_transmitter_t0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48392),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i5_1_lut_LC_3_16_7 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i5_1_lut_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i5_1_lut_LC_3_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i5_1_lut_LC_3_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20582),
            .lcout(\nx.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i0_LC_3_17_0 .C_ON=1'b1;
    defparam \nx.timer_1102__i0_LC_3_17_0 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i0_LC_3_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i0_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__28666),
            .in2(_gnd_net_),
            .in3(N__20571),
            .lcout(timer_0),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\nx.n10479 ),
            .clk(N__48385),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i1_LC_3_17_1 .C_ON=1'b1;
    defparam \nx.timer_1102__i1_LC_3_17_1 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i1_LC_3_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i1_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__20947),
            .in2(_gnd_net_),
            .in3(N__20568),
            .lcout(timer_1),
            .ltout(),
            .carryin(\nx.n10479 ),
            .carryout(\nx.n10480 ),
            .clk(N__48385),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i2_LC_3_17_2 .C_ON=1'b1;
    defparam \nx.timer_1102__i2_LC_3_17_2 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i2_LC_3_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i2_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__22693),
            .in2(_gnd_net_),
            .in3(N__20655),
            .lcout(timer_2),
            .ltout(),
            .carryin(\nx.n10480 ),
            .carryout(\nx.n10481 ),
            .clk(N__48385),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i3_LC_3_17_3 .C_ON=1'b1;
    defparam \nx.timer_1102__i3_LC_3_17_3 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i3_LC_3_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i3_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__20869),
            .in2(_gnd_net_),
            .in3(N__20652),
            .lcout(timer_3),
            .ltout(),
            .carryin(\nx.n10481 ),
            .carryout(\nx.n10482 ),
            .clk(N__48385),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i4_LC_3_17_4 .C_ON=1'b1;
    defparam \nx.timer_1102__i4_LC_3_17_4 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i4_LC_3_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i4_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__20803),
            .in2(_gnd_net_),
            .in3(N__20649),
            .lcout(timer_4),
            .ltout(),
            .carryin(\nx.n10482 ),
            .carryout(\nx.n10483 ),
            .clk(N__48385),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i5_LC_3_17_5 .C_ON=1'b1;
    defparam \nx.timer_1102__i5_LC_3_17_5 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i5_LC_3_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i5_LC_3_17_5  (
            .in0(_gnd_net_),
            .in1(N__20761),
            .in2(_gnd_net_),
            .in3(N__20646),
            .lcout(timer_5),
            .ltout(),
            .carryin(\nx.n10483 ),
            .carryout(\nx.n10484 ),
            .clk(N__48385),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i6_LC_3_17_6 .C_ON=1'b1;
    defparam \nx.timer_1102__i6_LC_3_17_6 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i6_LC_3_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i6_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__21277),
            .in2(_gnd_net_),
            .in3(N__20643),
            .lcout(timer_6),
            .ltout(),
            .carryin(\nx.n10484 ),
            .carryout(\nx.n10485 ),
            .clk(N__48385),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i7_LC_3_17_7 .C_ON=1'b1;
    defparam \nx.timer_1102__i7_LC_3_17_7 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i7_LC_3_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i7_LC_3_17_7  (
            .in0(_gnd_net_),
            .in1(N__22870),
            .in2(_gnd_net_),
            .in3(N__20640),
            .lcout(timer_7),
            .ltout(),
            .carryin(\nx.n10485 ),
            .carryout(\nx.n10486 ),
            .clk(N__48385),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i8_LC_3_18_0 .C_ON=1'b1;
    defparam \nx.timer_1102__i8_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i8_LC_3_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i8_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__21187),
            .in2(_gnd_net_),
            .in3(N__20637),
            .lcout(timer_8),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\nx.n10487 ),
            .clk(N__48393),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i9_LC_3_18_1 .C_ON=1'b1;
    defparam \nx.timer_1102__i9_LC_3_18_1 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i9_LC_3_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i9_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__22630),
            .in2(_gnd_net_),
            .in3(N__20634),
            .lcout(timer_9),
            .ltout(),
            .carryin(\nx.n10487 ),
            .carryout(\nx.n10488 ),
            .clk(N__48393),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i10_LC_3_18_2 .C_ON=1'b1;
    defparam \nx.timer_1102__i10_LC_3_18_2 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i10_LC_3_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i10_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(N__21082),
            .in2(_gnd_net_),
            .in3(N__20631),
            .lcout(timer_10),
            .ltout(),
            .carryin(\nx.n10488 ),
            .carryout(\nx.n10489 ),
            .clk(N__48393),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i11_LC_3_18_3 .C_ON=1'b1;
    defparam \nx.timer_1102__i11_LC_3_18_3 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i11_LC_3_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i11_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__22552),
            .in2(_gnd_net_),
            .in3(N__20628),
            .lcout(timer_11),
            .ltout(),
            .carryin(\nx.n10489 ),
            .carryout(\nx.n10490 ),
            .clk(N__48393),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i12_LC_3_18_4 .C_ON=1'b1;
    defparam \nx.timer_1102__i12_LC_3_18_4 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i12_LC_3_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i12_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(N__21016),
            .in2(_gnd_net_),
            .in3(N__20682),
            .lcout(timer_12),
            .ltout(),
            .carryin(\nx.n10490 ),
            .carryout(\nx.n10491 ),
            .clk(N__48393),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i13_LC_3_18_5 .C_ON=1'b1;
    defparam \nx.timer_1102__i13_LC_3_18_5 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i13_LC_3_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i13_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(N__22942),
            .in2(_gnd_net_),
            .in3(N__20679),
            .lcout(timer_13),
            .ltout(),
            .carryin(\nx.n10491 ),
            .carryout(\nx.n10492 ),
            .clk(N__48393),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i14_LC_3_18_6 .C_ON=1'b1;
    defparam \nx.timer_1102__i14_LC_3_18_6 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i14_LC_3_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i14_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__21439),
            .in2(_gnd_net_),
            .in3(N__20676),
            .lcout(timer_14),
            .ltout(),
            .carryin(\nx.n10492 ),
            .carryout(\nx.n10493 ),
            .clk(N__48393),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i15_LC_3_18_7 .C_ON=1'b1;
    defparam \nx.timer_1102__i15_LC_3_18_7 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i15_LC_3_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i15_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__21388),
            .in2(_gnd_net_),
            .in3(N__20673),
            .lcout(timer_15),
            .ltout(),
            .carryin(\nx.n10493 ),
            .carryout(\nx.n10494 ),
            .clk(N__48393),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i16_LC_3_19_0 .C_ON=1'b1;
    defparam \nx.timer_1102__i16_LC_3_19_0 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i16_LC_3_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i16_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__21337),
            .in2(_gnd_net_),
            .in3(N__20670),
            .lcout(timer_16),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\nx.n10495 ),
            .clk(N__48398),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i17_LC_3_19_1 .C_ON=1'b1;
    defparam \nx.timer_1102__i17_LC_3_19_1 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i17_LC_3_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i17_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__22729),
            .in2(_gnd_net_),
            .in3(N__20667),
            .lcout(timer_17),
            .ltout(),
            .carryin(\nx.n10495 ),
            .carryout(\nx.n10496 ),
            .clk(N__48398),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i18_LC_3_19_2 .C_ON=1'b1;
    defparam \nx.timer_1102__i18_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i18_LC_3_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i18_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__22783),
            .in2(_gnd_net_),
            .in3(N__20664),
            .lcout(timer_18),
            .ltout(),
            .carryin(\nx.n10496 ),
            .carryout(\nx.n10497 ),
            .clk(N__48398),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i19_LC_3_19_3 .C_ON=1'b1;
    defparam \nx.timer_1102__i19_LC_3_19_3 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i19_LC_3_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i19_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__25120),
            .in2(_gnd_net_),
            .in3(N__20661),
            .lcout(timer_19),
            .ltout(),
            .carryin(\nx.n10497 ),
            .carryout(\nx.n10498 ),
            .clk(N__48398),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i20_LC_3_19_4 .C_ON=1'b1;
    defparam \nx.timer_1102__i20_LC_3_19_4 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i20_LC_3_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i20_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__25168),
            .in2(_gnd_net_),
            .in3(N__20658),
            .lcout(timer_20),
            .ltout(),
            .carryin(\nx.n10498 ),
            .carryout(\nx.n10499 ),
            .clk(N__48398),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i21_LC_3_19_5 .C_ON=1'b1;
    defparam \nx.timer_1102__i21_LC_3_19_5 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i21_LC_3_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i21_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__22969),
            .in2(_gnd_net_),
            .in3(N__20709),
            .lcout(timer_21),
            .ltout(),
            .carryin(\nx.n10499 ),
            .carryout(\nx.n10500 ),
            .clk(N__48398),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i22_LC_3_19_6 .C_ON=1'b1;
    defparam \nx.timer_1102__i22_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i22_LC_3_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i22_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__24868),
            .in2(_gnd_net_),
            .in3(N__20706),
            .lcout(timer_22),
            .ltout(),
            .carryin(\nx.n10500 ),
            .carryout(\nx.n10501 ),
            .clk(N__48398),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i23_LC_3_19_7 .C_ON=1'b1;
    defparam \nx.timer_1102__i23_LC_3_19_7 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i23_LC_3_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i23_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__21598),
            .in2(_gnd_net_),
            .in3(N__20703),
            .lcout(timer_23),
            .ltout(),
            .carryin(\nx.n10501 ),
            .carryout(\nx.n10502 ),
            .clk(N__48398),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i24_LC_3_20_0 .C_ON=1'b1;
    defparam \nx.timer_1102__i24_LC_3_20_0 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i24_LC_3_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i24_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__21547),
            .in2(_gnd_net_),
            .in3(N__20700),
            .lcout(timer_24),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\nx.n10503 ),
            .clk(N__48403),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i25_LC_3_20_1 .C_ON=1'b1;
    defparam \nx.timer_1102__i25_LC_3_20_1 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i25_LC_3_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i25_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__22807),
            .in2(_gnd_net_),
            .in3(N__20697),
            .lcout(timer_25),
            .ltout(),
            .carryin(\nx.n10503 ),
            .carryout(\nx.n10504 ),
            .clk(N__48403),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i26_LC_3_20_2 .C_ON=1'b1;
    defparam \nx.timer_1102__i26_LC_3_20_2 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i26_LC_3_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i26_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__21481),
            .in2(_gnd_net_),
            .in3(N__20694),
            .lcout(timer_26),
            .ltout(),
            .carryin(\nx.n10504 ),
            .carryout(\nx.n10505 ),
            .clk(N__48403),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i27_LC_3_20_3 .C_ON=1'b1;
    defparam \nx.timer_1102__i27_LC_3_20_3 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i27_LC_3_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i27_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__21670),
            .in2(_gnd_net_),
            .in3(N__20691),
            .lcout(timer_27),
            .ltout(),
            .carryin(\nx.n10505 ),
            .carryout(\nx.n10506 ),
            .clk(N__48403),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i28_LC_3_20_4 .C_ON=1'b1;
    defparam \nx.timer_1102__i28_LC_3_20_4 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i28_LC_3_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i28_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__23029),
            .in2(_gnd_net_),
            .in3(N__20688),
            .lcout(timer_28),
            .ltout(),
            .carryin(\nx.n10506 ),
            .carryout(\nx.n10507 ),
            .clk(N__48403),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i29_LC_3_20_5 .C_ON=1'b1;
    defparam \nx.timer_1102__i29_LC_3_20_5 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i29_LC_3_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i29_LC_3_20_5  (
            .in0(_gnd_net_),
            .in1(N__22654),
            .in2(_gnd_net_),
            .in3(N__20685),
            .lcout(timer_29),
            .ltout(),
            .carryin(\nx.n10507 ),
            .carryout(\nx.n10508 ),
            .clk(N__48403),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i30_LC_3_20_6 .C_ON=1'b1;
    defparam \nx.timer_1102__i30_LC_3_20_6 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i30_LC_3_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i30_LC_3_20_6  (
            .in0(_gnd_net_),
            .in1(N__22444),
            .in2(_gnd_net_),
            .in3(N__20967),
            .lcout(timer_30),
            .ltout(),
            .carryin(\nx.n10508 ),
            .carryout(\nx.n10509 ),
            .clk(N__48403),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_1102__i31_LC_3_20_7 .C_ON=1'b0;
    defparam \nx.timer_1102__i31_LC_3_20_7 .SEQ_MODE=4'b1000;
    defparam \nx.timer_1102__i31_LC_3_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_1102__i31_LC_3_20_7  (
            .in0(_gnd_net_),
            .in1(N__21757),
            .in2(_gnd_net_),
            .in3(N__20964),
            .lcout(timer_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48403),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_2_LC_3_21_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_2_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_2_LC_3_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_2_LC_3_21_0  (
            .in0(_gnd_net_),
            .in1(N__28635),
            .in2(N__28677),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_21_0_),
            .carryout(\nx.n10422 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_3_lut_LC_3_21_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_3_lut_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_3_lut_LC_3_21_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \nx.sub_14_add_2_3_lut_LC_3_21_1  (
            .in0(N__20850),
            .in1(N__20961),
            .in2(N__20952),
            .in3(N__20910),
            .lcout(\nx.n11533 ),
            .ltout(),
            .carryin(\nx.n10422 ),
            .carryout(\nx.n10423 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_4_lut_LC_3_21_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_4_lut_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_4_lut_LC_3_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_4_lut_LC_3_21_2  (
            .in0(_gnd_net_),
            .in1(N__22764),
            .in2(N__22698),
            .in3(N__20886),
            .lcout(\nx.one_wire_N_528_2 ),
            .ltout(),
            .carryin(\nx.n10423 ),
            .carryout(\nx.n10424 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_5_lut_LC_3_21_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_5_lut_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_5_lut_LC_3_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_5_lut_LC_3_21_3  (
            .in0(_gnd_net_),
            .in1(N__20883),
            .in2(N__20877),
            .in3(N__20829),
            .lcout(\nx.one_wire_N_528_3 ),
            .ltout(),
            .carryin(\nx.n10424 ),
            .carryout(\nx.n10425 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_6_lut_LC_3_21_4 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_6_lut_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_6_lut_LC_3_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_6_lut_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(N__20826),
            .in2(N__20816),
            .in3(N__20775),
            .lcout(\nx.one_wire_N_528_4 ),
            .ltout(),
            .carryin(\nx.n10425 ),
            .carryout(\nx.n10426 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_7_lut_LC_3_21_5 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_7_lut_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_7_lut_LC_3_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_7_lut_LC_3_21_5  (
            .in0(_gnd_net_),
            .in1(N__20771),
            .in2(N__20742),
            .in3(N__20712),
            .lcout(\nx.one_wire_N_528_5 ),
            .ltout(),
            .carryin(\nx.n10426 ),
            .carryout(\nx.n10427 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_8_lut_LC_3_21_6 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_8_lut_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_8_lut_LC_3_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_8_lut_LC_3_21_6  (
            .in0(_gnd_net_),
            .in1(N__21281),
            .in2(N__21258),
            .in3(N__21231),
            .lcout(\nx.one_wire_N_528_6 ),
            .ltout(),
            .carryin(\nx.n10427 ),
            .carryout(\nx.n10428 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_9_lut_LC_3_21_7 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_9_lut_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_9_lut_LC_3_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_9_lut_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(N__23199),
            .in2(N__22881),
            .in3(N__21210),
            .lcout(\nx.one_wire_N_528_7 ),
            .ltout(),
            .carryin(\nx.n10428 ),
            .carryout(\nx.n10429 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_10_lut_LC_3_22_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_10_lut_LC_3_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_10_lut_LC_3_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_10_lut_LC_3_22_0  (
            .in0(_gnd_net_),
            .in1(N__21207),
            .in2(N__21197),
            .in3(N__21138),
            .lcout(\nx.one_wire_N_528_8 ),
            .ltout(),
            .carryin(bfn_3_22_0_),
            .carryout(\nx.n10430 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_11_lut_LC_3_22_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_11_lut_LC_3_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_11_lut_LC_3_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_11_lut_LC_3_22_1  (
            .in0(_gnd_net_),
            .in1(N__25074),
            .in2(N__22635),
            .in3(N__21099),
            .lcout(\nx.one_wire_N_528_9 ),
            .ltout(),
            .carryin(\nx.n10430 ),
            .carryout(\nx.n10431 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_12_lut_LC_3_22_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_12_lut_LC_3_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_12_lut_LC_3_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_12_lut_LC_3_22_2  (
            .in0(_gnd_net_),
            .in1(N__22596),
            .in2(N__21095),
            .in3(N__21033),
            .lcout(\nx.one_wire_N_528_10 ),
            .ltout(),
            .carryin(\nx.n10431 ),
            .carryout(\nx.n10432 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_13_lut_LC_3_22_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_13_lut_LC_3_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_13_lut_LC_3_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_13_lut_LC_3_22_3  (
            .in0(_gnd_net_),
            .in1(N__22911),
            .in2(N__22557),
            .in3(N__21030),
            .lcout(\nx.one_wire_N_528_11 ),
            .ltout(),
            .carryin(\nx.n10432 ),
            .carryout(\nx.n10433 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_14_lut_LC_3_22_4 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_14_lut_LC_3_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_14_lut_LC_3_22_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_14_lut_LC_3_22_4  (
            .in0(N__21027),
            .in1(N__21020),
            .in2(N__20997),
            .in3(N__20979),
            .lcout(\nx.n12945 ),
            .ltout(),
            .carryin(\nx.n10433 ),
            .carryout(\nx.n10434 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_15_lut_LC_3_22_5 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_15_lut_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_15_lut_LC_3_22_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_15_lut_LC_3_22_5  (
            .in0(N__20976),
            .in1(N__22890),
            .in2(N__22950),
            .in3(N__20970),
            .lcout(\nx.n12947 ),
            .ltout(),
            .carryin(\nx.n10434 ),
            .carryout(\nx.n10435 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_16_lut_LC_3_22_6 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_16_lut_LC_3_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_16_lut_LC_3_22_6 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_16_lut_LC_3_22_6  (
            .in0(N__21462),
            .in1(N__21456),
            .in2(N__21447),
            .in3(N__21420),
            .lcout(\nx.n12949 ),
            .ltout(),
            .carryin(\nx.n10435 ),
            .carryout(\nx.n10436 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_16_THRU_CRY_0_LC_3_22_7 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_16_THRU_CRY_0_LC_3_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_16_THRU_CRY_0_LC_3_22_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_16_THRU_CRY_0_LC_3_22_7  (
            .in0(_gnd_net_),
            .in1(N__45757),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10436 ),
            .carryout(\nx.n10436_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_17_lut_LC_3_23_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_17_lut_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_17_lut_LC_3_23_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_17_lut_LC_3_23_0  (
            .in0(N__21417),
            .in1(N__21411),
            .in2(N__21398),
            .in3(N__21369),
            .lcout(\nx.n12951 ),
            .ltout(),
            .carryin(bfn_3_23_0_),
            .carryout(\nx.n10437 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_18_lut_LC_3_23_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_18_lut_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_18_lut_LC_3_23_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_18_lut_LC_3_23_1  (
            .in0(N__21366),
            .in1(N__21360),
            .in2(N__21350),
            .in3(N__21321),
            .lcout(\nx.n12953 ),
            .ltout(),
            .carryin(\nx.n10437 ),
            .carryout(\nx.n10438 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_19_lut_LC_3_23_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_19_lut_LC_3_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_19_lut_LC_3_23_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_19_lut_LC_3_23_2  (
            .in0(N__21318),
            .in1(N__22737),
            .in2(N__22752),
            .in3(N__21312),
            .lcout(\nx.n12955 ),
            .ltout(),
            .carryin(\nx.n10438 ),
            .carryout(\nx.n10439 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_20_lut_LC_3_23_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_20_lut_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_20_lut_LC_3_23_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_20_lut_LC_3_23_3  (
            .in0(N__21309),
            .in1(N__23046),
            .in2(N__22788),
            .in3(N__21303),
            .lcout(\nx.n12957 ),
            .ltout(),
            .carryin(\nx.n10439 ),
            .carryout(\nx.n10440 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_21_lut_LC_3_23_4 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_21_lut_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_21_lut_LC_3_23_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_21_lut_LC_3_23_4  (
            .in0(N__21300),
            .in1(N__25124),
            .in2(N__25047),
            .in3(N__21294),
            .lcout(\nx.n12959 ),
            .ltout(),
            .carryin(\nx.n10440 ),
            .carryout(\nx.n10441 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_22_lut_LC_3_23_5 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_22_lut_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_22_lut_LC_3_23_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_22_lut_LC_3_23_5  (
            .in0(N__21291),
            .in1(N__24990),
            .in2(N__25179),
            .in3(N__21285),
            .lcout(\nx.n12961 ),
            .ltout(),
            .carryin(\nx.n10441 ),
            .carryout(\nx.n10442 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_22_THRU_CRY_0_LC_3_23_6 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_22_THRU_CRY_0_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_22_THRU_CRY_0_LC_3_23_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_22_THRU_CRY_0_LC_3_23_6  (
            .in0(_gnd_net_),
            .in1(N__45666),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10442 ),
            .carryout(\nx.n10442_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_22_THRU_CRY_1_LC_3_23_7 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_22_THRU_CRY_1_LC_3_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_22_THRU_CRY_1_LC_3_23_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_22_THRU_CRY_1_LC_3_23_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__45754),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10442_THRU_CRY_0_THRU_CO ),
            .carryout(\nx.n10442_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_23_lut_LC_3_24_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_23_lut_LC_3_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_23_lut_LC_3_24_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_23_lut_LC_3_24_0  (
            .in0(N__21651),
            .in1(N__22827),
            .in2(N__22974),
            .in3(N__21645),
            .lcout(\nx.n12963 ),
            .ltout(),
            .carryin(bfn_3_24_0_),
            .carryout(\nx.n10443 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_24_lut_LC_3_24_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_24_lut_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_24_lut_LC_3_24_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_24_lut_LC_3_24_1  (
            .in0(N__21642),
            .in1(N__24872),
            .in2(N__29262),
            .in3(N__21636),
            .lcout(\nx.n12965 ),
            .ltout(),
            .carryin(\nx.n10443 ),
            .carryout(\nx.n10444 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_25_lut_LC_3_24_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_25_lut_LC_3_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_25_lut_LC_3_24_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_25_lut_LC_3_24_2  (
            .in0(N__21633),
            .in1(N__21627),
            .in2(N__21612),
            .in3(N__21579),
            .lcout(\nx.n12967 ),
            .ltout(),
            .carryin(\nx.n10444 ),
            .carryout(\nx.n10445 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_26_lut_LC_3_24_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_26_lut_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_26_lut_LC_3_24_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_26_lut_LC_3_24_3  (
            .in0(N__21576),
            .in1(N__21567),
            .in2(N__21554),
            .in3(N__21528),
            .lcout(\nx.n12969 ),
            .ltout(),
            .carryin(\nx.n10445 ),
            .carryout(\nx.n10446 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_27_lut_LC_3_24_4 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_27_lut_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_27_lut_LC_3_24_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_27_lut_LC_3_24_4  (
            .in0(N__21525),
            .in1(N__23067),
            .in2(N__22815),
            .in3(N__21516),
            .lcout(\nx.n12971 ),
            .ltout(),
            .carryin(\nx.n10446 ),
            .carryout(\nx.n10447 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_28_lut_LC_3_24_5 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_28_lut_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_28_lut_LC_3_24_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_28_lut_LC_3_24_5  (
            .in0(N__21513),
            .in1(N__21507),
            .in2(N__21492),
            .in3(N__21465),
            .lcout(\nx.n12973 ),
            .ltout(),
            .carryin(\nx.n10447 ),
            .carryout(\nx.n10448 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_28_THRU_CRY_0_LC_3_24_6 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_28_THRU_CRY_0_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_28_THRU_CRY_0_LC_3_24_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_28_THRU_CRY_0_LC_3_24_6  (
            .in0(_gnd_net_),
            .in1(N__45635),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10448 ),
            .carryout(\nx.n10448_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_28_THRU_CRY_1_LC_3_24_7 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_28_THRU_CRY_1_LC_3_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_28_THRU_CRY_1_LC_3_24_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_28_THRU_CRY_1_LC_3_24_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__45750),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10448_THRU_CRY_0_THRU_CO ),
            .carryout(\nx.n10448_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_29_lut_LC_3_25_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_29_lut_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_29_lut_LC_3_25_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_29_lut_LC_3_25_0  (
            .in0(N__21801),
            .in1(N__21933),
            .in2(N__21675),
            .in3(N__21795),
            .lcout(\nx.n12975 ),
            .ltout(),
            .carryin(bfn_3_25_0_),
            .carryout(\nx.n10449 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_30_lut_LC_3_25_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_30_lut_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_30_lut_LC_3_25_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_30_lut_LC_3_25_1  (
            .in0(N__21792),
            .in1(N__23034),
            .in2(N__23097),
            .in3(N__21786),
            .lcout(\nx.n12977 ),
            .ltout(),
            .carryin(\nx.n10449 ),
            .carryout(\nx.n10450 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_31_lut_LC_3_25_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_31_lut_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_31_lut_LC_3_25_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_31_lut_LC_3_25_2  (
            .in0(N__21783),
            .in1(N__22662),
            .in2(N__22575),
            .in3(N__21777),
            .lcout(\nx.n12979 ),
            .ltout(),
            .carryin(\nx.n10450 ),
            .carryout(\nx.n10451 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_32_lut_LC_3_25_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_32_lut_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_32_lut_LC_3_25_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_32_lut_LC_3_25_3  (
            .in0(N__21774),
            .in1(N__22454),
            .in2(N__22473),
            .in3(N__21768),
            .lcout(\nx.n12981 ),
            .ltout(),
            .carryin(\nx.n10451 ),
            .carryout(\nx.n10452 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_33_lut_LC_3_25_4 .C_ON=1'b0;
    defparam \nx.sub_14_add_2_33_lut_LC_3_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_33_lut_LC_3_25_4 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \nx.sub_14_add_2_33_lut_LC_3_25_4  (
            .in0(N__21764),
            .in1(N__21738),
            .in2(N__21723),
            .in3(N__21714),
            .lcout(\nx.n7181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i27_LC_3_25_6 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i27_LC_3_25_6 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i27_LC_3_25_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i27_LC_3_25_6  (
            .in0(N__21942),
            .in1(N__21674),
            .in2(_gnd_net_),
            .in3(N__28876),
            .lcout(neo_pixel_transmitter_t0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48416),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i28_1_lut_LC_3_25_7 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i28_1_lut_LC_3_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i28_1_lut_LC_3_25_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i28_1_lut_LC_3_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21941),
            .lcout(\nx.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_2_lut_LC_3_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_2_lut_LC_3_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_2_lut_LC_3_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_2_lut_LC_3_26_0  (
            .in0(_gnd_net_),
            .in1(N__26162),
            .in2(_gnd_net_),
            .in3(N__21918),
            .lcout(\nx.n3077 ),
            .ltout(),
            .carryin(bfn_3_26_0_),
            .carryout(\nx.n10862 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_3_lut_LC_3_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_3_lut_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_3_lut_LC_3_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_3_lut_LC_3_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23485),
            .in3(N__21909),
            .lcout(\nx.n3076 ),
            .ltout(),
            .carryin(\nx.n10862 ),
            .carryout(\nx.n10863 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_4_lut_LC_3_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_4_lut_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_4_lut_LC_3_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_4_lut_LC_3_26_2  (
            .in0(_gnd_net_),
            .in1(N__45632),
            .in2(N__21906),
            .in3(N__21879),
            .lcout(\nx.n3075 ),
            .ltout(),
            .carryin(\nx.n10863 ),
            .carryout(\nx.n10864 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_5_lut_LC_3_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_5_lut_LC_3_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_5_lut_LC_3_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_5_lut_LC_3_26_3  (
            .in0(_gnd_net_),
            .in1(N__45090),
            .in2(N__21876),
            .in3(N__21843),
            .lcout(\nx.n3074 ),
            .ltout(),
            .carryin(\nx.n10864 ),
            .carryout(\nx.n10865 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_6_lut_LC_3_26_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_6_lut_LC_3_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_6_lut_LC_3_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_6_lut_LC_3_26_4  (
            .in0(_gnd_net_),
            .in1(N__45633),
            .in2(N__23193),
            .in3(N__21825),
            .lcout(\nx.n3073 ),
            .ltout(),
            .carryin(\nx.n10865 ),
            .carryout(\nx.n10866 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_7_lut_LC_3_26_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_7_lut_LC_3_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_7_lut_LC_3_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_7_lut_LC_3_26_5  (
            .in0(_gnd_net_),
            .in1(N__45091),
            .in2(N__23247),
            .in3(N__21816),
            .lcout(\nx.n3072 ),
            .ltout(),
            .carryin(\nx.n10866 ),
            .carryout(\nx.n10867 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_8_lut_LC_3_26_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_8_lut_LC_3_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_8_lut_LC_3_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_8_lut_LC_3_26_6  (
            .in0(_gnd_net_),
            .in1(N__45634),
            .in2(N__23601),
            .in3(N__21804),
            .lcout(\nx.n3071 ),
            .ltout(),
            .carryin(\nx.n10867 ),
            .carryout(\nx.n10868 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_9_lut_LC_3_26_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_9_lut_LC_3_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_9_lut_LC_3_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_9_lut_LC_3_26_7  (
            .in0(_gnd_net_),
            .in1(N__45092),
            .in2(N__31734),
            .in3(N__22110),
            .lcout(\nx.n3070 ),
            .ltout(),
            .carryin(\nx.n10868 ),
            .carryout(\nx.n10869 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_10_lut_LC_3_27_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_10_lut_LC_3_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_10_lut_LC_3_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_10_lut_LC_3_27_0  (
            .in0(_gnd_net_),
            .in1(N__45392),
            .in2(N__23535),
            .in3(N__22095),
            .lcout(\nx.n3069 ),
            .ltout(),
            .carryin(bfn_3_27_0_),
            .carryout(\nx.n10870 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_11_lut_LC_3_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_11_lut_LC_3_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_11_lut_LC_3_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_11_lut_LC_3_27_1  (
            .in0(_gnd_net_),
            .in1(N__45399),
            .in2(N__22092),
            .in3(N__22053),
            .lcout(\nx.n3068 ),
            .ltout(),
            .carryin(\nx.n10870 ),
            .carryout(\nx.n10871 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_12_lut_LC_3_27_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_12_lut_LC_3_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_12_lut_LC_3_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_12_lut_LC_3_27_2  (
            .in0(_gnd_net_),
            .in1(N__45393),
            .in2(N__23391),
            .in3(N__22041),
            .lcout(\nx.n3067 ),
            .ltout(),
            .carryin(\nx.n10871 ),
            .carryout(\nx.n10872 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_13_lut_LC_3_27_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_13_lut_LC_3_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_13_lut_LC_3_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_13_lut_LC_3_27_3  (
            .in0(_gnd_net_),
            .in1(N__45400),
            .in2(N__22038),
            .in3(N__21999),
            .lcout(\nx.n3066 ),
            .ltout(),
            .carryin(\nx.n10872 ),
            .carryout(\nx.n10873 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_14_lut_LC_3_27_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_14_lut_LC_3_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_14_lut_LC_3_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_14_lut_LC_3_27_4  (
            .in0(_gnd_net_),
            .in1(N__45394),
            .in2(N__23160),
            .in3(N__21984),
            .lcout(\nx.n3065 ),
            .ltout(),
            .carryin(\nx.n10873 ),
            .carryout(\nx.n10874 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_15_lut_LC_3_27_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_15_lut_LC_3_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_15_lut_LC_3_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_15_lut_LC_3_27_5  (
            .in0(_gnd_net_),
            .in1(N__45401),
            .in2(N__23318),
            .in3(N__21966),
            .lcout(\nx.n3064 ),
            .ltout(),
            .carryin(\nx.n10874 ),
            .carryout(\nx.n10875 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_16_lut_LC_3_27_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_16_lut_LC_3_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_16_lut_LC_3_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_16_lut_LC_3_27_6  (
            .in0(_gnd_net_),
            .in1(N__45395),
            .in2(N__23355),
            .in3(N__21948),
            .lcout(\nx.n3063 ),
            .ltout(),
            .carryin(\nx.n10875 ),
            .carryout(\nx.n10876 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_17_lut_LC_3_27_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_17_lut_LC_3_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_17_lut_LC_3_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_17_lut_LC_3_27_7  (
            .in0(_gnd_net_),
            .in1(N__27503),
            .in2(N__45670),
            .in3(N__21945),
            .lcout(\nx.n3062 ),
            .ltout(),
            .carryin(\nx.n10876 ),
            .carryout(\nx.n10877 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_18_lut_LC_3_28_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_18_lut_LC_3_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_18_lut_LC_3_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_18_lut_LC_3_28_0  (
            .in0(_gnd_net_),
            .in1(N__23729),
            .in2(N__45631),
            .in3(N__22179),
            .lcout(\nx.n3061 ),
            .ltout(),
            .carryin(bfn_3_28_0_),
            .carryout(\nx.n10878 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_19_lut_LC_3_28_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_19_lut_LC_3_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_19_lut_LC_3_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_19_lut_LC_3_28_1  (
            .in0(_gnd_net_),
            .in1(N__45322),
            .in2(N__25848),
            .in3(N__22176),
            .lcout(\nx.n3060 ),
            .ltout(),
            .carryin(\nx.n10878 ),
            .carryout(\nx.n10879 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_20_lut_LC_3_28_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_20_lut_LC_3_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_20_lut_LC_3_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_20_lut_LC_3_28_2  (
            .in0(_gnd_net_),
            .in1(N__45504),
            .in2(N__23846),
            .in3(N__22167),
            .lcout(\nx.n3059 ),
            .ltout(),
            .carryin(\nx.n10879 ),
            .carryout(\nx.n10880 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_21_lut_LC_3_28_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_21_lut_LC_3_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_21_lut_LC_3_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_21_lut_LC_3_28_3  (
            .in0(_gnd_net_),
            .in1(N__45323),
            .in2(N__23709),
            .in3(N__22164),
            .lcout(\nx.n3058 ),
            .ltout(),
            .carryin(\nx.n10880 ),
            .carryout(\nx.n10881 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_22_lut_LC_3_28_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_22_lut_LC_3_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_22_lut_LC_3_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_22_lut_LC_3_28_4  (
            .in0(_gnd_net_),
            .in1(N__45505),
            .in2(N__24057),
            .in3(N__22161),
            .lcout(\nx.n3057 ),
            .ltout(),
            .carryin(\nx.n10881 ),
            .carryout(\nx.n10882 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_23_lut_LC_3_28_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_23_lut_LC_3_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_23_lut_LC_3_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_23_lut_LC_3_28_5  (
            .in0(_gnd_net_),
            .in1(N__45324),
            .in2(N__23817),
            .in3(N__22158),
            .lcout(\nx.n3056 ),
            .ltout(),
            .carryin(\nx.n10882 ),
            .carryout(\nx.n10883 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_24_lut_LC_3_28_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_24_lut_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_24_lut_LC_3_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_24_lut_LC_3_28_6  (
            .in0(_gnd_net_),
            .in1(N__45506),
            .in2(N__23577),
            .in3(N__22143),
            .lcout(\nx.n3055 ),
            .ltout(),
            .carryin(\nx.n10883 ),
            .carryout(\nx.n10884 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_25_lut_LC_3_28_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_25_lut_LC_3_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_25_lut_LC_3_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_25_lut_LC_3_28_7  (
            .in0(_gnd_net_),
            .in1(N__45325),
            .in2(N__23282),
            .in3(N__22128),
            .lcout(\nx.n3054 ),
            .ltout(),
            .carryin(\nx.n10884 ),
            .carryout(\nx.n10885 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_26_lut_LC_3_29_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_26_lut_LC_3_29_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_26_lut_LC_3_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_26_lut_LC_3_29_0  (
            .in0(_gnd_net_),
            .in1(N__23456),
            .in2(N__45630),
            .in3(N__22296),
            .lcout(\nx.n3053 ),
            .ltout(),
            .carryin(bfn_3_29_0_),
            .carryout(\nx.n10886 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_27_lut_LC_3_29_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_27_lut_LC_3_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_27_lut_LC_3_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2076_27_lut_LC_3_29_1  (
            .in0(_gnd_net_),
            .in1(N__45317),
            .in2(N__23126),
            .in3(N__22287),
            .lcout(\nx.n3052 ),
            .ltout(),
            .carryin(\nx.n10886 ),
            .carryout(\nx.n10887 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_28_lut_LC_3_29_2 .C_ON=1'b0;
    defparam \nx.mod_5_add_2076_28_lut_LC_3_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_28_lut_LC_3_29_2 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_2076_28_lut_LC_3_29_2  (
            .in0(N__45318),
            .in1(N__25605),
            .in2(N__27465),
            .in3(N__22284),
            .lcout(\nx.n3083 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_138_LC_3_29_6 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_138_LC_3_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_138_LC_3_29_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_138_LC_3_29_6  (
            .in0(N__24968),
            .in1(N__31003),
            .in2(N__26559),
            .in3(N__36895),
            .lcout(\nx.n45_adj_707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2_3_lut_adj_36_LC_3_30_1 .C_ON=1'b0;
    defparam \nx.i2_3_lut_adj_36_LC_3_30_1 .SEQ_MODE=4'b0000;
    defparam \nx.i2_3_lut_adj_36_LC_3_30_1 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i2_3_lut_adj_36_LC_3_30_1  (
            .in0(_gnd_net_),
            .in1(N__32708),
            .in2(N__22516),
            .in3(N__22202),
            .lcout(),
            .ltout(\nx.n11_adj_628_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8_4_lut_LC_3_30_2 .C_ON=1'b0;
    defparam \nx.i8_4_lut_LC_3_30_2 .SEQ_MODE=4'b0000;
    defparam \nx.i8_4_lut_LC_3_30_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i8_4_lut_LC_3_30_2  (
            .in0(N__24653),
            .in1(N__24635),
            .in2(N__22251),
            .in3(N__22248),
            .lcout(\nx.n1334 ),
            .ltout(\nx.n1334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i945_3_lut_LC_3_30_3 .C_ON=1'b0;
    defparam \nx.mod_5_i945_3_lut_LC_3_30_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i945_3_lut_LC_3_30_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i945_3_lut_LC_3_30_3  (
            .in0(N__22242),
            .in1(_gnd_net_),
            .in2(N__22224),
            .in3(N__22221),
            .lcout(\nx.n1406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i880_3_lut_LC_3_30_4 .C_ON=1'b0;
    defparam \nx.mod_5_i880_3_lut_LC_3_30_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i880_3_lut_LC_3_30_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i880_3_lut_LC_3_30_4  (
            .in0(N__24533),
            .in1(N__22215),
            .in2(_gnd_net_),
            .in3(N__22364),
            .lcout(\nx.n1309 ),
            .ltout(\nx.n1309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i947_3_lut_LC_3_30_5 .C_ON=1'b0;
    defparam \nx.mod_5_i947_3_lut_LC_3_30_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i947_3_lut_LC_3_30_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i947_3_lut_LC_3_30_5  (
            .in0(_gnd_net_),
            .in1(N__22188),
            .in2(N__22182),
            .in3(N__24587),
            .lcout(\nx.n1408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i875_3_lut_LC_3_30_6 .C_ON=1'b0;
    defparam \nx.mod_5_i875_3_lut_LC_3_30_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i875_3_lut_LC_3_30_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i875_3_lut_LC_3_30_6  (
            .in0(_gnd_net_),
            .in1(N__22416),
            .in2(N__22404),
            .in3(N__22365),
            .lcout(\nx.n1304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i948_3_lut_LC_3_30_7 .C_ON=1'b0;
    defparam \nx.mod_5_i948_3_lut_LC_3_30_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i948_3_lut_LC_3_30_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i948_3_lut_LC_3_30_7  (
            .in0(N__22335),
            .in1(N__32709),
            .in2(_gnd_net_),
            .in3(N__24586),
            .lcout(\nx.n1409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_2_lut_LC_3_31_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_2_lut_LC_3_31_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_2_lut_LC_3_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_2_lut_LC_3_31_0  (
            .in0(_gnd_net_),
            .in1(N__24970),
            .in2(_gnd_net_),
            .in3(N__22329),
            .lcout(\nx.n1477 ),
            .ltout(),
            .carryin(bfn_3_31_0_),
            .carryout(\nx.n10582 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_3_lut_LC_3_31_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_3_lut_LC_3_31_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_3_lut_LC_3_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_3_lut_LC_3_31_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28247),
            .in3(N__22326),
            .lcout(\nx.n1476 ),
            .ltout(),
            .carryin(\nx.n10582 ),
            .carryout(\nx.n10583 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_4_lut_LC_3_31_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_4_lut_LC_3_31_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_4_lut_LC_3_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_4_lut_LC_3_31_2  (
            .in0(_gnd_net_),
            .in1(N__44926),
            .in2(N__26791),
            .in3(N__22323),
            .lcout(\nx.n1475 ),
            .ltout(),
            .carryin(\nx.n10583 ),
            .carryout(\nx.n10584 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_5_lut_LC_3_31_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_5_lut_LC_3_31_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_5_lut_LC_3_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_5_lut_LC_3_31_3  (
            .in0(_gnd_net_),
            .in1(N__44929),
            .in2(N__26850),
            .in3(N__22320),
            .lcout(\nx.n1474 ),
            .ltout(),
            .carryin(\nx.n10584 ),
            .carryout(\nx.n10585 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_6_lut_LC_3_31_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_6_lut_LC_3_31_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_6_lut_LC_3_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_6_lut_LC_3_31_4  (
            .in0(_gnd_net_),
            .in1(N__44927),
            .in2(N__26677),
            .in3(N__22317),
            .lcout(\nx.n1473 ),
            .ltout(),
            .carryin(\nx.n10585 ),
            .carryout(\nx.n10586 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_7_lut_LC_3_31_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_7_lut_LC_3_31_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_7_lut_LC_3_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_7_lut_LC_3_31_5  (
            .in0(_gnd_net_),
            .in1(N__44930),
            .in2(N__26721),
            .in3(N__22314),
            .lcout(\nx.n1472 ),
            .ltout(),
            .carryin(\nx.n10586 ),
            .carryout(\nx.n10587 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_8_lut_LC_3_31_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_8_lut_LC_3_31_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_8_lut_LC_3_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_8_lut_LC_3_31_6  (
            .in0(_gnd_net_),
            .in1(N__44928),
            .in2(N__24489),
            .in3(N__22311),
            .lcout(\nx.n1471 ),
            .ltout(),
            .carryin(\nx.n10587 ),
            .carryout(\nx.n10588 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_9_lut_LC_3_31_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_9_lut_LC_3_31_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_9_lut_LC_3_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_9_lut_LC_3_31_7  (
            .in0(_gnd_net_),
            .in1(N__44931),
            .in2(N__26462),
            .in3(N__22533),
            .lcout(\nx.n1470 ),
            .ltout(),
            .carryin(\nx.n10588 ),
            .carryout(\nx.n10589 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_10_lut_LC_3_32_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_10_lut_LC_3_32_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_10_lut_LC_3_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_10_lut_LC_3_32_0  (
            .in0(_gnd_net_),
            .in1(N__44828),
            .in2(N__24903),
            .in3(N__22530),
            .lcout(\nx.n1469 ),
            .ltout(),
            .carryin(bfn_3_32_0_),
            .carryout(\nx.n10590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_11_lut_LC_3_32_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_11_lut_LC_3_32_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_11_lut_LC_3_32_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_11_lut_LC_3_32_1  (
            .in0(_gnd_net_),
            .in1(N__26761),
            .in2(N__45279),
            .in3(N__22527),
            .lcout(\nx.n1468 ),
            .ltout(),
            .carryin(\nx.n10590 ),
            .carryout(\nx.n10591 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_12_lut_LC_3_32_2 .C_ON=1'b0;
    defparam \nx.mod_5_add_1004_12_lut_LC_3_32_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_12_lut_LC_3_32_2 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1004_12_lut_LC_3_32_2  (
            .in0(N__44832),
            .in1(N__22482),
            .in2(N__28203),
            .in3(N__22524),
            .lcout(\nx.n1499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i941_3_lut_LC_3_32_4 .C_ON=1'b0;
    defparam \nx.mod_5_i941_3_lut_LC_3_32_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i941_3_lut_LC_3_32_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i941_3_lut_LC_3_32_4  (
            .in0(_gnd_net_),
            .in1(N__22521),
            .in2(N__22491),
            .in3(N__24590),
            .lcout(\nx.n1402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_4_lut_adj_37_LC_3_32_5 .C_ON=1'b0;
    defparam \nx.i6_4_lut_adj_37_LC_3_32_5 .SEQ_MODE=4'b0000;
    defparam \nx.i6_4_lut_adj_37_LC_3_32_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i6_4_lut_adj_37_LC_3_32_5  (
            .in0(N__22481),
            .in1(N__26455),
            .in2(N__26765),
            .in3(N__24898),
            .lcout(\nx.n16_adj_629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i31_1_lut_LC_4_16_0 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i31_1_lut_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i31_1_lut_LC_4_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i31_1_lut_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22424),
            .lcout(\nx.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i30_LC_4_16_4 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i30_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i30_LC_4_16_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i30_LC_4_16_4  (
            .in0(N__22455),
            .in1(N__22425),
            .in2(_gnd_net_),
            .in3(N__28842),
            .lcout(neo_pixel_transmitter_t0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48399),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i15_LC_4_17_1.C_ON=1'b0;
    defparam neopxl_color_prev_i15_LC_4_17_1.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i15_LC_4_17_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 neopxl_color_prev_i15_LC_4_17_1 (
            .in0(N__26651),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(neopxl_color_prev_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48388),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i3_1_lut_LC_4_17_3 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i3_1_lut_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i3_1_lut_LC_4_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i3_1_lut_LC_4_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22673),
            .lcout(\nx.n31_adj_650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i18_1_lut_LC_4_17_5 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i18_1_lut_LC_4_17_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i18_1_lut_LC_4_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i18_1_lut_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22706),
            .lcout(\nx.n16_adj_661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i17_LC_4_17_6 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i17_LC_4_17_6 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i17_LC_4_17_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i17_LC_4_17_6  (
            .in0(_gnd_net_),
            .in1(N__28843),
            .in2(N__22710),
            .in3(N__22736),
            .lcout(neo_pixel_transmitter_t0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48388),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i2_LC_4_17_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i2_LC_4_17_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i2_LC_4_17_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i2_LC_4_17_7  (
            .in0(N__22674),
            .in1(N__22694),
            .in2(N__28873),
            .in3(_gnd_net_),
            .lcout(neo_pixel_transmitter_t0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48388),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_18_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_18_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_18_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_18_0  (
            .in0(N__28833),
            .in1(N__22661),
            .in2(_gnd_net_),
            .in3(N__22584),
            .lcout(neo_pixel_transmitter_t0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48400),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i9_LC_4_18_2 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i9_LC_4_18_2 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i9_LC_4_18_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i9_LC_4_18_2  (
            .in0(N__28834),
            .in1(N__22631),
            .in2(_gnd_net_),
            .in3(N__25086),
            .lcout(neo_pixel_transmitter_t0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48400),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i11_1_lut_LC_4_18_3 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i11_1_lut_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i11_1_lut_LC_4_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i11_1_lut_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22611),
            .lcout(\nx.n23_adj_617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i30_1_lut_LC_4_18_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i30_1_lut_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i30_1_lut_LC_4_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i30_1_lut_LC_4_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22583),
            .lcout(\nx.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i11_LC_4_18_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i11_LC_4_18_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i11_LC_4_18_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i11_LC_4_18_7  (
            .in0(N__22553),
            .in1(N__28835),
            .in2(_gnd_net_),
            .in3(N__22923),
            .lcout(neo_pixel_transmitter_t0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48400),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i21_LC_4_19_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i21_LC_4_19_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i21_LC_4_19_0 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i21_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(N__28850),
            .in2(N__22839),
            .in3(N__22970),
            .lcout(neo_pixel_transmitter_t0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_1 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_1 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_1  (
            .in0(N__22899),
            .in1(N__22943),
            .in2(_gnd_net_),
            .in3(N__28855),
            .lcout(neo_pixel_transmitter_t0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i12_1_lut_LC_4_19_3 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i12_1_lut_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i12_1_lut_LC_4_19_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \nx.sub_14_inv_0_i12_1_lut_LC_4_19_3  (
            .in0(N__22922),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\nx.n22_adj_618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i14_1_lut_LC_4_19_4 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i14_1_lut_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i14_1_lut_LC_4_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i14_1_lut_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22898),
            .lcout(\nx.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i7_LC_4_19_5 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i7_LC_4_19_5 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i7_LC_4_19_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i7_LC_4_19_5  (
            .in0(N__23214),
            .in1(N__22877),
            .in2(_gnd_net_),
            .in3(N__28856),
            .lcout(neo_pixel_transmitter_t0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48404),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9312_3_lut_LC_4_19_6 .C_ON=1'b0;
    defparam \nx.i9312_3_lut_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9312_3_lut_LC_4_19_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \nx.i9312_3_lut_LC_4_19_6  (
            .in0(N__26647),
            .in1(N__23979),
            .in2(_gnd_net_),
            .in3(N__43160),
            .lcout(\nx.n13159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i22_1_lut_LC_4_19_7 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i22_1_lut_LC_4_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i22_1_lut_LC_4_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i22_1_lut_LC_4_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22835),
            .lcout(\nx.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_0  (
            .in0(_gnd_net_),
            .in1(N__22808),
            .in2(N__23079),
            .in3(N__28851),
            .lcout(neo_pixel_transmitter_t0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48408),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i18_LC_4_20_1 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i18_LC_4_20_1 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i18_LC_4_20_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i18_LC_4_20_1  (
            .in0(N__23055),
            .in1(N__22784),
            .in2(N__28875),
            .in3(_gnd_net_),
            .lcout(neo_pixel_transmitter_t0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48408),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i29_1_lut_LC_4_20_2 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i29_1_lut_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i29_1_lut_LC_4_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i29_1_lut_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23006),
            .lcout(\nx.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i26_1_lut_LC_4_20_3 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i26_1_lut_LC_4_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i26_1_lut_LC_4_20_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \nx.sub_14_inv_0_i26_1_lut_LC_4_20_3  (
            .in0(_gnd_net_),
            .in1(N__23075),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\nx.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i19_1_lut_LC_4_20_4 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i19_1_lut_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i19_1_lut_LC_4_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i19_1_lut_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23054),
            .lcout(\nx.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i28_LC_4_20_5 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i28_LC_4_20_5 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i28_LC_4_20_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i28_LC_4_20_5  (
            .in0(N__23030),
            .in1(_gnd_net_),
            .in2(N__23010),
            .in3(N__28878),
            .lcout(neo_pixel_transmitter_t0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48408),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_86_LC_4_20_7 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_86_LC_4_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_86_LC_4_20_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_86_LC_4_20_7  (
            .in0(N__25372),
            .in1(N__31906),
            .in2(N__30368),
            .in3(N__25492),
            .lcout(\nx.n43_adj_677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_93_LC_4_21_0 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_93_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_93_LC_4_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_93_LC_4_21_0  (
            .in0(N__23182),
            .in1(N__23143),
            .in2(N__23311),
            .in3(N__23233),
            .lcout(\nx.n44_adj_681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2022_3_lut_LC_4_21_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2022_3_lut_LC_4_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2022_3_lut_LC_4_21_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2022_3_lut_LC_4_21_1  (
            .in0(_gnd_net_),
            .in1(N__25452),
            .in2(N__25470),
            .in3(N__31858),
            .lcout(\nx.n2995 ),
            .ltout(\nx.n2995_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_3_lut_adj_94_LC_4_21_2 .C_ON=1'b0;
    defparam \nx.i7_3_lut_adj_94_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i7_3_lut_adj_94_LC_4_21_2 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i7_3_lut_adj_94_LC_4_21_2  (
            .in0(_gnd_net_),
            .in1(N__26171),
            .in2(N__22998),
            .in3(N__23492),
            .lcout(),
            .ltout(\nx.n33_adj_682_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i22_4_lut_adj_98_LC_4_21_3 .C_ON=1'b0;
    defparam \nx.i22_4_lut_adj_98_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.i22_4_lut_adj_98_LC_4_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i22_4_lut_adj_98_LC_4_21_3  (
            .in0(N__22995),
            .in1(N__23386),
            .in2(N__22989),
            .in3(N__31732),
            .lcout(\nx.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2032_3_lut_LC_4_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2032_3_lut_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2032_3_lut_LC_4_21_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2032_3_lut_LC_4_21_4  (
            .in0(_gnd_net_),
            .in1(N__25326),
            .in2(N__31875),
            .in3(N__25346),
            .lcout(\nx.n3005 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i8_1_lut_LC_4_21_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i8_1_lut_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i8_1_lut_LC_4_21_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \nx.sub_14_inv_0_i8_1_lut_LC_4_21_6  (
            .in0(N__23213),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\nx.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9508_3_lut_LC_4_21_7 .C_ON=1'b0;
    defparam \nx.i9508_3_lut_LC_4_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.i9508_3_lut_LC_4_21_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.i9508_3_lut_LC_4_21_7  (
            .in0(_gnd_net_),
            .in1(N__25356),
            .in2(N__25382),
            .in3(N__31854),
            .lcout(\nx.n3006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2013_3_lut_LC_4_22_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2013_3_lut_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2013_3_lut_LC_4_22_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \nx.mod_5_i2013_3_lut_LC_4_22_0  (
            .in0(N__25632),
            .in1(N__31838),
            .in2(_gnd_net_),
            .in3(N__29589),
            .lcout(\nx.n2986 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1958_3_lut_LC_4_22_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1958_3_lut_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1958_3_lut_LC_4_22_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1958_3_lut_LC_4_22_1  (
            .in0(_gnd_net_),
            .in1(N__27173),
            .in2(N__27147),
            .in3(N__30301),
            .lcout(\nx.n2899 ),
            .ltout(\nx.n2899_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9504_3_lut_LC_4_22_2 .C_ON=1'b0;
    defparam \nx.i9504_3_lut_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9504_3_lut_LC_4_22_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.i9504_3_lut_LC_4_22_2  (
            .in0(_gnd_net_),
            .in1(N__31837),
            .in2(N__23163),
            .in3(N__25548),
            .lcout(\nx.n2998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1953_3_lut_LC_4_22_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1953_3_lut_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1953_3_lut_LC_4_22_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1953_3_lut_LC_4_22_3  (
            .in0(_gnd_net_),
            .in1(N__27285),
            .in2(N__27258),
            .in3(N__30302),
            .lcout(\nx.n2894 ),
            .ltout(\nx.n2894_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_87_LC_4_22_4 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_87_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_87_LC_4_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_87_LC_4_22_4  (
            .in0(N__29650),
            .in1(N__27543),
            .in2(N__23130),
            .in3(N__29518),
            .lcout(\nx.n40_adj_678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2012_3_lut_LC_4_22_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2012_3_lut_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2012_3_lut_LC_4_22_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i2012_3_lut_LC_4_22_6  (
            .in0(_gnd_net_),
            .in1(N__31839),
            .in2(N__29967),
            .in3(N__25620),
            .lcout(\nx.n2985 ),
            .ltout(\nx.n2985_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_95_LC_4_22_7 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_95_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_95_LC_4_22_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_95_LC_4_22_7  (
            .in0(N__25601),
            .in1(N__23263),
            .in2(N__23463),
            .in3(N__23443),
            .lcout(\nx.n40_adj_683 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i22_4_lut_adj_92_LC_4_23_0 .C_ON=1'b0;
    defparam \nx.i22_4_lut_adj_92_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.i22_4_lut_adj_92_LC_4_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i22_4_lut_adj_92_LC_4_23_0  (
            .in0(N__29450),
            .in1(N__29707),
            .in2(N__23415),
            .in3(N__23361),
            .lcout(),
            .ltout(\nx.n47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i24_4_lut_LC_4_23_1 .C_ON=1'b0;
    defparam \nx.i24_4_lut_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.i24_4_lut_LC_4_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i24_4_lut_LC_4_23_1  (
            .in0(N__25221),
            .in1(N__23403),
            .in2(N__23397),
            .in3(N__30462),
            .lcout(\nx.n2918 ),
            .ltout(\nx.n2918_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2027_3_lut_LC_4_23_2 .C_ON=1'b0;
    defparam \nx.mod_5_i2027_3_lut_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2027_3_lut_LC_4_23_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2027_3_lut_LC_4_23_2  (
            .in0(_gnd_net_),
            .in1(N__25245),
            .in2(N__23394),
            .in3(N__25268),
            .lcout(\nx.n3000 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_3_lut_LC_4_23_3 .C_ON=1'b0;
    defparam \nx.i13_3_lut_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.i13_3_lut_LC_4_23_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \nx.i13_3_lut_LC_4_23_3  (
            .in0(_gnd_net_),
            .in1(N__27579),
            .in2(N__30409),
            .in3(N__29956),
            .lcout(\nx.n38_adj_676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2023_3_lut_LC_4_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2023_3_lut_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2023_3_lut_LC_4_23_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i2023_3_lut_LC_4_23_4  (
            .in0(N__31834),
            .in1(_gnd_net_),
            .in2(N__25506),
            .in3(N__25479),
            .lcout(\nx.n2996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9502_3_lut_LC_4_23_5 .C_ON=1'b0;
    defparam \nx.i9502_3_lut_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9502_3_lut_LC_4_23_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.i9502_3_lut_LC_4_23_5  (
            .in0(N__25538),
            .in1(_gnd_net_),
            .in2(N__25518),
            .in3(N__31833),
            .lcout(\nx.n2997 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2018_3_lut_LC_4_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2018_3_lut_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2018_3_lut_LC_4_23_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.mod_5_i2018_3_lut_LC_4_23_6  (
            .in0(N__31836),
            .in1(N__29528),
            .in2(_gnd_net_),
            .in3(N__25680),
            .lcout(\nx.n2991 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2014_3_lut_LC_4_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i2014_3_lut_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2014_3_lut_LC_4_23_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2014_3_lut_LC_4_23_7  (
            .in0(_gnd_net_),
            .in1(N__25641),
            .in2(N__30495),
            .in3(N__31835),
            .lcout(\nx.n2987 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9506_3_lut_LC_4_24_0 .C_ON=1'b0;
    defparam \nx.i9506_3_lut_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.i9506_3_lut_LC_4_24_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.i9506_3_lut_LC_4_24_0  (
            .in0(_gnd_net_),
            .in1(N__25317),
            .in2(N__31863),
            .in3(N__29451),
            .lcout(\nx.n3004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2029_3_lut_LC_4_24_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2029_3_lut_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2029_3_lut_LC_4_24_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2029_3_lut_LC_4_24_1  (
            .in0(_gnd_net_),
            .in1(N__30361),
            .in2(N__25302),
            .in3(N__31822),
            .lcout(\nx.n3002 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2016_3_lut_LC_4_24_2 .C_ON=1'b0;
    defparam \nx.mod_5_i2016_3_lut_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2016_3_lut_LC_4_24_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i2016_3_lut_LC_4_24_2  (
            .in0(N__29571),
            .in1(_gnd_net_),
            .in2(N__31865),
            .in3(N__25659),
            .lcout(\nx.n2989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2017_3_lut_LC_4_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2017_3_lut_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2017_3_lut_LC_4_24_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2017_3_lut_LC_4_24_3  (
            .in0(_gnd_net_),
            .in1(N__27542),
            .in2(N__25671),
            .in3(N__31826),
            .lcout(\nx.n2990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2015_3_lut_LC_4_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2015_3_lut_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2015_3_lut_LC_4_24_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2015_3_lut_LC_4_24_4  (
            .in0(_gnd_net_),
            .in1(N__30144),
            .in2(N__31866),
            .in3(N__25650),
            .lcout(\nx.n2988 ),
            .ltout(\nx.n2988_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_100_LC_4_24_5 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_100_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_100_LC_4_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_100_LC_4_24_5  (
            .in0(N__24043),
            .in1(N__23695),
            .in2(N__23550),
            .in3(N__23803),
            .lcout(\nx.n41_adj_686 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2021_3_lut_LC_4_24_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2021_3_lut_LC_4_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2021_3_lut_LC_4_24_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2021_3_lut_LC_4_24_6  (
            .in0(_gnd_net_),
            .in1(N__25440),
            .in2(N__31864),
            .in3(N__29874),
            .lcout(\nx.n2994 ),
            .ltout(\nx.n2994_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_97_LC_4_24_7 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_97_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_97_LC_4_24_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_97_LC_4_24_7  (
            .in0(N__23828),
            .in1(N__25841),
            .in2(N__23538),
            .in3(N__23521),
            .lcout(\nx.n42_adj_684 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2036_3_lut_LC_4_25_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2036_3_lut_LC_4_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2036_3_lut_LC_4_25_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i2036_3_lut_LC_4_25_0  (
            .in0(N__25212),
            .in1(N__26134),
            .in2(_gnd_net_),
            .in3(N__31859),
            .lcout(\nx.n3009 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2019_3_lut_LC_4_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2019_3_lut_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2019_3_lut_LC_4_25_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2019_3_lut_LC_4_25_1  (
            .in0(_gnd_net_),
            .in1(N__29652),
            .in2(N__31876),
            .in3(N__25428),
            .lcout(\nx.n2992 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2083_3_lut_LC_4_25_2 .C_ON=1'b0;
    defparam \nx.mod_5_i2083_3_lut_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2083_3_lut_LC_4_25_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i2083_3_lut_LC_4_25_2  (
            .in0(N__27456),
            .in1(_gnd_net_),
            .in2(N__23813),
            .in3(N__23787),
            .lcout(\nx.n3088 ),
            .ltout(\nx.n3088_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_104_LC_4_25_3 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_104_LC_4_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_104_LC_4_25_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_104_LC_4_25_3  (
            .in0(N__24004),
            .in1(N__23776),
            .in2(N__23751),
            .in3(N__24277),
            .lcout(\nx.n44_adj_690 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2088_3_lut_LC_4_25_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2088_3_lut_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2088_3_lut_LC_4_25_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2088_3_lut_LC_4_25_5  (
            .in0(_gnd_net_),
            .in1(N__23739),
            .in2(N__23730),
            .in3(N__27452),
            .lcout(\nx.n3093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2085_3_lut_LC_4_25_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2085_3_lut_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2085_3_lut_LC_4_25_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2085_3_lut_LC_4_25_6  (
            .in0(_gnd_net_),
            .in1(N__23705),
            .in2(N__27464),
            .in3(N__23682),
            .lcout(\nx.n3090 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_121_LC_4_25_7 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_121_LC_4_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_121_LC_4_25_7 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \nx.i1_4_lut_adj_121_LC_4_25_7  (
            .in0(N__23673),
            .in1(N__27311),
            .in2(N__24236),
            .in3(N__23661),
            .lcout(\nx.n12355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_122_LC_4_26_1 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_122_LC_4_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_122_LC_4_26_1 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \nx.i1_4_lut_adj_122_LC_4_26_1  (
            .in0(N__25733),
            .in1(N__24237),
            .in2(N__23652),
            .in3(N__23637),
            .lcout(),
            .ltout(\nx.n12357_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_123_LC_4_26_2 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_123_LC_4_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_123_LC_4_26_2 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \nx.i1_4_lut_adj_123_LC_4_26_2  (
            .in0(N__24238),
            .in1(N__25808),
            .in2(N__23631),
            .in3(N__23628),
            .lcout(),
            .ltout(\nx.n12359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_124_LC_4_26_3 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_124_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_124_LC_4_26_3 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \nx.i1_4_lut_adj_124_LC_4_26_3  (
            .in0(N__25794),
            .in1(N__23616),
            .in2(N__23604),
            .in3(N__24239),
            .lcout(),
            .ltout(\nx.n12361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_125_LC_4_26_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_125_LC_4_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_125_LC_4_26_4 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \nx.i1_4_lut_adj_125_LC_4_26_4  (
            .in0(N__24240),
            .in1(N__24303),
            .in2(N__24291),
            .in3(N__24281),
            .lcout(),
            .ltout(\nx.n12363_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_126_LC_4_26_5 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_126_LC_4_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_126_LC_4_26_5 .LUT_INIT=16'b1111101111111000;
    LogicCell40 \nx.i1_4_lut_adj_126_LC_4_26_5  (
            .in0(N__24261),
            .in1(N__24241),
            .in2(N__24249),
            .in3(N__24014),
            .lcout(),
            .ltout(\nx.n12365_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_127_LC_4_26_6 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_127_LC_4_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_127_LC_4_26_6 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \nx.i1_4_lut_adj_127_LC_4_26_6  (
            .in0(N__24242),
            .in1(N__24101),
            .in2(N__24087),
            .in3(N__24084),
            .lcout(\nx.n12367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2084_3_lut_LC_4_26_7 .C_ON=1'b0;
    defparam \nx.mod_5_i2084_3_lut_LC_4_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2084_3_lut_LC_4_26_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2084_3_lut_LC_4_26_7  (
            .in0(_gnd_net_),
            .in1(N__24053),
            .in2(N__24027),
            .in3(N__27463),
            .lcout(\nx.n3089 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.bit_ctr__i0_LC_4_27_0 .C_ON=1'b1;
    defparam \nx.bit_ctr__i0_LC_4_27_0 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i0_LC_4_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i0_LC_4_27_0  (
            .in0(_gnd_net_),
            .in1(N__23959),
            .in2(_gnd_net_),
            .in3(N__23943),
            .lcout(\nx.bit_ctr_0 ),
            .ltout(),
            .carryin(bfn_4_27_0_),
            .carryout(\nx.n10391 ),
            .clk(N__48423),
            .ce(N__24840),
            .sr(N__24768));
    defparam \nx.bit_ctr__i1_LC_4_27_1 .C_ON=1'b1;
    defparam \nx.bit_ctr__i1_LC_4_27_1 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i1_LC_4_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i1_LC_4_27_1  (
            .in0(_gnd_net_),
            .in1(N__23927),
            .in2(_gnd_net_),
            .in3(N__23916),
            .lcout(\nx.bit_ctr_1 ),
            .ltout(),
            .carryin(\nx.n10391 ),
            .carryout(\nx.n10392 ),
            .clk(N__48423),
            .ce(N__24840),
            .sr(N__24768));
    defparam \nx.bit_ctr__i2_LC_4_27_2 .C_ON=1'b1;
    defparam \nx.bit_ctr__i2_LC_4_27_2 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i2_LC_4_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i2_LC_4_27_2  (
            .in0(_gnd_net_),
            .in1(N__23903),
            .in2(_gnd_net_),
            .in3(N__23892),
            .lcout(\nx.bit_ctr_2 ),
            .ltout(),
            .carryin(\nx.n10392 ),
            .carryout(\nx.n10393 ),
            .clk(N__48423),
            .ce(N__24840),
            .sr(N__24768));
    defparam \nx.bit_ctr__i3_LC_4_27_3 .C_ON=1'b1;
    defparam \nx.bit_ctr__i3_LC_4_27_3 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i3_LC_4_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i3_LC_4_27_3  (
            .in0(_gnd_net_),
            .in1(N__23877),
            .in2(_gnd_net_),
            .in3(N__23850),
            .lcout(\nx.bit_ctr_3 ),
            .ltout(),
            .carryin(\nx.n10393 ),
            .carryout(\nx.n10394 ),
            .clk(N__48423),
            .ce(N__24840),
            .sr(N__24768));
    defparam \nx.bit_ctr__i4_LC_4_27_4 .C_ON=1'b1;
    defparam \nx.bit_ctr__i4_LC_4_27_4 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i4_LC_4_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i4_LC_4_27_4  (
            .in0(_gnd_net_),
            .in1(N__24356),
            .in2(_gnd_net_),
            .in3(N__24330),
            .lcout(\nx.bit_ctr_4 ),
            .ltout(),
            .carryin(\nx.n10394 ),
            .carryout(\nx.n10395 ),
            .clk(N__48423),
            .ce(N__24840),
            .sr(N__24768));
    defparam \nx.bit_ctr__i5_LC_4_27_5 .C_ON=1'b1;
    defparam \nx.bit_ctr__i5_LC_4_27_5 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i5_LC_4_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i5_LC_4_27_5  (
            .in0(_gnd_net_),
            .in1(N__26170),
            .in2(_gnd_net_),
            .in3(N__24327),
            .lcout(\nx.bit_ctr_5 ),
            .ltout(),
            .carryin(\nx.n10395 ),
            .carryout(\nx.n10396 ),
            .clk(N__48423),
            .ce(N__24840),
            .sr(N__24768));
    defparam \nx.bit_ctr__i6_LC_4_27_6 .C_ON=1'b1;
    defparam \nx.bit_ctr__i6_LC_4_27_6 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i6_LC_4_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i6_LC_4_27_6  (
            .in0(_gnd_net_),
            .in1(N__26119),
            .in2(_gnd_net_),
            .in3(N__24324),
            .lcout(\nx.bit_ctr_6 ),
            .ltout(),
            .carryin(\nx.n10396 ),
            .carryout(\nx.n10397 ),
            .clk(N__48423),
            .ce(N__24840),
            .sr(N__24768));
    defparam \nx.bit_ctr__i7_LC_4_27_7 .C_ON=1'b1;
    defparam \nx.bit_ctr__i7_LC_4_27_7 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i7_LC_4_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i7_LC_4_27_7  (
            .in0(_gnd_net_),
            .in1(N__29808),
            .in2(_gnd_net_),
            .in3(N__24321),
            .lcout(\nx.bit_ctr_7 ),
            .ltout(),
            .carryin(\nx.n10397 ),
            .carryout(\nx.n10398 ),
            .clk(N__48423),
            .ce(N__24840),
            .sr(N__24768));
    defparam \nx.bit_ctr__i8_LC_4_28_0 .C_ON=1'b1;
    defparam \nx.bit_ctr__i8_LC_4_28_0 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i8_LC_4_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i8_LC_4_28_0  (
            .in0(_gnd_net_),
            .in1(N__28523),
            .in2(_gnd_net_),
            .in3(N__24318),
            .lcout(\nx.bit_ctr_8 ),
            .ltout(),
            .carryin(bfn_4_28_0_),
            .carryout(\nx.n10399 ),
            .clk(N__48426),
            .ce(N__24844),
            .sr(N__24778));
    defparam \nx.bit_ctr__i9_LC_4_28_1 .C_ON=1'b1;
    defparam \nx.bit_ctr__i9_LC_4_28_1 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i9_LC_4_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i9_LC_4_28_1  (
            .in0(_gnd_net_),
            .in1(N__35881),
            .in2(_gnd_net_),
            .in3(N__24315),
            .lcout(\nx.bit_ctr_9 ),
            .ltout(),
            .carryin(\nx.n10399 ),
            .carryout(\nx.n10400 ),
            .clk(N__48426),
            .ce(N__24844),
            .sr(N__24778));
    defparam \nx.bit_ctr__i10_LC_4_28_2 .C_ON=1'b1;
    defparam \nx.bit_ctr__i10_LC_4_28_2 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i10_LC_4_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i10_LC_4_28_2  (
            .in0(_gnd_net_),
            .in1(N__37859),
            .in2(_gnd_net_),
            .in3(N__24312),
            .lcout(\nx.bit_ctr_10 ),
            .ltout(),
            .carryin(\nx.n10400 ),
            .carryout(\nx.n10401 ),
            .clk(N__48426),
            .ce(N__24844),
            .sr(N__24778));
    defparam \nx.bit_ctr__i11_LC_4_28_3 .C_ON=1'b1;
    defparam \nx.bit_ctr__i11_LC_4_28_3 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i11_LC_4_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i11_LC_4_28_3  (
            .in0(_gnd_net_),
            .in1(N__41258),
            .in2(_gnd_net_),
            .in3(N__24309),
            .lcout(\nx.bit_ctr_11 ),
            .ltout(),
            .carryin(\nx.n10401 ),
            .carryout(\nx.n10402 ),
            .clk(N__48426),
            .ce(N__24844),
            .sr(N__24778));
    defparam \nx.bit_ctr__i12_LC_4_28_4 .C_ON=1'b1;
    defparam \nx.bit_ctr__i12_LC_4_28_4 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i12_LC_4_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i12_LC_4_28_4  (
            .in0(_gnd_net_),
            .in1(N__43539),
            .in2(_gnd_net_),
            .in3(N__24306),
            .lcout(\nx.bit_ctr_12 ),
            .ltout(),
            .carryin(\nx.n10402 ),
            .carryout(\nx.n10403 ),
            .clk(N__48426),
            .ce(N__24844),
            .sr(N__24778));
    defparam \nx.bit_ctr__i13_LC_4_28_5 .C_ON=1'b1;
    defparam \nx.bit_ctr__i13_LC_4_28_5 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i13_LC_4_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i13_LC_4_28_5  (
            .in0(_gnd_net_),
            .in1(N__39828),
            .in2(_gnd_net_),
            .in3(N__24402),
            .lcout(\nx.bit_ctr_13 ),
            .ltout(),
            .carryin(\nx.n10403 ),
            .carryout(\nx.n10404 ),
            .clk(N__48426),
            .ce(N__24844),
            .sr(N__24778));
    defparam \nx.bit_ctr__i14_LC_4_28_6 .C_ON=1'b1;
    defparam \nx.bit_ctr__i14_LC_4_28_6 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i14_LC_4_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i14_LC_4_28_6  (
            .in0(_gnd_net_),
            .in1(N__36901),
            .in2(_gnd_net_),
            .in3(N__24399),
            .lcout(\nx.bit_ctr_14 ),
            .ltout(),
            .carryin(\nx.n10404 ),
            .carryout(\nx.n10405 ),
            .clk(N__48426),
            .ce(N__24844),
            .sr(N__24778));
    defparam \nx.bit_ctr__i15_LC_4_28_7 .C_ON=1'b1;
    defparam \nx.bit_ctr__i15_LC_4_28_7 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i15_LC_4_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i15_LC_4_28_7  (
            .in0(_gnd_net_),
            .in1(N__34064),
            .in2(_gnd_net_),
            .in3(N__24396),
            .lcout(\nx.bit_ctr_15 ),
            .ltout(),
            .carryin(\nx.n10405 ),
            .carryout(\nx.n10406 ),
            .clk(N__48426),
            .ce(N__24844),
            .sr(N__24778));
    defparam \nx.bit_ctr__i16_LC_4_29_0 .C_ON=1'b1;
    defparam \nx.bit_ctr__i16_LC_4_29_0 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i16_LC_4_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i16_LC_4_29_0  (
            .in0(_gnd_net_),
            .in1(N__30096),
            .in2(_gnd_net_),
            .in3(N__24393),
            .lcout(\nx.bit_ctr_16 ),
            .ltout(),
            .carryin(bfn_4_29_0_),
            .carryout(\nx.n10407 ),
            .clk(N__48432),
            .ce(N__24846),
            .sr(N__24783));
    defparam \nx.bit_ctr__i17_LC_4_29_1 .C_ON=1'b1;
    defparam \nx.bit_ctr__i17_LC_4_29_1 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i17_LC_4_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i17_LC_4_29_1  (
            .in0(_gnd_net_),
            .in1(N__32745),
            .in2(_gnd_net_),
            .in3(N__24390),
            .lcout(\nx.bit_ctr_17 ),
            .ltout(),
            .carryin(\nx.n10407 ),
            .carryout(\nx.n10408 ),
            .clk(N__48432),
            .ce(N__24846),
            .sr(N__24783));
    defparam \nx.bit_ctr__i18_LC_4_29_2 .C_ON=1'b1;
    defparam \nx.bit_ctr__i18_LC_4_29_2 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i18_LC_4_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i18_LC_4_29_2  (
            .in0(_gnd_net_),
            .in1(N__34952),
            .in2(_gnd_net_),
            .in3(N__24387),
            .lcout(\nx.bit_ctr_18 ),
            .ltout(),
            .carryin(\nx.n10408 ),
            .carryout(\nx.n10409 ),
            .clk(N__48432),
            .ce(N__24846),
            .sr(N__24783));
    defparam \nx.bit_ctr__i19_LC_4_29_3 .C_ON=1'b1;
    defparam \nx.bit_ctr__i19_LC_4_29_3 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i19_LC_4_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i19_LC_4_29_3  (
            .in0(_gnd_net_),
            .in1(N__30995),
            .in2(_gnd_net_),
            .in3(N__24384),
            .lcout(\nx.bit_ctr_19 ),
            .ltout(),
            .carryin(\nx.n10409 ),
            .carryout(\nx.n10410 ),
            .clk(N__48432),
            .ce(N__24846),
            .sr(N__24783));
    defparam \nx.bit_ctr__i20_LC_4_29_4 .C_ON=1'b1;
    defparam \nx.bit_ctr__i20_LC_4_29_4 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i20_LC_4_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i20_LC_4_29_4  (
            .in0(_gnd_net_),
            .in1(N__30836),
            .in2(_gnd_net_),
            .in3(N__24381),
            .lcout(\nx.bit_ctr_20 ),
            .ltout(),
            .carryin(\nx.n10410 ),
            .carryout(\nx.n10411 ),
            .clk(N__48432),
            .ce(N__24846),
            .sr(N__24783));
    defparam \nx.bit_ctr__i21_LC_4_29_5 .C_ON=1'b1;
    defparam \nx.bit_ctr__i21_LC_4_29_5 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i21_LC_4_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i21_LC_4_29_5  (
            .in0(_gnd_net_),
            .in1(N__24969),
            .in2(_gnd_net_),
            .in3(N__24378),
            .lcout(\nx.bit_ctr_21 ),
            .ltout(),
            .carryin(\nx.n10411 ),
            .carryout(\nx.n10412 ),
            .clk(N__48432),
            .ce(N__24846),
            .sr(N__24783));
    defparam \nx.bit_ctr__i22_LC_4_29_6 .C_ON=1'b1;
    defparam \nx.bit_ctr__i22_LC_4_29_6 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i22_LC_4_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i22_LC_4_29_6  (
            .in0(_gnd_net_),
            .in1(N__32710),
            .in2(_gnd_net_),
            .in3(N__24468),
            .lcout(\nx.bit_ctr_22 ),
            .ltout(),
            .carryin(\nx.n10412 ),
            .carryout(\nx.n10413 ),
            .clk(N__48432),
            .ce(N__24846),
            .sr(N__24783));
    defparam \nx.bit_ctr__i23_LC_4_29_7 .C_ON=1'b1;
    defparam \nx.bit_ctr__i23_LC_4_29_7 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i23_LC_4_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i23_LC_4_29_7  (
            .in0(_gnd_net_),
            .in1(N__24534),
            .in2(_gnd_net_),
            .in3(N__24465),
            .lcout(\nx.bit_ctr_23 ),
            .ltout(),
            .carryin(\nx.n10413 ),
            .carryout(\nx.n10414 ),
            .clk(N__48432),
            .ce(N__24846),
            .sr(N__24783));
    defparam \nx.bit_ctr__i24_LC_4_30_0 .C_ON=1'b1;
    defparam \nx.bit_ctr__i24_LC_4_30_0 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i24_LC_4_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i24_LC_4_30_0  (
            .in0(_gnd_net_),
            .in1(N__24444),
            .in2(_gnd_net_),
            .in3(N__24423),
            .lcout(\nx.bit_ctr_24 ),
            .ltout(),
            .carryin(bfn_4_30_0_),
            .carryout(\nx.n10415 ),
            .clk(N__48437),
            .ce(N__24845),
            .sr(N__24779));
    defparam \nx.bit_ctr__i25_LC_4_30_1 .C_ON=1'b1;
    defparam \nx.bit_ctr__i25_LC_4_30_1 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i25_LC_4_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i25_LC_4_30_1  (
            .in0(_gnd_net_),
            .in1(N__26219),
            .in2(_gnd_net_),
            .in3(N__24420),
            .lcout(\nx.bit_ctr_25 ),
            .ltout(),
            .carryin(\nx.n10415 ),
            .carryout(\nx.n10416 ),
            .clk(N__48437),
            .ce(N__24845),
            .sr(N__24779));
    defparam \nx.bit_ctr__i26_LC_4_30_2 .C_ON=1'b1;
    defparam \nx.bit_ctr__i26_LC_4_30_2 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i26_LC_4_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i26_LC_4_30_2  (
            .in0(_gnd_net_),
            .in1(N__28056),
            .in2(_gnd_net_),
            .in3(N__24417),
            .lcout(\nx.bit_ctr_26 ),
            .ltout(),
            .carryin(\nx.n10416 ),
            .carryout(\nx.n10417 ),
            .clk(N__48437),
            .ce(N__24845),
            .sr(N__24779));
    defparam \nx.bit_ctr__i27_LC_4_30_3 .C_ON=1'b1;
    defparam \nx.bit_ctr__i27_LC_4_30_3 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i27_LC_4_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i27_LC_4_30_3  (
            .in0(_gnd_net_),
            .in1(N__27732),
            .in2(_gnd_net_),
            .in3(N__24414),
            .lcout(\nx.bit_ctr_27 ),
            .ltout(),
            .carryin(\nx.n10417 ),
            .carryout(\nx.n10418 ),
            .clk(N__48437),
            .ce(N__24845),
            .sr(N__24779));
    defparam \nx.bit_ctr__i28_LC_4_30_4 .C_ON=1'b1;
    defparam \nx.bit_ctr__i28_LC_4_30_4 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i28_LC_4_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i28_LC_4_30_4  (
            .in0(_gnd_net_),
            .in1(N__27678),
            .in2(_gnd_net_),
            .in3(N__24411),
            .lcout(\nx.bit_ctr_28 ),
            .ltout(),
            .carryin(\nx.n10418 ),
            .carryout(\nx.n10419 ),
            .clk(N__48437),
            .ce(N__24845),
            .sr(N__24779));
    defparam \nx.bit_ctr__i29_LC_4_30_5 .C_ON=1'b1;
    defparam \nx.bit_ctr__i29_LC_4_30_5 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i29_LC_4_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i29_LC_4_30_5  (
            .in0(_gnd_net_),
            .in1(N__26504),
            .in2(_gnd_net_),
            .in3(N__24408),
            .lcout(\nx.bit_ctr_29 ),
            .ltout(),
            .carryin(\nx.n10419 ),
            .carryout(\nx.n10420 ),
            .clk(N__48437),
            .ce(N__24845),
            .sr(N__24779));
    defparam \nx.bit_ctr__i30_LC_4_30_6 .C_ON=1'b1;
    defparam \nx.bit_ctr__i30_LC_4_30_6 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i30_LC_4_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i30_LC_4_30_6  (
            .in0(_gnd_net_),
            .in1(N__26437),
            .in2(_gnd_net_),
            .in3(N__24405),
            .lcout(\nx.bit_ctr_30 ),
            .ltout(),
            .carryin(\nx.n10420 ),
            .carryout(\nx.n10421 ),
            .clk(N__48437),
            .ce(N__24845),
            .sr(N__24779));
    defparam \nx.bit_ctr__i31_LC_4_30_7 .C_ON=1'b0;
    defparam \nx.bit_ctr__i31_LC_4_30_7 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i31_LC_4_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i31_LC_4_30_7  (
            .in0(_gnd_net_),
            .in1(N__26557),
            .in2(_gnd_net_),
            .in3(N__24849),
            .lcout(\nx.bit_ctr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48437),
            .ce(N__24845),
            .sr(N__24779));
    defparam \nx.mod_5_i946_3_lut_LC_4_31_0 .C_ON=1'b0;
    defparam \nx.mod_5_i946_3_lut_LC_4_31_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i946_3_lut_LC_4_31_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i946_3_lut_LC_4_31_0  (
            .in0(_gnd_net_),
            .in1(N__24738),
            .in2(N__24708),
            .in3(N__24581),
            .lcout(\nx.n1407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i944_3_lut_LC_4_31_1 .C_ON=1'b0;
    defparam \nx.mod_5_i944_3_lut_LC_4_31_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i944_3_lut_LC_4_31_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i944_3_lut_LC_4_31_1  (
            .in0(_gnd_net_),
            .in1(N__24696),
            .in2(N__24591),
            .in3(N__24687),
            .lcout(\nx.n1405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i942_3_lut_LC_4_31_2 .C_ON=1'b0;
    defparam \nx.mod_5_i942_3_lut_LC_4_31_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i942_3_lut_LC_4_31_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i942_3_lut_LC_4_31_2  (
            .in0(_gnd_net_),
            .in1(N__24666),
            .in2(N__24657),
            .in3(N__24580),
            .lcout(\nx.n1403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i943_3_lut_LC_4_31_4 .C_ON=1'b0;
    defparam \nx.mod_5_i943_3_lut_LC_4_31_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i943_3_lut_LC_4_31_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i943_3_lut_LC_4_31_4  (
            .in0(_gnd_net_),
            .in1(N__24636),
            .in2(N__24603),
            .in3(N__24585),
            .lcout(\nx.n1404 ),
            .ltout(\nx.n1404_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_3_lut_adj_38_LC_4_31_5 .C_ON=1'b0;
    defparam \nx.i3_3_lut_adj_38_LC_4_31_5 .SEQ_MODE=4'b0000;
    defparam \nx.i3_3_lut_adj_38_LC_4_31_5 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i3_3_lut_adj_38_LC_4_31_5  (
            .in0(_gnd_net_),
            .in1(N__24971),
            .in2(N__24546),
            .in3(N__28243),
            .lcout(\nx.n13_adj_631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_137_LC_4_31_6 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_137_LC_4_31_6 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_137_LC_4_31_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_137_LC_4_31_6  (
            .in0(N__34074),
            .in1(N__24541),
            .in2(N__26505),
            .in3(N__43548),
            .lcout(\nx.n47_adj_706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1010_3_lut_LC_4_32_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1010_3_lut_LC_4_32_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1010_3_lut_LC_4_32_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1010_3_lut_LC_4_32_1  (
            .in0(_gnd_net_),
            .in1(N__24488),
            .in2(N__28202),
            .in3(N__24474),
            .lcout(\nx.n1503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1016_3_lut_LC_4_32_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1016_3_lut_LC_4_32_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1016_3_lut_LC_4_32_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i1016_3_lut_LC_4_32_2  (
            .in0(N__24975),
            .in1(N__24939),
            .in2(_gnd_net_),
            .in3(N__28182),
            .lcout(\nx.n1509 ),
            .ltout(\nx.n1509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6448_2_lut_LC_4_32_3 .C_ON=1'b0;
    defparam \nx.i6448_2_lut_LC_4_32_3 .SEQ_MODE=4'b0000;
    defparam \nx.i6448_2_lut_LC_4_32_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \nx.i6448_2_lut_LC_4_32_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24933),
            .in3(N__30837),
            .lcout(\nx.n9672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8_3_lut_LC_4_32_4 .C_ON=1'b0;
    defparam \nx.i8_3_lut_LC_4_32_4 .SEQ_MODE=4'b0000;
    defparam \nx.i8_3_lut_LC_4_32_4 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \nx.i8_3_lut_LC_4_32_4  (
            .in0(_gnd_net_),
            .in1(N__26792),
            .in2(N__26684),
            .in3(N__24930),
            .lcout(),
            .ltout(\nx.n18_adj_630_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_LC_4_32_5 .C_ON=1'b0;
    defparam \nx.i9_4_lut_LC_4_32_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_LC_4_32_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_LC_4_32_5  (
            .in0(N__26719),
            .in1(N__26848),
            .in2(N__24924),
            .in3(N__24921),
            .lcout(\nx.n1433 ),
            .ltout(\nx.n1433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1008_3_lut_LC_4_32_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1008_3_lut_LC_4_32_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1008_3_lut_LC_4_32_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1008_3_lut_LC_4_32_6  (
            .in0(_gnd_net_),
            .in1(N__24915),
            .in2(N__24906),
            .in3(N__24902),
            .lcout(\nx.n1501 ),
            .ltout(\nx.n1501_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_4_lut_adj_39_LC_4_32_7 .C_ON=1'b0;
    defparam \nx.i7_4_lut_adj_39_LC_4_32_7 .SEQ_MODE=4'b0000;
    defparam \nx.i7_4_lut_adj_39_LC_4_32_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i7_4_lut_adj_39_LC_4_32_7  (
            .in0(N__28351),
            .in1(N__31016),
            .in2(N__24885),
            .in3(N__24882),
            .lcout(\nx.n18_adj_632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i22_LC_5_16_2 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i22_LC_5_16_2 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i22_LC_5_16_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i22_LC_5_16_2  (
            .in0(N__24876),
            .in1(N__29276),
            .in2(_gnd_net_),
            .in3(N__28865),
            .lcout(neo_pixel_transmitter_t0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48405),
            .ce(),
            .sr(_gnd_net_));
    defparam i9323_3_lut_LC_5_17_0.C_ON=1'b0;
    defparam i9323_3_lut_LC_5_17_0.SEQ_MODE=4'b0000;
    defparam i9323_3_lut_LC_5_17_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i9323_3_lut_LC_5_17_0 (
            .in0(N__49091),
            .in1(N__47015),
            .in2(_gnd_net_),
            .in3(N__48993),
            .lcout(n13170),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9324_3_lut_LC_5_17_2.C_ON=1'b0;
    defparam i9324_3_lut_LC_5_17_2.SEQ_MODE=4'b0000;
    defparam i9324_3_lut_LC_5_17_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 i9324_3_lut_LC_5_17_2 (
            .in0(N__39149),
            .in1(N__47084),
            .in2(_gnd_net_),
            .in3(N__48992),
            .lcout(n13171),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i19_LC_5_17_6 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i19_LC_5_17_6 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i19_LC_5_17_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i19_LC_5_17_6  (
            .in0(N__25128),
            .in1(N__28866),
            .in2(_gnd_net_),
            .in3(N__25059),
            .lcout(neo_pixel_transmitter_t0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48394),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_1__bdd_4_lut_9609_LC_5_18_1.C_ON=1'b0;
    defparam current_pin_1__bdd_4_lut_9609_LC_5_18_1.SEQ_MODE=4'b0000;
    defparam current_pin_1__bdd_4_lut_9609_LC_5_18_1.LUT_INIT=16'b1010111111000000;
    LogicCell40 current_pin_1__bdd_4_lut_9609_LC_5_18_1 (
            .in0(N__25101),
            .in1(N__25092),
            .in2(N__50574),
            .in3(N__50356),
            .lcout(n13450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i10_1_lut_LC_5_18_4 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i10_1_lut_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i10_1_lut_LC_5_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i10_1_lut_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25085),
            .lcout(\nx.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i20_1_lut_LC_5_18_7 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i20_1_lut_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i20_1_lut_LC_5_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i20_1_lut_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25058),
            .lcout(\nx.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i6_LC_5_19_0.C_ON=1'b0;
    defparam neopxl_color_prev_i6_LC_5_19_0.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i6_LC_5_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 neopxl_color_prev_i6_LC_5_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40758),
            .lcout(neopxl_color_prev_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48409),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_3_lut_adj_19_LC_5_19_1 .C_ON=1'b0;
    defparam \nx.i6_3_lut_adj_19_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.i6_3_lut_adj_19_LC_5_19_1 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i6_3_lut_adj_19_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__28543),
            .in2(N__29069),
            .in3(N__31454),
            .lcout(\nx.n29_adj_607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_5_19_2.C_ON=1'b0;
    defparam i3_4_lut_LC_5_19_2.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_5_19_2.LUT_INIT=16'b0110111111110110;
    LogicCell40 i3_4_lut_LC_5_19_2 (
            .in0(N__25029),
            .in1(N__40757),
            .in2(N__26652),
            .in3(N__25023),
            .lcout(n11_adj_775),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i13_LC_5_19_4.C_ON=1'b0;
    defparam neopxl_color_prev_i13_LC_5_19_4.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i13_LC_5_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 neopxl_color_prev_i13_LC_5_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28915),
            .lcout(neopxl_color_prev_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48409),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i21_1_lut_LC_5_19_5 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i21_1_lut_LC_5_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i21_1_lut_LC_5_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i21_1_lut_LC_5_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25148),
            .lcout(\nx.n13_adj_649 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1896_3_lut_LC_5_19_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1896_3_lut_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1896_3_lut_LC_5_19_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1896_3_lut_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(N__29033),
            .in2(N__29013),
            .in3(N__36569),
            .lcout(\nx.n2805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i20_LC_5_19_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i20_LC_5_19_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i20_LC_5_19_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i20_LC_5_19_7  (
            .in0(N__25175),
            .in1(N__25149),
            .in2(_gnd_net_),
            .in3(N__28877),
            .lcout(neo_pixel_transmitter_t0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48409),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_26_LC_5_20_0 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_26_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_26_LC_5_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_26_LC_5_20_0  (
            .in0(N__27121),
            .in1(N__27271),
            .in2(N__26953),
            .in3(N__29668),
            .lcout(\nx.n39_adj_614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1891_rep_18_3_lut_LC_5_20_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1891_rep_18_3_lut_LC_5_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1891_rep_18_3_lut_LC_5_20_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1891_rep_18_3_lut_LC_5_20_1  (
            .in0(N__29244),
            .in1(_gnd_net_),
            .in2(N__36593),
            .in3(N__31599),
            .lcout(\nx.n2800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1900_3_lut_LC_5_20_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1900_3_lut_LC_5_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1900_3_lut_LC_5_20_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1900_3_lut_LC_5_20_2  (
            .in0(N__28491),
            .in1(N__28544),
            .in2(_gnd_net_),
            .in3(N__36565),
            .lcout(\nx.n2809 ),
            .ltout(\nx.n2809_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_3_lut_adj_25_LC_5_20_3 .C_ON=1'b0;
    defparam \nx.i7_3_lut_adj_25_LC_5_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.i7_3_lut_adj_25_LC_5_20_3 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \nx.i7_3_lut_adj_25_LC_5_20_3  (
            .in0(N__29826),
            .in1(_gnd_net_),
            .in2(N__25140),
            .in3(N__29890),
            .lcout(),
            .ltout(\nx.n31_adj_613_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_LC_5_20_4 .C_ON=1'b0;
    defparam \nx.i20_4_lut_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_LC_5_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i20_4_lut_LC_5_20_4  (
            .in0(N__26986),
            .in1(N__27163),
            .in2(N__25137),
            .in3(N__25134),
            .lcout(\nx.n44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1956_3_lut_LC_5_20_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1956_3_lut_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1956_3_lut_LC_5_20_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1956_3_lut_LC_5_20_5  (
            .in0(_gnd_net_),
            .in1(N__27094),
            .in2(N__30303),
            .in3(N__27072),
            .lcout(\nx.n2897 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1966_3_lut_LC_5_20_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1966_3_lut_LC_5_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1966_3_lut_LC_5_20_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1966_3_lut_LC_5_20_6  (
            .in0(N__26987),
            .in1(_gnd_net_),
            .in2(N__26970),
            .in3(N__30286),
            .lcout(\nx.n2907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1963_3_lut_LC_5_21_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1963_3_lut_LC_5_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1963_3_lut_LC_5_21_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1963_3_lut_LC_5_21_0  (
            .in0(_gnd_net_),
            .in1(N__26892),
            .in2(N__26919),
            .in3(N__30294),
            .lcout(\nx.n2904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1955_3_lut_LC_5_21_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1955_3_lut_LC_5_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1955_3_lut_LC_5_21_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1955_3_lut_LC_5_21_1  (
            .in0(_gnd_net_),
            .in1(N__27059),
            .in2(N__30305),
            .in3(N__27042),
            .lcout(\nx.n2896 ),
            .ltout(\nx.n2896_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_3_lut_adj_84_LC_5_21_2 .C_ON=1'b0;
    defparam \nx.i7_3_lut_adj_84_LC_5_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i7_3_lut_adj_84_LC_5_21_2 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i7_3_lut_adj_84_LC_5_21_2  (
            .in0(_gnd_net_),
            .in1(N__26135),
            .in2(N__25236),
            .in3(N__29777),
            .lcout(\nx.n32_adj_674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1965_3_lut_LC_5_21_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1965_3_lut_LC_5_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1965_3_lut_LC_5_21_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1965_3_lut_LC_5_21_3  (
            .in0(N__26931),
            .in1(_gnd_net_),
            .in2(N__30304),
            .in3(N__26957),
            .lcout(\nx.n2906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1960_3_lut_LC_5_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1960_3_lut_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1960_3_lut_LC_5_21_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1960_3_lut_LC_5_21_4  (
            .in0(_gnd_net_),
            .in1(N__27186),
            .in2(N__27216),
            .in3(N__30293),
            .lcout(\nx.n2901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1957_3_lut_LC_5_21_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1957_3_lut_LC_5_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1957_3_lut_LC_5_21_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1957_3_lut_LC_5_21_5  (
            .in0(_gnd_net_),
            .in1(N__27131),
            .in2(N__30306),
            .in3(N__27108),
            .lcout(\nx.n2898 ),
            .ltout(\nx.n2898_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_85_LC_5_21_6 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_85_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_85_LC_5_21_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_85_LC_5_21_6  (
            .in0(N__25342),
            .in1(N__25258),
            .in2(N__25233),
            .in3(N__25415),
            .lcout(),
            .ltout(\nx.n42_adj_675_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i21_4_lut_adj_88_LC_5_21_7 .C_ON=1'b0;
    defparam \nx.i21_4_lut_adj_88_LC_5_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.i21_4_lut_adj_88_LC_5_21_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i21_4_lut_adj_88_LC_5_21_7  (
            .in0(N__25559),
            .in1(N__29872),
            .in2(N__25230),
            .in3(N__25227),
            .lcout(\nx.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_2_lut_LC_5_22_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_2_lut_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_2_lut_LC_5_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_2_lut_LC_5_22_0  (
            .in0(_gnd_net_),
            .in1(N__26136),
            .in2(_gnd_net_),
            .in3(N__25200),
            .lcout(\nx.n2977 ),
            .ltout(),
            .carryin(bfn_5_22_0_),
            .carryout(\nx.n10837 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_3_lut_LC_5_22_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_3_lut_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_3_lut_LC_5_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_3_lut_LC_5_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29781),
            .in3(N__25182),
            .lcout(\nx.n2976 ),
            .ltout(),
            .carryin(\nx.n10837 ),
            .carryout(\nx.n10838 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_4_lut_LC_5_22_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_4_lut_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_4_lut_LC_5_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_4_lut_LC_5_22_2  (
            .in0(_gnd_net_),
            .in1(N__45557),
            .in2(N__25419),
            .in3(N__25386),
            .lcout(\nx.n2975 ),
            .ltout(),
            .carryin(\nx.n10838 ),
            .carryout(\nx.n10839 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_5_lut_LC_5_22_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_5_lut_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_5_lut_LC_5_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_5_lut_LC_5_22_3  (
            .in0(_gnd_net_),
            .in1(N__45563),
            .in2(N__25383),
            .in3(N__25350),
            .lcout(\nx.n2974 ),
            .ltout(),
            .carryin(\nx.n10839 ),
            .carryout(\nx.n10840 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_6_lut_LC_5_22_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_6_lut_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_6_lut_LC_5_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_6_lut_LC_5_22_4  (
            .in0(_gnd_net_),
            .in1(N__45558),
            .in2(N__25347),
            .in3(N__25320),
            .lcout(\nx.n2973 ),
            .ltout(),
            .carryin(\nx.n10840 ),
            .carryout(\nx.n10841 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_7_lut_LC_5_22_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_7_lut_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_7_lut_LC_5_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_7_lut_LC_5_22_5  (
            .in0(_gnd_net_),
            .in1(N__29443),
            .in2(N__45730),
            .in3(N__25308),
            .lcout(\nx.n2972 ),
            .ltout(),
            .carryin(\nx.n10841 ),
            .carryout(\nx.n10842 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_8_lut_LC_5_22_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_8_lut_LC_5_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_8_lut_LC_5_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_8_lut_LC_5_22_6  (
            .in0(_gnd_net_),
            .in1(N__45562),
            .in2(N__31913),
            .in3(N__25305),
            .lcout(\nx.n2971 ),
            .ltout(),
            .carryin(\nx.n10842 ),
            .carryout(\nx.n10843 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_9_lut_LC_5_22_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_9_lut_LC_5_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_9_lut_LC_5_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_9_lut_LC_5_22_7  (
            .in0(_gnd_net_),
            .in1(N__45564),
            .in2(N__30369),
            .in3(N__25290),
            .lcout(\nx.n2970 ),
            .ltout(),
            .carryin(\nx.n10843 ),
            .carryout(\nx.n10844 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_10_lut_LC_5_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_10_lut_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_10_lut_LC_5_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_10_lut_LC_5_23_0  (
            .in0(_gnd_net_),
            .in1(N__45551),
            .in2(N__30410),
            .in3(N__25272),
            .lcout(\nx.n2969 ),
            .ltout(),
            .carryin(bfn_5_23_0_),
            .carryout(\nx.n10845 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_11_lut_LC_5_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_11_lut_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_11_lut_LC_5_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_11_lut_LC_5_23_1  (
            .in0(_gnd_net_),
            .in1(N__45659),
            .in2(N__25269),
            .in3(N__25239),
            .lcout(\nx.n2968 ),
            .ltout(),
            .carryin(\nx.n10845 ),
            .carryout(\nx.n10846 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_12_lut_LC_5_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_12_lut_LC_5_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_12_lut_LC_5_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_12_lut_LC_5_23_2  (
            .in0(_gnd_net_),
            .in1(N__45552),
            .in2(N__29714),
            .in3(N__25566),
            .lcout(\nx.n2967 ),
            .ltout(),
            .carryin(\nx.n10846 ),
            .carryout(\nx.n10847 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_13_lut_LC_5_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_13_lut_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_13_lut_LC_5_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_13_lut_LC_5_23_3  (
            .in0(_gnd_net_),
            .in1(N__45660),
            .in2(N__25563),
            .in3(N__25542),
            .lcout(\nx.n2966 ),
            .ltout(),
            .carryin(\nx.n10847 ),
            .carryout(\nx.n10848 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_14_lut_LC_5_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_14_lut_LC_5_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_14_lut_LC_5_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_14_lut_LC_5_23_4  (
            .in0(_gnd_net_),
            .in1(N__45553),
            .in2(N__25539),
            .in3(N__25509),
            .lcout(\nx.n2965 ),
            .ltout(),
            .carryin(\nx.n10848 ),
            .carryout(\nx.n10849 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_15_lut_LC_5_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_15_lut_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_15_lut_LC_5_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_15_lut_LC_5_23_5  (
            .in0(_gnd_net_),
            .in1(N__45661),
            .in2(N__25505),
            .in3(N__25473),
            .lcout(\nx.n2964 ),
            .ltout(),
            .carryin(\nx.n10849 ),
            .carryout(\nx.n10850 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_16_lut_LC_5_23_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_16_lut_LC_5_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_16_lut_LC_5_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_16_lut_LC_5_23_6  (
            .in0(_gnd_net_),
            .in1(N__25469),
            .in2(N__45753),
            .in3(N__25443),
            .lcout(\nx.n2963 ),
            .ltout(),
            .carryin(\nx.n10850 ),
            .carryout(\nx.n10851 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_17_lut_LC_5_23_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_17_lut_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_17_lut_LC_5_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_17_lut_LC_5_23_7  (
            .in0(_gnd_net_),
            .in1(N__45665),
            .in2(N__29873),
            .in3(N__25434),
            .lcout(\nx.n2962 ),
            .ltout(),
            .carryin(\nx.n10851 ),
            .carryout(\nx.n10852 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_18_lut_LC_5_24_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_18_lut_LC_5_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_18_lut_LC_5_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_18_lut_LC_5_24_0  (
            .in0(_gnd_net_),
            .in1(N__45540),
            .in2(N__25869),
            .in3(N__25431),
            .lcout(\nx.n2961 ),
            .ltout(),
            .carryin(bfn_5_24_0_),
            .carryout(\nx.n10853 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_19_lut_LC_5_24_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_19_lut_LC_5_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_19_lut_LC_5_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_19_lut_LC_5_24_1  (
            .in0(_gnd_net_),
            .in1(N__45565),
            .in2(N__29651),
            .in3(N__25422),
            .lcout(\nx.n2960 ),
            .ltout(),
            .carryin(\nx.n10853 ),
            .carryout(\nx.n10854 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_20_lut_LC_5_24_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_20_lut_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_20_lut_LC_5_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_20_lut_LC_5_24_2  (
            .in0(_gnd_net_),
            .in1(N__45541),
            .in2(N__29529),
            .in3(N__25674),
            .lcout(\nx.n2959 ),
            .ltout(),
            .carryin(\nx.n10854 ),
            .carryout(\nx.n10855 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_21_lut_LC_5_24_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_21_lut_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_21_lut_LC_5_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_21_lut_LC_5_24_3  (
            .in0(_gnd_net_),
            .in1(N__45566),
            .in2(N__27541),
            .in3(N__25662),
            .lcout(\nx.n2958 ),
            .ltout(),
            .carryin(\nx.n10855 ),
            .carryout(\nx.n10856 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_22_lut_LC_5_24_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_22_lut_LC_5_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_22_lut_LC_5_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_22_lut_LC_5_24_4  (
            .in0(_gnd_net_),
            .in1(N__45542),
            .in2(N__29570),
            .in3(N__25653),
            .lcout(\nx.n2957 ),
            .ltout(),
            .carryin(\nx.n10856 ),
            .carryout(\nx.n10857 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_23_lut_LC_5_24_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_23_lut_LC_5_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_23_lut_LC_5_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_23_lut_LC_5_24_5  (
            .in0(_gnd_net_),
            .in1(N__45567),
            .in2(N__30143),
            .in3(N__25644),
            .lcout(\nx.n2956 ),
            .ltout(),
            .carryin(\nx.n10857 ),
            .carryout(\nx.n10858 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_24_lut_LC_5_24_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_24_lut_LC_5_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_24_lut_LC_5_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_24_lut_LC_5_24_6  (
            .in0(_gnd_net_),
            .in1(N__45543),
            .in2(N__30488),
            .in3(N__25635),
            .lcout(\nx.n2955 ),
            .ltout(),
            .carryin(\nx.n10858 ),
            .carryout(\nx.n10859 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_25_lut_LC_5_24_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_25_lut_LC_5_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_25_lut_LC_5_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_25_lut_LC_5_24_7  (
            .in0(_gnd_net_),
            .in1(N__29585),
            .in2(N__45729),
            .in3(N__25623),
            .lcout(\nx.n2954 ),
            .ltout(),
            .carryin(\nx.n10859 ),
            .carryout(\nx.n10860 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_26_lut_LC_5_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_26_lut_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_26_lut_LC_5_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_26_lut_LC_5_25_0  (
            .in0(_gnd_net_),
            .in1(N__29966),
            .in2(N__45727),
            .in3(N__25611),
            .lcout(\nx.n2953 ),
            .ltout(),
            .carryin(bfn_5_25_0_),
            .carryout(\nx.n10861 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_27_lut_LC_5_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_add_2009_27_lut_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_27_lut_LC_5_25_1 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_2009_27_lut_LC_5_25_1  (
            .in0(N__45526),
            .in1(N__31867),
            .in2(N__27578),
            .in3(N__25608),
            .lcout(\nx.n2984 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2020_3_lut_LC_5_25_2 .C_ON=1'b0;
    defparam \nx.mod_5_i2020_3_lut_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2020_3_lut_LC_5_25_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i2020_3_lut_LC_5_25_2  (
            .in0(N__25584),
            .in1(_gnd_net_),
            .in2(N__31877),
            .in3(N__25868),
            .lcout(\nx.n2993 ),
            .ltout(\nx.n2993_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2087_3_lut_LC_5_25_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2087_3_lut_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2087_3_lut_LC_5_25_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2087_3_lut_LC_5_25_3  (
            .in0(_gnd_net_),
            .in1(N__25827),
            .in2(N__25815),
            .in3(N__27458),
            .lcout(\nx.n3092 ),
            .ltout(\nx.n3092_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i23_4_lut_adj_106_LC_5_25_4 .C_ON=1'b0;
    defparam \nx.i23_4_lut_adj_106_LC_5_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.i23_4_lut_adj_106_LC_5_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i23_4_lut_adj_106_LC_5_25_4  (
            .in0(N__25793),
            .in1(N__25713),
            .in2(N__25764),
            .in3(N__25761),
            .lcout(\nx.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_2_lut_LC_5_25_7 .C_ON=1'b0;
    defparam \nx.i9_2_lut_LC_5_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.i9_2_lut_LC_5_25_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i9_2_lut_LC_5_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27307),
            .in3(N__25729),
            .lcout(\nx.n36_adj_687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_2_lut_LC_5_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_2_lut_LC_5_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_2_lut_LC_5_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_2_lut_LC_5_26_0  (
            .in0(_gnd_net_),
            .in1(N__26230),
            .in2(_gnd_net_),
            .in3(N__25695),
            .lcout(\nx.n1077 ),
            .ltout(),
            .carryin(bfn_5_26_0_),
            .carryout(\nx.n10468 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_3_lut_LC_5_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_3_lut_LC_5_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_3_lut_LC_5_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_3_lut_LC_5_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26253),
            .in3(N__25692),
            .lcout(\nx.n1076 ),
            .ltout(),
            .carryin(\nx.n10468 ),
            .carryout(\nx.n10469 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_4_lut_LC_5_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_4_lut_LC_5_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_4_lut_LC_5_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_4_lut_LC_5_26_2  (
            .in0(_gnd_net_),
            .in1(N__26391),
            .in2(N__45704),
            .in3(N__25689),
            .lcout(\nx.n1075 ),
            .ltout(),
            .carryin(\nx.n10469 ),
            .carryout(\nx.n10470 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_5_lut_LC_5_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_5_lut_LC_5_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_5_lut_LC_5_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_5_lut_LC_5_26_3  (
            .in0(_gnd_net_),
            .in1(N__45501),
            .in2(N__26316),
            .in3(N__25686),
            .lcout(\nx.n1074 ),
            .ltout(),
            .carryin(\nx.n10470 ),
            .carryout(\nx.n10471 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_6_lut_LC_5_26_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_6_lut_LC_5_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_6_lut_LC_5_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_6_lut_LC_5_26_4  (
            .in0(_gnd_net_),
            .in1(N__45525),
            .in2(N__27767),
            .in3(N__25683),
            .lcout(\nx.n1073 ),
            .ltout(),
            .carryin(\nx.n10471 ),
            .carryout(\nx.n10472 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_7_lut_LC_5_26_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_7_lut_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_7_lut_LC_5_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_7_lut_LC_5_26_5  (
            .in0(_gnd_net_),
            .in1(N__45502),
            .in2(N__26082),
            .in3(N__25983),
            .lcout(\nx.n1072 ),
            .ltout(),
            .carryin(\nx.n10472 ),
            .carryout(\nx.n10473 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_8_lut_LC_5_26_6 .C_ON=1'b0;
    defparam \nx.mod_5_add_736_8_lut_LC_5_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_8_lut_LC_5_26_6 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_736_8_lut_LC_5_26_6  (
            .in0(N__45503),
            .in1(N__26048),
            .in2(N__27891),
            .in3(N__25980),
            .lcout(\nx.n1103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_2_lut_LC_5_26_7 .C_ON=1'b0;
    defparam \nx.mod_5_add_1272_2_lut_LC_5_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_2_lut_LC_5_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_2_lut_LC_5_26_7  (
            .in0(_gnd_net_),
            .in1(N__45497),
            .in2(_gnd_net_),
            .in3(N__32763),
            .lcout(\nx.n1877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_136_LC_5_27_0 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_136_LC_5_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_136_LC_5_27_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_136_LC_5_27_0  (
            .in0(N__35880),
            .in1(N__27737),
            .in2(N__26235),
            .in3(N__37881),
            .lcout(\nx.n46_adj_705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i742_3_lut_LC_5_27_1 .C_ON=1'b0;
    defparam \nx.mod_5_i742_3_lut_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i742_3_lut_LC_5_27_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i742_3_lut_LC_5_27_1  (
            .in0(N__25941),
            .in1(N__26390),
            .in2(_gnd_net_),
            .in3(N__26046),
            .lcout(\nx.n1107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9571_2_lut_LC_5_27_2 .C_ON=1'b0;
    defparam \nx.i9571_2_lut_LC_5_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9571_2_lut_LC_5_27_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \nx.i9571_2_lut_LC_5_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27972),
            .in3(N__30639),
            .lcout(\nx.n1007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i740_3_lut_LC_5_27_3 .C_ON=1'b0;
    defparam \nx.mod_5_i740_3_lut_LC_5_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i740_3_lut_LC_5_27_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i740_3_lut_LC_5_27_3  (
            .in0(_gnd_net_),
            .in1(N__25902),
            .in2(N__27768),
            .in3(N__26047),
            .lcout(\nx.n1105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1219_3_lut_LC_5_27_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1219_3_lut_LC_5_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1219_3_lut_LC_5_27_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1219_3_lut_LC_5_27_4  (
            .in0(_gnd_net_),
            .in1(N__34887),
            .in2(N__34916),
            .in3(N__35148),
            .lcout(\nx.n1808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7853_3_lut_LC_5_27_5 .C_ON=1'b0;
    defparam \nx.i7853_3_lut_LC_5_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.i7853_3_lut_LC_5_27_5 .LUT_INIT=16'b1111000011110011;
    LogicCell40 \nx.i7853_3_lut_LC_5_27_5  (
            .in0(_gnd_net_),
            .in1(N__27956),
            .in2(N__30645),
            .in3(N__27971),
            .lcout(),
            .ltout(\nx.n11617_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_4_lut_LC_5_27_6 .C_ON=1'b0;
    defparam \nx.i4_4_lut_LC_5_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.i4_4_lut_LC_5_27_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \nx.i4_4_lut_LC_5_27_6  (
            .in0(N__26389),
            .in1(N__26181),
            .in2(N__26364),
            .in3(N__27884),
            .lcout(\nx.n1037 ),
            .ltout(\nx.n1037_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i743_3_lut_LC_5_27_7 .C_ON=1'b0;
    defparam \nx.mod_5_i743_3_lut_LC_5_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i743_3_lut_LC_5_27_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i743_3_lut_LC_5_27_7  (
            .in0(_gnd_net_),
            .in1(N__26361),
            .in2(N__26355),
            .in3(N__26249),
            .lcout(\nx.n1108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i741_3_lut_LC_5_28_0 .C_ON=1'b0;
    defparam \nx.mod_5_i741_3_lut_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i741_3_lut_LC_5_28_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i741_3_lut_LC_5_28_0  (
            .in0(N__26315),
            .in1(N__26301),
            .in2(_gnd_net_),
            .in3(N__26044),
            .lcout(\nx.n1106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i676_3_lut_LC_5_28_2 .C_ON=1'b0;
    defparam \nx.mod_5_i676_3_lut_LC_5_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i676_3_lut_LC_5_28_2 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \nx.mod_5_i676_3_lut_LC_5_28_2  (
            .in0(N__30625),
            .in1(N__28023),
            .in2(N__28070),
            .in3(_gnd_net_),
            .lcout(\nx.n1009 ),
            .ltout(\nx.n1009_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2_3_lut_LC_5_28_3 .C_ON=1'b0;
    defparam \nx.i2_3_lut_LC_5_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.i2_3_lut_LC_5_28_3 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \nx.i2_3_lut_LC_5_28_3  (
            .in0(_gnd_net_),
            .in1(N__26223),
            .in2(N__26184),
            .in3(N__26075),
            .lcout(\nx.n7_adj_616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_139_LC_5_28_4 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_139_LC_5_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_139_LC_5_28_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_139_LC_5_28_4  (
            .in0(N__27689),
            .in1(N__26169),
            .in2(N__41268),
            .in3(N__26118),
            .lcout(\nx.n44_adj_708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i672_3_lut_LC_5_28_5 .C_ON=1'b0;
    defparam \nx.mod_5_i672_3_lut_LC_5_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i672_3_lut_LC_5_28_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \nx.mod_5_i672_3_lut_LC_5_28_5  (
            .in0(_gnd_net_),
            .in1(N__30627),
            .in2(N__27939),
            .in3(N__27915),
            .lcout(\nx.n1005 ),
            .ltout(\nx.n1005_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i739_3_lut_LC_5_28_6 .C_ON=1'b0;
    defparam \nx.mod_5_i739_3_lut_LC_5_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i739_3_lut_LC_5_28_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i739_3_lut_LC_5_28_6  (
            .in0(_gnd_net_),
            .in1(N__26064),
            .in2(N__26055),
            .in3(N__26045),
            .lcout(\nx.n1104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i675_3_lut_LC_5_28_7 .C_ON=1'b0;
    defparam \nx.mod_5_i675_3_lut_LC_5_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i675_3_lut_LC_5_28_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i675_3_lut_LC_5_28_7  (
            .in0(_gnd_net_),
            .in1(N__28013),
            .in2(N__27999),
            .in3(N__30626),
            .lcout(\nx.n1008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_158_LC_5_29_0 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_158_LC_5_29_0 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_158_LC_5_29_0 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \nx.i1_2_lut_adj_158_LC_5_29_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27736),
            .in3(N__27816),
            .lcout(\nx.n7082 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9585_4_lut_LC_5_29_1 .C_ON=1'b0;
    defparam \nx.i9585_4_lut_LC_5_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9585_4_lut_LC_5_29_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \nx.i9585_4_lut_LC_5_29_1  (
            .in0(N__27873),
            .in1(N__27853),
            .in2(N__27825),
            .in3(N__26573),
            .lcout(\nx.n13064 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9228_4_lut_LC_5_29_2 .C_ON=1'b0;
    defparam \nx.i9228_4_lut_LC_5_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9228_4_lut_LC_5_29_2 .LUT_INIT=16'b1100001101101001;
    LogicCell40 \nx.i9228_4_lut_LC_5_29_2  (
            .in0(N__27724),
            .in1(N__27674),
            .in2(N__27636),
            .in3(N__27815),
            .lcout(\nx.n7342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_29_LC_5_29_3 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_29_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_29_LC_5_29_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \nx.i1_2_lut_adj_29_LC_5_29_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27682),
            .in3(N__27631),
            .lcout(),
            .ltout(\nx.n7084_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_27_LC_5_29_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_27_LC_5_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_27_LC_5_29_4 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \nx.i1_4_lut_adj_27_LC_5_29_4  (
            .in0(N__27723),
            .in1(N__26572),
            .in2(N__26373),
            .in3(N__27841),
            .lcout(\nx.n838 ),
            .ltout(\nx.n838_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_3_lut_4_lut_adj_143_LC_5_29_5 .C_ON=1'b0;
    defparam \nx.i1_3_lut_4_lut_adj_143_LC_5_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.i1_3_lut_4_lut_adj_143_LC_5_29_5 .LUT_INIT=16'b0000000001111011;
    LogicCell40 \nx.i1_3_lut_4_lut_adj_143_LC_5_29_5  (
            .in0(N__27728),
            .in1(N__28052),
            .in2(N__26370),
            .in3(N__27983),
            .lcout(),
            .ltout(\nx.n12595_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_28_LC_5_29_6 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_28_LC_5_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_28_LC_5_29_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \nx.i1_4_lut_adj_28_LC_5_29_6  (
            .in0(N__27794),
            .in1(N__27905),
            .in2(N__26367),
            .in3(N__27931),
            .lcout(\nx.n10994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i605_4_lut_LC_5_29_7 .C_ON=1'b0;
    defparam \nx.mod_5_i605_4_lut_LC_5_29_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i605_4_lut_LC_5_29_7 .LUT_INIT=16'b1111111000000001;
    LogicCell40 \nx.mod_5_i605_4_lut_LC_5_29_7  (
            .in0(N__27872),
            .in1(N__27854),
            .in2(N__27824),
            .in3(N__26574),
            .lcout(\nx.n906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6377_2_lut_LC_5_30_0 .C_ON=1'b0;
    defparam \nx.i6377_2_lut_LC_5_30_0 .SEQ_MODE=4'b0000;
    defparam \nx.i6377_2_lut_LC_5_30_0 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \nx.i6377_2_lut_LC_5_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26558),
            .in3(N__26428),
            .lcout(\nx.n608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_3_lut_LC_5_30_1 .C_ON=1'b0;
    defparam \nx.i1_3_lut_LC_5_30_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_3_lut_LC_5_30_1 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \nx.i1_3_lut_LC_5_30_1  (
            .in0(_gnd_net_),
            .in1(N__26548),
            .in2(N__26438),
            .in3(N__26497),
            .lcout(\nx.n9618 ),
            .ltout(\nx.n9618_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9471_4_lut_4_lut_LC_5_30_2 .C_ON=1'b0;
    defparam \nx.i9471_4_lut_4_lut_LC_5_30_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9471_4_lut_4_lut_LC_5_30_2 .LUT_INIT=16'b1010001001101100;
    LogicCell40 \nx.i9471_4_lut_4_lut_LC_5_30_2  (
            .in0(N__26498),
            .in1(N__26432),
            .in2(N__26613),
            .in3(N__26552),
            .lcout(\nx.n708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7854_rep_2_3_lut_4_lut_LC_5_30_3 .C_ON=1'b0;
    defparam \nx.i7854_rep_2_3_lut_4_lut_LC_5_30_3 .SEQ_MODE=4'b0000;
    defparam \nx.i7854_rep_2_3_lut_4_lut_LC_5_30_3 .LUT_INIT=16'b0010001000101000;
    LogicCell40 \nx.i7854_rep_2_3_lut_4_lut_LC_5_30_3  (
            .in0(N__27666),
            .in1(N__26499),
            .in2(N__26610),
            .in3(N__26518),
            .lcout(\nx.n11738 ),
            .ltout(\nx.n11738_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_LC_5_30_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_LC_5_30_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_LC_5_30_4 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \nx.i1_4_lut_LC_5_30_4  (
            .in0(N__26609),
            .in1(N__26522),
            .in2(N__26595),
            .in3(N__26591),
            .lcout(\nx.n739 ),
            .ltout(\nx.n739_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i538_3_lut_LC_5_30_5 .C_ON=1'b0;
    defparam \nx.mod_5_i538_3_lut_LC_5_30_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i538_3_lut_LC_5_30_5 .LUT_INIT=16'b1010101010100101;
    LogicCell40 \nx.mod_5_i538_3_lut_LC_5_30_5  (
            .in0(N__26592),
            .in1(_gnd_net_),
            .in2(N__26583),
            .in3(N__26580),
            .lcout(\nx.n807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6508_rep_3_2_lut_3_lut_LC_5_30_6 .C_ON=1'b0;
    defparam \nx.i6508_rep_3_2_lut_3_lut_LC_5_30_6 .SEQ_MODE=4'b0000;
    defparam \nx.i6508_rep_3_2_lut_3_lut_LC_5_30_6 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \nx.i6508_rep_3_2_lut_3_lut_LC_5_30_6  (
            .in0(_gnd_net_),
            .in1(N__26553),
            .in2(N__26523),
            .in3(N__26433),
            .lcout(),
            .ltout(\nx.n11771_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9479_4_lut_LC_5_30_7 .C_ON=1'b0;
    defparam \nx.i9479_4_lut_LC_5_30_7 .SEQ_MODE=4'b0000;
    defparam \nx.i9479_4_lut_LC_5_30_7 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \nx.i9479_4_lut_LC_5_30_7  (
            .in0(N__27667),
            .in1(N__26500),
            .in2(N__26475),
            .in3(N__27627),
            .lcout(\nx.n11559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1009_3_lut_LC_5_31_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1009_3_lut_LC_5_31_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1009_3_lut_LC_5_31_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1009_3_lut_LC_5_31_0  (
            .in0(_gnd_net_),
            .in1(N__26472),
            .in2(N__26463),
            .in3(N__28186),
            .lcout(\nx.n1502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_adj_135_LC_5_31_1 .C_ON=1'b0;
    defparam \nx.i20_4_lut_adj_135_LC_5_31_1 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_adj_135_LC_5_31_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i20_4_lut_adj_135_LC_5_31_1  (
            .in0(N__29827),
            .in1(N__30846),
            .in2(N__30115),
            .in3(N__26439),
            .lcout(\nx.n48_adj_704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1013_3_lut_LC_5_31_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1013_3_lut_LC_5_31_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1013_3_lut_LC_5_31_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1013_3_lut_LC_5_31_2  (
            .in0(_gnd_net_),
            .in1(N__26849),
            .in2(N__26829),
            .in3(N__28188),
            .lcout(\nx.n1506 ),
            .ltout(\nx.n1506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_40_LC_5_31_3 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_40_LC_5_31_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_40_LC_5_31_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_adj_40_LC_5_31_3  (
            .in0(N__28279),
            .in1(N__28937),
            .in2(N__26817),
            .in3(N__26814),
            .lcout(\nx.n20_adj_634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1014_3_lut_LC_5_31_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1014_3_lut_LC_5_31_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1014_3_lut_LC_5_31_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1014_3_lut_LC_5_31_4  (
            .in0(_gnd_net_),
            .in1(N__26808),
            .in2(N__26799),
            .in3(N__28187),
            .lcout(\nx.n1507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1007_3_lut_LC_5_32_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1007_3_lut_LC_5_32_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1007_3_lut_LC_5_32_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1007_3_lut_LC_5_32_4  (
            .in0(_gnd_net_),
            .in1(N__26766),
            .in2(N__28207),
            .in3(N__26742),
            .lcout(\nx.n1500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1011_3_lut_LC_5_32_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1011_3_lut_LC_5_32_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1011_3_lut_LC_5_32_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1011_3_lut_LC_5_32_6  (
            .in0(N__26733),
            .in1(_gnd_net_),
            .in2(N__28208),
            .in3(N__26720),
            .lcout(\nx.n1504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1012_3_lut_LC_5_32_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1012_3_lut_LC_5_32_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1012_3_lut_LC_5_32_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1012_3_lut_LC_5_32_7  (
            .in0(_gnd_net_),
            .in1(N__26700),
            .in2(N__26688),
            .in3(N__28195),
            .lcout(\nx.n1505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i15_LC_6_16_1.C_ON=1'b0;
    defparam neopxl_color_i15_LC_6_16_1.SEQ_MODE=4'b1000;
    defparam neopxl_color_i15_LC_6_16_1.LUT_INIT=16'b1111011100010000;
    LogicCell40 neopxl_color_i15_LC_6_16_1 (
            .in0(N__50075),
            .in1(N__49843),
            .in2(N__49600),
            .in3(N__26646),
            .lcout(neopxl_color_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48410),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1830_3_lut_LC_6_18_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1830_3_lut_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1830_3_lut_LC_6_18_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1830_3_lut_LC_6_18_0  (
            .in0(_gnd_net_),
            .in1(N__35826),
            .in2(N__36209),
            .in3(N__33441),
            .lcout(\nx.n2707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1823_3_lut_LC_6_18_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1823_3_lut_LC_6_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1823_3_lut_LC_6_18_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1823_3_lut_LC_6_18_1  (
            .in0(_gnd_net_),
            .in1(N__37668),
            .in2(N__33588),
            .in3(N__36206),
            .lcout(\nx.n2700 ),
            .ltout(\nx.n2700_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_21_LC_6_18_2 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_21_LC_6_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_21_LC_6_18_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_21_LC_6_18_2  (
            .in0(N__28969),
            .in1(N__29032),
            .in2(N__26856),
            .in3(N__29101),
            .lcout(\nx.n40_adj_609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1831_3_lut_LC_6_18_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1831_3_lut_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1831_3_lut_LC_6_18_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1831_3_lut_LC_6_18_3  (
            .in0(_gnd_net_),
            .in1(N__35928),
            .in2(N__33459),
            .in3(N__36199),
            .lcout(\nx.n2708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1829_3_lut_LC_6_18_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1829_3_lut_LC_6_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1829_3_lut_LC_6_18_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1829_3_lut_LC_6_18_4  (
            .in0(_gnd_net_),
            .in1(N__33426),
            .in2(N__36210),
            .in3(N__39423),
            .lcout(\nx.n2706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1892_3_lut_LC_6_18_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1892_3_lut_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1892_3_lut_LC_6_18_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1892_3_lut_LC_6_18_6  (
            .in0(_gnd_net_),
            .in1(N__28953),
            .in2(N__28976),
            .in3(N__36575),
            .lcout(\nx.n2801 ),
            .ltout(\nx.n2801_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_42_LC_6_18_7 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_42_LC_6_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_42_LC_6_18_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_42_LC_6_18_7  (
            .in0(N__27202),
            .in1(N__26911),
            .in2(N__26853),
            .in3(N__27095),
            .lcout(\nx.n42_adj_635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1893_3_lut_LC_6_19_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1893_3_lut_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1893_3_lut_LC_6_19_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1893_3_lut_LC_6_19_0  (
            .in0(_gnd_net_),
            .in1(N__28986),
            .in2(N__36590),
            .in3(N__31482),
            .lcout(\nx.n2802 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1887_3_lut_LC_6_19_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1887_3_lut_LC_6_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1887_3_lut_LC_6_19_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1887_3_lut_LC_6_19_1  (
            .in0(_gnd_net_),
            .in1(N__31282),
            .in2(N__29184),
            .in3(N__36550),
            .lcout(\nx.n2796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1898_3_lut_LC_6_19_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1898_3_lut_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1898_3_lut_LC_6_19_2 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.mod_5_i1898_3_lut_LC_6_19_2  (
            .in0(N__36549),
            .in1(N__29082),
            .in2(N__29106),
            .in3(_gnd_net_),
            .lcout(\nx.n2807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1890_rep_19_3_lut_LC_6_19_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1890_rep_19_3_lut_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1890_rep_19_3_lut_LC_6_19_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1890_rep_19_3_lut_LC_6_19_3  (
            .in0(_gnd_net_),
            .in1(N__29211),
            .in2(N__29232),
            .in3(N__36548),
            .lcout(\nx.n2799 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_LC_6_19_4 .C_ON=1'b0;
    defparam \nx.i14_4_lut_LC_6_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_LC_6_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_LC_6_19_4  (
            .in0(N__31537),
            .in1(N__33853),
            .in2(N__31286),
            .in3(N__31312),
            .lcout(),
            .ltout(\nx.n37_adj_608_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_LC_6_19_5 .C_ON=1'b0;
    defparam \nx.i19_4_lut_LC_6_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_LC_6_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_LC_6_19_5  (
            .in0(N__26880),
            .in1(N__29167),
            .in2(N__26874),
            .in3(N__31564),
            .lcout(),
            .ltout(\nx.n42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i22_4_lut_LC_6_19_6 .C_ON=1'b0;
    defparam \nx.i22_4_lut_LC_6_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.i22_4_lut_LC_6_19_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i22_4_lut_LC_6_19_6  (
            .in0(N__31491),
            .in1(N__26871),
            .in2(N__26865),
            .in3(N__33978),
            .lcout(\nx.n2720 ),
            .ltout(\nx.n2720_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1885_3_lut_LC_6_19_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1885_3_lut_LC_6_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1885_3_lut_LC_6_19_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1885_3_lut_LC_6_19_7  (
            .in0(_gnd_net_),
            .in1(N__31538),
            .in2(N__26862),
            .in3(N__29130),
            .lcout(\nx.n2794 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1886_3_lut_LC_6_20_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1886_3_lut_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1886_3_lut_LC_6_20_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1886_3_lut_LC_6_20_0  (
            .in0(_gnd_net_),
            .in1(N__29171),
            .in2(N__29142),
            .in3(N__36554),
            .lcout(\nx.n2795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1879_3_lut_LC_6_20_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1879_3_lut_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1879_3_lut_LC_6_20_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1879_3_lut_LC_6_20_1  (
            .in0(N__31688),
            .in1(_gnd_net_),
            .in2(N__36591),
            .in3(N__29298),
            .lcout(\nx.n2788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1888_3_lut_LC_6_20_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1888_3_lut_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1888_3_lut_LC_6_20_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1888_3_lut_LC_6_20_2  (
            .in0(_gnd_net_),
            .in1(N__29193),
            .in2(N__31515),
            .in3(N__36564),
            .lcout(\nx.n2797 ),
            .ltout(\nx.n2797_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_49_LC_6_20_3 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_49_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_49_LC_6_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_49_LC_6_20_3  (
            .in0(N__36043),
            .in1(N__30442),
            .in2(N__26859),
            .in3(N__29470),
            .lcout(\nx.n41_adj_643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1889_3_lut_LC_6_20_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1889_3_lut_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1889_3_lut_LC_6_20_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1889_3_lut_LC_6_20_4  (
            .in0(_gnd_net_),
            .in1(N__29202),
            .in2(N__33813),
            .in3(N__36556),
            .lcout(\nx.n2798 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1897_rep_21_3_lut_LC_6_20_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1897_rep_21_3_lut_LC_6_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1897_rep_21_3_lut_LC_6_20_5 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.mod_5_i1897_rep_21_3_lut_LC_6_20_5  (
            .in0(N__36560),
            .in1(N__29043),
            .in2(N__29073),
            .in3(_gnd_net_),
            .lcout(\nx.n2806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1899_rep_16_3_lut_LC_6_20_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1899_rep_16_3_lut_LC_6_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1899_rep_16_3_lut_LC_6_20_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \nx.mod_5_i1899_rep_16_3_lut_LC_6_20_6  (
            .in0(_gnd_net_),
            .in1(N__36555),
            .in2(N__29118),
            .in3(N__31455),
            .lcout(\nx.n2808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1894_3_lut_LC_6_20_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1894_3_lut_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1894_3_lut_LC_6_20_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1894_3_lut_LC_6_20_7  (
            .in0(_gnd_net_),
            .in1(N__28995),
            .in2(N__36592),
            .in3(N__31569),
            .lcout(\nx.n2803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_2_lut_LC_6_21_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_2_lut_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_2_lut_LC_6_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_2_lut_LC_6_21_0  (
            .in0(_gnd_net_),
            .in1(N__29828),
            .in2(_gnd_net_),
            .in3(N__27030),
            .lcout(\nx.n2877 ),
            .ltout(),
            .carryin(bfn_6_21_0_),
            .carryout(\nx.n10813 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_3_lut_LC_6_21_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_3_lut_LC_6_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_3_lut_LC_6_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_3_lut_LC_6_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27020),
            .in3(N__26991),
            .lcout(\nx.n2876 ),
            .ltout(),
            .carryin(\nx.n10813 ),
            .carryout(\nx.n10814 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_4_lut_LC_6_21_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_4_lut_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_4_lut_LC_6_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_4_lut_LC_6_21_2  (
            .in0(_gnd_net_),
            .in1(N__45554),
            .in2(N__26988),
            .in3(N__26961),
            .lcout(\nx.n2875 ),
            .ltout(),
            .carryin(\nx.n10814 ),
            .carryout(\nx.n10815 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_5_lut_LC_6_21_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_5_lut_LC_6_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_5_lut_LC_6_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_5_lut_LC_6_21_3  (
            .in0(_gnd_net_),
            .in1(N__45656),
            .in2(N__26958),
            .in3(N__26925),
            .lcout(\nx.n2874 ),
            .ltout(),
            .carryin(\nx.n10815 ),
            .carryout(\nx.n10816 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_6_lut_LC_6_21_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_6_lut_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_6_lut_LC_6_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_6_lut_LC_6_21_4  (
            .in0(_gnd_net_),
            .in1(N__45555),
            .in2(N__29474),
            .in3(N__26922),
            .lcout(\nx.n2873 ),
            .ltout(),
            .carryin(\nx.n10816 ),
            .carryout(\nx.n10817 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_7_lut_LC_6_21_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_7_lut_LC_6_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_7_lut_LC_6_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_7_lut_LC_6_21_5  (
            .in0(_gnd_net_),
            .in1(N__45657),
            .in2(N__26918),
            .in3(N__26886),
            .lcout(\nx.n2872 ),
            .ltout(),
            .carryin(\nx.n10817 ),
            .carryout(\nx.n10818 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_8_lut_LC_6_21_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_8_lut_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_8_lut_LC_6_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_8_lut_LC_6_21_6  (
            .in0(_gnd_net_),
            .in1(N__45556),
            .in2(N__36047),
            .in3(N__26883),
            .lcout(\nx.n2871 ),
            .ltout(),
            .carryin(\nx.n10818 ),
            .carryout(\nx.n10819 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_9_lut_LC_6_21_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_9_lut_LC_6_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_9_lut_LC_6_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_9_lut_LC_6_21_7  (
            .in0(_gnd_net_),
            .in1(N__45658),
            .in2(N__30446),
            .in3(N__27219),
            .lcout(\nx.n2870 ),
            .ltout(),
            .carryin(\nx.n10819 ),
            .carryout(\nx.n10820 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_10_lut_LC_6_22_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_10_lut_LC_6_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_10_lut_LC_6_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_10_lut_LC_6_22_0  (
            .in0(_gnd_net_),
            .in1(N__45547),
            .in2(N__27215),
            .in3(N__27180),
            .lcout(\nx.n2869 ),
            .ltout(),
            .carryin(bfn_6_22_0_),
            .carryout(\nx.n10821 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_11_lut_LC_6_22_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_11_lut_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_11_lut_LC_6_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_11_lut_LC_6_22_1  (
            .in0(_gnd_net_),
            .in1(N__45645),
            .in2(N__29738),
            .in3(N__27177),
            .lcout(\nx.n2868 ),
            .ltout(),
            .carryin(\nx.n10821 ),
            .carryout(\nx.n10822 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_12_lut_LC_6_22_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_12_lut_LC_6_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_12_lut_LC_6_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_12_lut_LC_6_22_2  (
            .in0(_gnd_net_),
            .in1(N__45548),
            .in2(N__27174),
            .in3(N__27135),
            .lcout(\nx.n2867 ),
            .ltout(),
            .carryin(\nx.n10822 ),
            .carryout(\nx.n10823 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_13_lut_LC_6_22_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_13_lut_LC_6_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_13_lut_LC_6_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_13_lut_LC_6_22_3  (
            .in0(_gnd_net_),
            .in1(N__45646),
            .in2(N__27132),
            .in3(N__27102),
            .lcout(\nx.n2866 ),
            .ltout(),
            .carryin(\nx.n10823 ),
            .carryout(\nx.n10824 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_14_lut_LC_6_22_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_14_lut_LC_6_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_14_lut_LC_6_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_14_lut_LC_6_22_4  (
            .in0(_gnd_net_),
            .in1(N__45549),
            .in2(N__27099),
            .in3(N__27063),
            .lcout(\nx.n2865 ),
            .ltout(),
            .carryin(\nx.n10824 ),
            .carryout(\nx.n10825 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_15_lut_LC_6_22_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_15_lut_LC_6_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_15_lut_LC_6_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_15_lut_LC_6_22_5  (
            .in0(_gnd_net_),
            .in1(N__45647),
            .in2(N__27060),
            .in3(N__27036),
            .lcout(\nx.n2864 ),
            .ltout(),
            .carryin(\nx.n10825 ),
            .carryout(\nx.n10826 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_16_lut_LC_6_22_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_16_lut_LC_6_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_16_lut_LC_6_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_16_lut_LC_6_22_6  (
            .in0(_gnd_net_),
            .in1(N__45550),
            .in2(N__29903),
            .in3(N__27033),
            .lcout(\nx.n2863 ),
            .ltout(),
            .carryin(\nx.n10826 ),
            .carryout(\nx.n10827 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_17_lut_LC_6_22_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_17_lut_LC_6_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_17_lut_LC_6_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_17_lut_LC_6_22_7  (
            .in0(_gnd_net_),
            .in1(N__45648),
            .in2(N__27284),
            .in3(N__27246),
            .lcout(\nx.n2862 ),
            .ltout(),
            .carryin(\nx.n10827 ),
            .carryout(\nx.n10828 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_18_lut_LC_6_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_18_lut_LC_6_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_18_lut_LC_6_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_18_lut_LC_6_23_0  (
            .in0(_gnd_net_),
            .in1(N__45530),
            .in2(N__29681),
            .in3(N__27243),
            .lcout(\nx.n2861 ),
            .ltout(),
            .carryin(bfn_6_23_0_),
            .carryout(\nx.n10829 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_19_lut_LC_6_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_19_lut_LC_6_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_19_lut_LC_6_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_19_lut_LC_6_23_1  (
            .in0(_gnd_net_),
            .in1(N__45533),
            .in2(N__29427),
            .in3(N__27240),
            .lcout(\nx.n2860 ),
            .ltout(),
            .carryin(\nx.n10829 ),
            .carryout(\nx.n10830 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_20_lut_LC_6_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_20_lut_LC_6_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_20_lut_LC_6_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_20_lut_LC_6_23_2  (
            .in0(_gnd_net_),
            .in1(N__45531),
            .in2(N__29396),
            .in3(N__27237),
            .lcout(\nx.n2859 ),
            .ltout(),
            .carryin(\nx.n10830 ),
            .carryout(\nx.n10831 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_21_lut_LC_6_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_21_lut_LC_6_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_21_lut_LC_6_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_21_lut_LC_6_23_3  (
            .in0(_gnd_net_),
            .in1(N__45534),
            .in2(N__29412),
            .in3(N__27234),
            .lcout(\nx.n2858 ),
            .ltout(),
            .carryin(\nx.n10831 ),
            .carryout(\nx.n10832 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_22_lut_LC_6_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_22_lut_LC_6_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_22_lut_LC_6_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_22_lut_LC_6_23_4  (
            .in0(_gnd_net_),
            .in1(N__45532),
            .in2(N__30329),
            .in3(N__27231),
            .lcout(\nx.n2857 ),
            .ltout(),
            .carryin(\nx.n10832 ),
            .carryout(\nx.n10833 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_23_lut_LC_6_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_23_lut_LC_6_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_23_lut_LC_6_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_23_lut_LC_6_23_5  (
            .in0(_gnd_net_),
            .in1(N__45535),
            .in2(N__29934),
            .in3(N__27228),
            .lcout(\nx.n2856 ),
            .ltout(),
            .carryin(\nx.n10833 ),
            .carryout(\nx.n10834 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_24_lut_LC_6_23_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_24_lut_LC_6_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_24_lut_LC_6_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_24_lut_LC_6_23_6  (
            .in0(_gnd_net_),
            .in1(N__29618),
            .in2(N__45728),
            .in3(N__27225),
            .lcout(\nx.n2855 ),
            .ltout(),
            .carryin(\nx.n10834 ),
            .carryout(\nx.n10835 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_25_lut_LC_6_23_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_25_lut_LC_6_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_25_lut_LC_6_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_25_lut_LC_6_23_7  (
            .in0(_gnd_net_),
            .in1(N__45539),
            .in2(N__36465),
            .in3(N__27222),
            .lcout(\nx.n2854 ),
            .ltout(),
            .carryin(\nx.n10835 ),
            .carryout(\nx.n10836 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_26_lut_LC_6_24_0 .C_ON=1'b0;
    defparam \nx.mod_5_add_1942_26_lut_LC_6_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_26_lut_LC_6_24_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1942_26_lut_LC_6_24_0  (
            .in0(N__45338),
            .in1(N__29370),
            .in2(N__30283),
            .in3(N__27582),
            .lcout(\nx.n2885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1882_3_lut_LC_6_24_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1882_3_lut_LC_6_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1882_3_lut_LC_6_24_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1882_3_lut_LC_6_24_1  (
            .in0(_gnd_net_),
            .in1(N__29325),
            .in2(N__33906),
            .in3(N__36595),
            .lcout(\nx.n2791 ),
            .ltout(\nx.n2791_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1949_3_lut_LC_6_24_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1949_3_lut_LC_6_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1949_3_lut_LC_6_24_2 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.mod_5_i1949_3_lut_LC_6_24_2  (
            .in0(N__30246),
            .in1(N__27558),
            .in2(N__27552),
            .in3(_gnd_net_),
            .lcout(\nx.n2890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1819_3_lut_LC_6_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1819_3_lut_LC_6_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1819_3_lut_LC_6_24_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1819_3_lut_LC_6_24_3  (
            .in0(_gnd_net_),
            .in1(N__33753),
            .in2(N__37704),
            .in3(N__36208),
            .lcout(\nx.n2696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1950_3_lut_LC_6_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1950_3_lut_LC_6_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1950_3_lut_LC_6_24_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1950_3_lut_LC_6_24_4  (
            .in0(_gnd_net_),
            .in1(N__29397),
            .in2(N__30284),
            .in3(N__27549),
            .lcout(\nx.n2891 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1880_3_lut_LC_6_24_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1880_3_lut_LC_6_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1880_3_lut_LC_6_24_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1880_3_lut_LC_6_24_5  (
            .in0(_gnd_net_),
            .in1(N__36594),
            .in2(N__31668),
            .in3(N__29310),
            .lcout(\nx.n2789 ),
            .ltout(\nx.n2789_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1947_3_lut_LC_6_24_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1947_3_lut_LC_6_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1947_3_lut_LC_6_24_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.mod_5_i1947_3_lut_LC_6_24_6  (
            .in0(N__30250),
            .in1(N__27513),
            .in2(N__27507),
            .in3(_gnd_net_),
            .lcout(\nx.n2888 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_LC_6_25_0 .C_ON=1'b0;
    defparam \nx.i1_2_lut_LC_6_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_LC_6_25_0 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i1_2_lut_LC_6_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30573),
            .in3(N__30519),
            .lcout(\nx.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2089_3_lut_LC_6_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2089_3_lut_LC_6_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2089_3_lut_LC_6_25_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2089_3_lut_LC_6_25_1  (
            .in0(_gnd_net_),
            .in1(N__27504),
            .in2(N__27480),
            .in3(N__27457),
            .lcout(\nx.n3094 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_64_LC_6_25_3 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_64_LC_6_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_64_LC_6_25_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_64_LC_6_25_3  (
            .in0(N__30547),
            .in1(N__30687),
            .in2(N__27777),
            .in3(N__32409),
            .lcout(),
            .ltout(\nx.n28_adj_660_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_81_LC_6_25_4 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_81_LC_6_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_81_LC_6_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_81_LC_6_25_4  (
            .in0(N__32449),
            .in1(N__27594),
            .in2(N__27609),
            .in3(N__27606),
            .lcout(\nx.n1928 ),
            .ltout(\nx.n1928_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9586_1_lut_LC_6_25_5 .C_ON=1'b0;
    defparam \nx.i9586_1_lut_LC_6_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9586_1_lut_LC_6_25_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \nx.i9586_1_lut_LC_6_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27600),
            .in3(_gnd_net_),
            .lcout(\nx.n13435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1283_3_lut_LC_6_25_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1283_3_lut_LC_6_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1283_3_lut_LC_6_25_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1283_3_lut_LC_6_25_7  (
            .in0(_gnd_net_),
            .in1(N__32538),
            .in2(N__32511),
            .in3(N__32887),
            .lcout(\nx.n1904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1287_3_lut_LC_6_26_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1287_3_lut_LC_6_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1287_3_lut_LC_6_26_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1287_3_lut_LC_6_26_0  (
            .in0(N__32643),
            .in1(_gnd_net_),
            .in2(N__32900),
            .in3(N__32662),
            .lcout(\nx.n1908 ),
            .ltout(\nx.n1908_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_55_LC_6_26_1 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_55_LC_6_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_55_LC_6_26_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_adj_55_LC_6_26_1  (
            .in0(N__30658),
            .in1(N__30007),
            .in2(N__27597),
            .in3(N__32356),
            .lcout(\nx.n24_adj_648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1286_3_lut_LC_6_26_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1286_3_lut_LC_6_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1286_3_lut_LC_6_26_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1286_3_lut_LC_6_26_2  (
            .in0(_gnd_net_),
            .in1(N__32607),
            .in2(N__32899),
            .in3(N__32624),
            .lcout(\nx.n1907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1288_3_lut_LC_6_26_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1288_3_lut_LC_6_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1288_3_lut_LC_6_26_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1288_3_lut_LC_6_26_3  (
            .in0(N__27588),
            .in1(N__32764),
            .in2(_gnd_net_),
            .in3(N__32874),
            .lcout(\nx.n1909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_16_LC_6_26_4 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_16_LC_6_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_16_LC_6_26_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_16_LC_6_26_4  (
            .in0(N__32588),
            .in1(N__32623),
            .in2(N__32400),
            .in3(N__27744),
            .lcout(\nx.n1829 ),
            .ltout(\nx.n1829_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1282_3_lut_LC_6_26_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1282_3_lut_LC_6_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1282_3_lut_LC_6_26_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \nx.mod_5_i1282_3_lut_LC_6_26_5  (
            .in0(N__32486),
            .in1(N__32472),
            .in2(N__27783),
            .in3(_gnd_net_),
            .lcout(\nx.n1903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1285_3_lut_LC_6_26_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1285_3_lut_LC_6_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1285_3_lut_LC_6_26_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i1285_3_lut_LC_6_26_6  (
            .in0(N__32878),
            .in1(_gnd_net_),
            .in2(N__32592),
            .in3(N__32568),
            .lcout(\nx.n1906 ),
            .ltout(\nx.n1906_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_3_lut_LC_6_26_7 .C_ON=1'b0;
    defparam \nx.i7_3_lut_LC_6_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.i7_3_lut_LC_6_26_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i7_3_lut_LC_6_26_7  (
            .in0(_gnd_net_),
            .in1(N__30108),
            .in2(N__27780),
            .in3(N__30061),
            .lcout(\nx.n22_adj_605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9569_2_lut_LC_6_27_0 .C_ON=1'b0;
    defparam \nx.i9569_2_lut_LC_6_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.i9569_2_lut_LC_6_27_0 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \nx.i9569_2_lut_LC_6_27_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27957),
            .in3(N__30643),
            .lcout(\nx.n1006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1215_3_lut_LC_6_27_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1215_3_lut_LC_6_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1215_3_lut_LC_6_27_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1215_3_lut_LC_6_27_1  (
            .in0(_gnd_net_),
            .in1(N__34716),
            .in2(N__34749),
            .in3(N__35151),
            .lcout(\nx.n1804 ),
            .ltout(\nx.n1804_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_3_lut_adj_132_LC_6_27_2 .C_ON=1'b0;
    defparam \nx.i5_3_lut_adj_132_LC_6_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.i5_3_lut_adj_132_LC_6_27_2 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i5_3_lut_adj_132_LC_6_27_2  (
            .in0(_gnd_net_),
            .in1(N__32769),
            .in2(N__27750),
            .in3(N__32666),
            .lcout(),
            .ltout(\nx.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_15_LC_6_27_3 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_15_LC_6_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_15_LC_6_27_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_15_LC_6_27_3  (
            .in0(N__34613),
            .in1(N__32530),
            .in2(N__27747),
            .in3(N__30861),
            .lcout(\nx.n26_adj_600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2045_2_lut_3_lut_LC_6_27_4 .C_ON=1'b0;
    defparam \nx.i2045_2_lut_3_lut_LC_6_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.i2045_2_lut_3_lut_LC_6_27_4 .LUT_INIT=16'b1100000000001100;
    LogicCell40 \nx.i2045_2_lut_3_lut_LC_6_27_4  (
            .in0(_gnd_net_),
            .in1(N__27738),
            .in2(N__27690),
            .in3(N__27635),
            .lcout(\nx.n5260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1278_3_lut_LC_6_27_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1278_3_lut_LC_6_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1278_3_lut_LC_6_27_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1278_3_lut_LC_6_27_5  (
            .in0(N__33020),
            .in1(_gnd_net_),
            .in2(N__33000),
            .in3(N__32882),
            .lcout(\nx.n1899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_2_lut_LC_6_28_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_2_lut_LC_6_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_2_lut_LC_6_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_2_lut_LC_6_28_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28071),
            .in3(N__28017),
            .lcout(\nx.n977 ),
            .ltout(),
            .carryin(bfn_6_28_0_),
            .carryout(\nx.n10474 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_3_lut_LC_6_28_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_3_lut_LC_6_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_3_lut_LC_6_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_3_lut_LC_6_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28014),
            .in3(N__27990),
            .lcout(\nx.n976 ),
            .ltout(),
            .carryin(\nx.n10474 ),
            .carryout(\nx.n10475 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_4_lut_LC_6_28_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_4_lut_LC_6_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_4_lut_LC_6_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_4_lut_LC_6_28_2  (
            .in0(_gnd_net_),
            .in1(N__45099),
            .in2(N__27987),
            .in3(N__27960),
            .lcout(\nx.n975 ),
            .ltout(),
            .carryin(\nx.n10475 ),
            .carryout(\nx.n10476 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_5_lut_LC_6_28_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_5_lut_LC_6_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_5_lut_LC_6_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_5_lut_LC_6_28_3  (
            .in0(_gnd_net_),
            .in1(N__45104),
            .in2(N__27798),
            .in3(N__27942),
            .lcout(\nx.n974 ),
            .ltout(),
            .carryin(\nx.n10476 ),
            .carryout(\nx.n10477 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_6_lut_LC_6_28_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_6_lut_LC_6_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_6_lut_LC_6_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_6_lut_LC_6_28_4  (
            .in0(_gnd_net_),
            .in1(N__45100),
            .in2(N__27938),
            .in3(N__27909),
            .lcout(\nx.n973 ),
            .ltout(),
            .carryin(\nx.n10477 ),
            .carryout(\nx.n10478 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_7_lut_LC_6_28_5 .C_ON=1'b0;
    defparam \nx.mod_5_add_669_7_lut_LC_6_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_7_lut_LC_6_28_5 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_669_7_lut_LC_6_28_5  (
            .in0(N__27906),
            .in1(N__30597),
            .in2(N__45496),
            .in3(N__27894),
            .lcout(\nx.n4_adj_596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1152_3_lut_LC_6_28_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1152_3_lut_LC_6_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1152_3_lut_LC_6_28_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1152_3_lut_LC_6_28_6  (
            .in0(N__30957),
            .in1(N__31005),
            .in2(_gnd_net_),
            .in3(N__34480),
            .lcout(\nx.n1709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i606_3_lut_LC_6_28_7 .C_ON=1'b0;
    defparam \nx.mod_5_i606_3_lut_LC_6_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i606_3_lut_LC_6_28_7 .LUT_INIT=16'b1111000011000011;
    LogicCell40 \nx.mod_5_i606_3_lut_LC_6_28_7  (
            .in0(_gnd_net_),
            .in1(N__27871),
            .in2(N__27855),
            .in3(N__27823),
            .lcout(\nx.n11674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_41_LC_6_29_0 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_41_LC_6_29_0 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_41_LC_6_29_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_41_LC_6_29_0  (
            .in0(N__28475),
            .in1(N__28143),
            .in2(N__28398),
            .in3(N__28098),
            .lcout(\nx.n1532 ),
            .ltout(\nx.n1532_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1078_3_lut_LC_6_29_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1078_3_lut_LC_6_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1078_3_lut_LC_6_29_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1078_3_lut_LC_6_29_1  (
            .in0(_gnd_net_),
            .in1(N__28397),
            .in2(N__28089),
            .in3(N__28371),
            .lcout(\nx.n1603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1081_3_lut_LC_6_29_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1081_3_lut_LC_6_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1081_3_lut_LC_6_29_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1081_3_lut_LC_6_29_2  (
            .in0(N__28476),
            .in1(_gnd_net_),
            .in2(N__28455),
            .in3(N__33263),
            .lcout(\nx.n1606 ),
            .ltout(\nx.n1606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_54_LC_6_29_3 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_54_LC_6_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_54_LC_6_29_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_54_LC_6_29_3  (
            .in0(N__31156),
            .in1(N__28077),
            .in2(N__28086),
            .in3(N__30801),
            .lcout(),
            .ltout(\nx.n22_adj_647_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_80_LC_6_29_4 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_80_LC_6_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_80_LC_6_29_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_80_LC_6_29_4  (
            .in0(N__33172),
            .in1(N__30910),
            .in2(N__28083),
            .in3(N__33321),
            .lcout(\nx.n1631 ),
            .ltout(\nx.n1631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1147_3_lut_LC_6_29_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1147_3_lut_LC_6_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1147_3_lut_LC_6_29_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1147_3_lut_LC_6_29_5  (
            .in0(_gnd_net_),
            .in1(N__33203),
            .in2(N__28080),
            .in3(N__30876),
            .lcout(\nx.n1704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1082_3_lut_LC_6_29_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1082_3_lut_LC_6_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1082_3_lut_LC_6_29_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1082_3_lut_LC_6_29_6  (
            .in0(_gnd_net_),
            .in1(N__28110),
            .in2(N__28128),
            .in3(N__33262),
            .lcout(\nx.n1607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1079_3_lut_LC_6_29_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1079_3_lut_LC_6_29_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1079_3_lut_LC_6_29_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1079_3_lut_LC_6_29_7  (
            .in0(N__28410),
            .in1(_gnd_net_),
            .in2(N__33275),
            .in3(N__28437),
            .lcout(\nx.n1604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_4_lut_LC_6_30_0 .C_ON=1'b0;
    defparam \nx.i7_4_lut_LC_6_30_0 .SEQ_MODE=4'b0000;
    defparam \nx.i7_4_lut_LC_6_30_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i7_4_lut_LC_6_30_0  (
            .in0(N__31109),
            .in1(N__33385),
            .in2(N__31070),
            .in3(N__31089),
            .lcout(\nx.n19_adj_602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1076_3_lut_LC_6_30_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1076_3_lut_LC_6_30_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1076_3_lut_LC_6_30_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1076_3_lut_LC_6_30_1  (
            .in0(_gnd_net_),
            .in1(N__28355),
            .in2(N__33272),
            .in3(N__28335),
            .lcout(\nx.n1601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1075_3_lut_LC_6_30_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1075_3_lut_LC_6_30_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1075_3_lut_LC_6_30_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1075_3_lut_LC_6_30_2  (
            .in0(N__28323),
            .in1(_gnd_net_),
            .in2(N__28302),
            .in3(N__33255),
            .lcout(\nx.n1600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1015_3_lut_LC_6_30_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1015_3_lut_LC_6_30_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1015_3_lut_LC_6_30_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1015_3_lut_LC_6_30_3  (
            .in0(_gnd_net_),
            .in1(N__28248),
            .in2(N__28224),
            .in3(N__28209),
            .lcout(\nx.n1508 ),
            .ltout(\nx.n1508_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_2_lut_LC_6_30_4 .C_ON=1'b0;
    defparam \nx.i5_2_lut_LC_6_30_4 .SEQ_MODE=4'b0000;
    defparam \nx.i5_2_lut_LC_6_30_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i5_2_lut_LC_6_30_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28146),
            .in3(N__28433),
            .lcout(\nx.n16_adj_633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_3_lut_adj_91_LC_6_30_5 .C_ON=1'b0;
    defparam \nx.i7_3_lut_adj_91_LC_6_30_5 .SEQ_MODE=4'b0000;
    defparam \nx.i7_3_lut_adj_91_LC_6_30_5 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \nx.i7_3_lut_adj_91_LC_6_30_5  (
            .in0(_gnd_net_),
            .in1(N__35063),
            .in2(N__35425),
            .in3(N__35185),
            .lcout(\nx.n20_adj_680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1074_3_lut_LC_6_30_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1074_3_lut_LC_6_30_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1074_3_lut_LC_6_30_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1074_3_lut_LC_6_30_6  (
            .in0(_gnd_net_),
            .in1(N__28287),
            .in2(N__28263),
            .in3(N__33251),
            .lcout(\nx.n1599 ),
            .ltout(\nx.n1599_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1141_3_lut_LC_6_30_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1141_3_lut_LC_6_30_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1141_3_lut_LC_6_30_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1141_3_lut_LC_6_30_7  (
            .in0(_gnd_net_),
            .in1(N__34499),
            .in2(N__28137),
            .in3(N__31098),
            .lcout(\nx.n1698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_2_lut_LC_6_31_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_2_lut_LC_6_31_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_2_lut_LC_6_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_2_lut_LC_6_31_0  (
            .in0(_gnd_net_),
            .in1(N__30845),
            .in2(_gnd_net_),
            .in3(N__28134),
            .lcout(\nx.n1577 ),
            .ltout(),
            .carryin(bfn_6_31_0_),
            .carryout(\nx.n10592 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_3_lut_LC_6_31_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_3_lut_LC_6_31_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_3_lut_LC_6_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_3_lut_LC_6_31_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33362),
            .in3(N__28131),
            .lcout(\nx.n1576 ),
            .ltout(),
            .carryin(\nx.n10592 ),
            .carryout(\nx.n10593 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_4_lut_LC_6_31_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_4_lut_LC_6_31_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_4_lut_LC_6_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_4_lut_LC_6_31_2  (
            .in0(_gnd_net_),
            .in1(N__44869),
            .in2(N__28127),
            .in3(N__28101),
            .lcout(\nx.n1575 ),
            .ltout(),
            .carryin(\nx.n10593 ),
            .carryout(\nx.n10594 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_5_lut_LC_6_31_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_5_lut_LC_6_31_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_5_lut_LC_6_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_5_lut_LC_6_31_3  (
            .in0(_gnd_net_),
            .in1(N__44923),
            .in2(N__28474),
            .in3(N__28443),
            .lcout(\nx.n1574 ),
            .ltout(),
            .carryin(\nx.n10594 ),
            .carryout(\nx.n10595 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_6_lut_LC_6_31_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_6_lut_LC_6_31_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_6_lut_LC_6_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_6_lut_LC_6_31_4  (
            .in0(_gnd_net_),
            .in1(N__44870),
            .in2(N__33308),
            .in3(N__28440),
            .lcout(\nx.n1573 ),
            .ltout(),
            .carryin(\nx.n10595 ),
            .carryout(\nx.n10596 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_7_lut_LC_6_31_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_7_lut_LC_6_31_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_7_lut_LC_6_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_7_lut_LC_6_31_5  (
            .in0(_gnd_net_),
            .in1(N__44924),
            .in2(N__28432),
            .in3(N__28401),
            .lcout(\nx.n1572 ),
            .ltout(),
            .carryin(\nx.n10596 ),
            .carryout(\nx.n10597 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_8_lut_LC_6_31_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_8_lut_LC_6_31_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_8_lut_LC_6_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_8_lut_LC_6_31_6  (
            .in0(_gnd_net_),
            .in1(N__44871),
            .in2(N__28393),
            .in3(N__28362),
            .lcout(\nx.n1571 ),
            .ltout(),
            .carryin(\nx.n10597 ),
            .carryout(\nx.n10598 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_9_lut_LC_6_31_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_9_lut_LC_6_31_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_9_lut_LC_6_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_9_lut_LC_6_31_7  (
            .in0(_gnd_net_),
            .in1(N__44925),
            .in2(N__31032),
            .in3(N__28359),
            .lcout(\nx.n1570 ),
            .ltout(),
            .carryin(\nx.n10598 ),
            .carryout(\nx.n10599 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_10_lut_LC_6_32_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_10_lut_LC_6_32_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_10_lut_LC_6_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_10_lut_LC_6_32_0  (
            .in0(_gnd_net_),
            .in1(N__44483),
            .in2(N__28356),
            .in3(N__28326),
            .lcout(\nx.n1569 ),
            .ltout(),
            .carryin(bfn_6_32_0_),
            .carryout(\nx.n10600 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_11_lut_LC_6_32_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_11_lut_LC_6_32_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_11_lut_LC_6_32_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_11_lut_LC_6_32_1  (
            .in0(_gnd_net_),
            .in1(N__44486),
            .in2(N__28322),
            .in3(N__28290),
            .lcout(\nx.n1568 ),
            .ltout(),
            .carryin(\nx.n10600 ),
            .carryout(\nx.n10601 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_12_lut_LC_6_32_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_12_lut_LC_6_32_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_12_lut_LC_6_32_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1071_12_lut_LC_6_32_2  (
            .in0(_gnd_net_),
            .in1(N__44484),
            .in2(N__28286),
            .in3(N__28251),
            .lcout(\nx.n1567 ),
            .ltout(),
            .carryin(\nx.n10601 ),
            .carryout(\nx.n10602 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_13_lut_LC_6_32_3 .C_ON=1'b0;
    defparam \nx.mod_5_add_1071_13_lut_LC_6_32_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_13_lut_LC_6_32_3 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1071_13_lut_LC_6_32_3  (
            .in0(N__44485),
            .in1(N__28941),
            .in2(N__33276),
            .in3(N__28920),
            .lcout(\nx.n1598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i0_LC_7_16_5.C_ON=1'b0;
    defparam pin_output_i0_i0_LC_7_16_5.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i0_LC_7_16_5.LUT_INIT=16'b0101000011011000;
    LogicCell40 pin_output_i0_i0_LC_7_16_5 (
            .in0(N__31254),
            .in1(N__35472),
            .in2(N__28613),
            .in3(N__46536),
            .lcout(pin_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48411),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1825_3_lut_LC_7_17_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1825_3_lut_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1825_3_lut_LC_7_17_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1825_3_lut_LC_7_17_0  (
            .in0(N__36687),
            .in1(_gnd_net_),
            .in2(N__33615),
            .in3(N__36207),
            .lcout(\nx.n2702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i13_LC_7_17_1.C_ON=1'b0;
    defparam neopxl_color_i13_LC_7_17_1.SEQ_MODE=4'b1000;
    defparam neopxl_color_i13_LC_7_17_1.LUT_INIT=16'b1101111100000100;
    LogicCell40 neopxl_color_i13_LC_7_17_1 (
            .in0(N__49842),
            .in1(N__49593),
            .in2(N__50077),
            .in3(N__28897),
            .lcout(neopxl_color_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48406),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i0_LC_7_17_2 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i0_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i0_LC_7_17_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i0_LC_7_17_2  (
            .in0(N__28874),
            .in1(N__28673),
            .in2(_gnd_net_),
            .in3(N__28647),
            .lcout(neo_pixel_transmitter_t0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48406),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i1_LC_7_17_4.C_ON=1'b0;
    defparam pin_output_i0_i1_LC_7_17_4.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i1_LC_7_17_4.LUT_INIT=16'b0101000011011000;
    LogicCell40 pin_output_i0_i1_LC_7_17_4 (
            .in0(N__31242),
            .in1(N__33105),
            .in2(N__28571),
            .in3(N__46515),
            .lcout(pin_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48406),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i1_1_lut_LC_7_18_0 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i1_1_lut_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i1_1_lut_LC_7_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i1_1_lut_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28646),
            .lcout(\nx.n33_adj_652 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9299_3_lut_LC_7_18_4.C_ON=1'b0;
    defparam i9299_3_lut_LC_7_18_4.SEQ_MODE=4'b0000;
    defparam i9299_3_lut_LC_7_18_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i9299_3_lut_LC_7_18_4 (
            .in0(N__28612),
            .in1(N__28564),
            .in2(_gnd_net_),
            .in3(N__49041),
            .lcout(n13146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_2_lut_LC_7_19_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_2_lut_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_2_lut_LC_7_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_2_lut_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__28548),
            .in2(_gnd_net_),
            .in3(N__28479),
            .lcout(\nx.n2777 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\nx.n10790 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_3_lut_LC_7_19_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_3_lut_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_3_lut_LC_7_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_3_lut_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31453),
            .in3(N__29109),
            .lcout(\nx.n2776 ),
            .ltout(),
            .carryin(\nx.n10790 ),
            .carryout(\nx.n10791 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_4_lut_LC_7_19_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_4_lut_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_4_lut_LC_7_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_4_lut_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__45695),
            .in2(N__29105),
            .in3(N__29076),
            .lcout(\nx.n2775 ),
            .ltout(),
            .carryin(\nx.n10791 ),
            .carryout(\nx.n10792 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_5_lut_LC_7_19_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_5_lut_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_5_lut_LC_7_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_5_lut_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__45698),
            .in2(N__29068),
            .in3(N__29037),
            .lcout(\nx.n2774 ),
            .ltout(),
            .carryin(\nx.n10792 ),
            .carryout(\nx.n10793 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_6_lut_LC_7_19_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_6_lut_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_6_lut_LC_7_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_6_lut_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__45696),
            .in2(N__29034),
            .in3(N__29001),
            .lcout(\nx.n2773 ),
            .ltout(),
            .carryin(\nx.n10793 ),
            .carryout(\nx.n10794 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_7_lut_LC_7_19_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_7_lut_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_7_lut_LC_7_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_7_lut_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__45699),
            .in2(N__36081),
            .in3(N__28998),
            .lcout(\nx.n2772 ),
            .ltout(),
            .carryin(\nx.n10794 ),
            .carryout(\nx.n10795 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_8_lut_LC_7_19_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_8_lut_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_8_lut_LC_7_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_8_lut_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__45697),
            .in2(N__31568),
            .in3(N__28989),
            .lcout(\nx.n2771 ),
            .ltout(),
            .carryin(\nx.n10795 ),
            .carryout(\nx.n10796 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_9_lut_LC_7_19_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_9_lut_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_9_lut_LC_7_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_9_lut_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__45700),
            .in2(N__31481),
            .in3(N__28980),
            .lcout(\nx.n2770 ),
            .ltout(),
            .carryin(\nx.n10796 ),
            .carryout(\nx.n10797 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_10_lut_LC_7_20_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_10_lut_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_10_lut_LC_7_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_10_lut_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__45016),
            .in2(N__28977),
            .in3(N__28944),
            .lcout(\nx.n2769 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\nx.n10798 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_11_lut_LC_7_20_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_11_lut_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_11_lut_LC_7_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_11_lut_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__45649),
            .in2(N__31598),
            .in3(N__29235),
            .lcout(\nx.n2768 ),
            .ltout(),
            .carryin(\nx.n10798 ),
            .carryout(\nx.n10799 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_12_lut_LC_7_20_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_12_lut_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_12_lut_LC_7_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_12_lut_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(N__45017),
            .in2(N__29231),
            .in3(N__29205),
            .lcout(\nx.n2767 ),
            .ltout(),
            .carryin(\nx.n10799 ),
            .carryout(\nx.n10800 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_13_lut_LC_7_20_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_13_lut_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_13_lut_LC_7_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_13_lut_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(N__45650),
            .in2(N__33809),
            .in3(N__29196),
            .lcout(\nx.n2766 ),
            .ltout(),
            .carryin(\nx.n10800 ),
            .carryout(\nx.n10801 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_14_lut_LC_7_20_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_14_lut_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_14_lut_LC_7_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_14_lut_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(N__31511),
            .in2(N__45752),
            .in3(N__29187),
            .lcout(\nx.n2765 ),
            .ltout(),
            .carryin(\nx.n10801 ),
            .carryout(\nx.n10802 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_15_lut_LC_7_20_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_15_lut_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_15_lut_LC_7_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_15_lut_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__45654),
            .in2(N__31287),
            .in3(N__29175),
            .lcout(\nx.n2764 ),
            .ltout(),
            .carryin(\nx.n10802 ),
            .carryout(\nx.n10803 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_16_lut_LC_7_20_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_16_lut_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_16_lut_LC_7_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_16_lut_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__45018),
            .in2(N__29172),
            .in3(N__29133),
            .lcout(\nx.n2763 ),
            .ltout(),
            .carryin(\nx.n10803 ),
            .carryout(\nx.n10804 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_17_lut_LC_7_20_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_17_lut_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_17_lut_LC_7_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_17_lut_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(N__45655),
            .in2(N__31542),
            .in3(N__29124),
            .lcout(\nx.n2762 ),
            .ltout(),
            .carryin(\nx.n10804 ),
            .carryout(\nx.n10805 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_18_lut_LC_7_21_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_18_lut_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_18_lut_LC_7_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_18_lut_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__31316),
            .in2(N__45751),
            .in3(N__29121),
            .lcout(\nx.n2761 ),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\nx.n10806 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_19_lut_LC_7_21_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_19_lut_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_19_lut_LC_7_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_19_lut_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__45642),
            .in2(N__33858),
            .in3(N__29328),
            .lcout(\nx.n2760 ),
            .ltout(),
            .carryin(\nx.n10806 ),
            .carryout(\nx.n10807 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_20_lut_LC_7_21_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_20_lut_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_20_lut_LC_7_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_20_lut_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(N__45691),
            .in2(N__33902),
            .in3(N__29316),
            .lcout(\nx.n2759 ),
            .ltout(),
            .carryin(\nx.n10807 ),
            .carryout(\nx.n10808 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_21_lut_LC_7_21_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_21_lut_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_21_lut_LC_7_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_21_lut_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__45643),
            .in2(N__31628),
            .in3(N__29313),
            .lcout(\nx.n2758 ),
            .ltout(),
            .carryin(\nx.n10808 ),
            .carryout(\nx.n10809 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_22_lut_LC_7_21_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_22_lut_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_22_lut_LC_7_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_22_lut_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(N__45692),
            .in2(N__31667),
            .in3(N__29301),
            .lcout(\nx.n2757 ),
            .ltout(),
            .carryin(\nx.n10809 ),
            .carryout(\nx.n10810 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_23_lut_LC_7_21_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_23_lut_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_23_lut_LC_7_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_23_lut_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__45644),
            .in2(N__31692),
            .in3(N__29292),
            .lcout(\nx.n2756 ),
            .ltout(),
            .carryin(\nx.n10810 ),
            .carryout(\nx.n10811 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_24_lut_LC_7_21_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_24_lut_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_24_lut_LC_7_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_24_lut_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(N__45693),
            .in2(N__36636),
            .in3(N__29289),
            .lcout(\nx.n2755 ),
            .ltout(),
            .carryin(\nx.n10811 ),
            .carryout(\nx.n10812 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_25_lut_LC_7_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_add_1875_25_lut_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_25_lut_LC_7_21_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_1875_25_lut_LC_7_21_7  (
            .in0(N__45694),
            .in1(N__36601),
            .in2(N__33789),
            .in3(N__29286),
            .lcout(\nx.n2786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_70_LC_7_22_0 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_70_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_70_LC_7_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_adj_70_LC_7_22_0  (
            .in0(N__32182),
            .in1(N__34375),
            .in2(N__34339),
            .in3(N__32129),
            .lcout(\nx.n25_adj_666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i23_1_lut_LC_7_22_1 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i23_1_lut_LC_7_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i23_1_lut_LC_7_22_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \nx.sub_14_inv_0_i23_1_lut_LC_7_22_1  (
            .in0(N__29283),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\nx.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1884_3_lut_LC_7_22_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1884_3_lut_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1884_3_lut_LC_7_22_2 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \nx.mod_5_i1884_3_lut_LC_7_22_2  (
            .in0(N__31317),
            .in1(N__36596),
            .in2(N__29547),
            .in3(_gnd_net_),
            .lcout(\nx.n2793 ),
            .ltout(\nx.n2793_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1951_3_lut_LC_7_22_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1951_3_lut_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1951_3_lut_LC_7_22_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1951_3_lut_LC_7_22_3  (
            .in0(_gnd_net_),
            .in1(N__29538),
            .in2(N__29532),
            .in3(N__30251),
            .lcout(\nx.n2892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1881_3_lut_LC_7_22_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1881_3_lut_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1881_3_lut_LC_7_22_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1881_3_lut_LC_7_22_4  (
            .in0(N__29493),
            .in1(_gnd_net_),
            .in2(N__31629),
            .in3(N__36600),
            .lcout(\nx.n2790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1883_3_lut_LC_7_22_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1883_3_lut_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1883_3_lut_LC_7_22_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1883_3_lut_LC_7_22_5  (
            .in0(N__33857),
            .in1(_gnd_net_),
            .in2(N__36605),
            .in3(N__29487),
            .lcout(\nx.n2792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9505_3_lut_LC_7_22_6 .C_ON=1'b0;
    defparam \nx.i9505_3_lut_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9505_3_lut_LC_7_22_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.i9505_3_lut_LC_7_22_6  (
            .in0(_gnd_net_),
            .in1(N__29481),
            .in2(N__30285),
            .in3(N__29475),
            .lcout(\nx.n2905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_63_LC_7_22_7 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_63_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_63_LC_7_22_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_63_LC_7_22_7  (
            .in0(N__41060),
            .in1(N__41153),
            .in2(N__41427),
            .in3(N__43199),
            .lcout(\nx.n33_adj_659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_33_LC_7_23_0 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_33_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_33_LC_7_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_33_LC_7_23_0  (
            .in0(N__29423),
            .in1(N__29408),
            .in2(N__29395),
            .in3(N__30322),
            .lcout(),
            .ltout(\nx.n38_adj_625_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_43_LC_7_23_1 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_43_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_43_LC_7_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_43_LC_7_23_1  (
            .in0(N__29369),
            .in1(N__36457),
            .in2(N__29355),
            .in3(N__29916),
            .lcout(),
            .ltout(\nx.n43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i23_4_lut_LC_7_23_2 .C_ON=1'b0;
    defparam \nx.i23_4_lut_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.i23_4_lut_LC_7_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i23_4_lut_LC_7_23_2  (
            .in0(N__29352),
            .in1(N__29340),
            .in2(N__29331),
            .in3(N__29988),
            .lcout(\nx.n2819 ),
            .ltout(\nx.n2819_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1945_3_lut_LC_7_23_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1945_3_lut_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1945_3_lut_LC_7_23_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1945_3_lut_LC_7_23_3  (
            .in0(N__29976),
            .in1(_gnd_net_),
            .in2(N__29970),
            .in3(N__36458),
            .lcout(\nx.n2886 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2_2_lut_LC_7_23_4 .C_ON=1'b0;
    defparam \nx.i2_2_lut_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.i2_2_lut_LC_7_23_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i2_2_lut_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29933),
            .in3(N__29617),
            .lcout(\nx.n26_adj_615 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1954_3_lut_LC_7_23_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1954_3_lut_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1954_3_lut_LC_7_23_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1954_3_lut_LC_7_23_5  (
            .in0(_gnd_net_),
            .in1(N__29910),
            .in2(N__30255),
            .in3(N__29904),
            .lcout(\nx.n2895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1968_3_lut_LC_7_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1968_3_lut_LC_7_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1968_3_lut_LC_7_23_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1968_3_lut_LC_7_23_6  (
            .in0(N__29841),
            .in1(N__29829),
            .in2(_gnd_net_),
            .in3(N__30211),
            .lcout(\nx.n2909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1959_3_lut_LC_7_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1959_3_lut_LC_7_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1959_3_lut_LC_7_23_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1959_3_lut_LC_7_23_7  (
            .in0(_gnd_net_),
            .in1(N__29745),
            .in2(N__30256),
            .in3(N__29739),
            .lcout(\nx.n2900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1952_3_lut_LC_7_24_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1952_3_lut_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1952_3_lut_LC_7_24_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1952_3_lut_LC_7_24_0  (
            .in0(_gnd_net_),
            .in1(N__29688),
            .in2(N__30275),
            .in3(N__29682),
            .lcout(\nx.n2893 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1946_3_lut_LC_7_24_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1946_3_lut_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1946_3_lut_LC_7_24_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1946_3_lut_LC_7_24_2  (
            .in0(_gnd_net_),
            .in1(N__29619),
            .in2(N__30277),
            .in3(N__29595),
            .lcout(\nx.n2887 ),
            .ltout(\nx.n2887_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_90_LC_7_24_3 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_90_LC_7_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_90_LC_7_24_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_90_LC_7_24_3  (
            .in0(N__29563),
            .in1(N__30481),
            .in2(N__30465),
            .in3(N__30130),
            .lcout(\nx.n39_adj_679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1961_3_lut_LC_7_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1961_3_lut_LC_7_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1961_3_lut_LC_7_24_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1961_3_lut_LC_7_24_4  (
            .in0(_gnd_net_),
            .in1(N__30450),
            .in2(N__30274),
            .in3(N__30423),
            .lcout(\nx.n2902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1962_3_lut_LC_7_24_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1962_3_lut_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1962_3_lut_LC_7_24_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1962_3_lut_LC_7_24_5  (
            .in0(_gnd_net_),
            .in1(N__30378),
            .in2(N__36048),
            .in3(N__30227),
            .lcout(\nx.n2903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1948_3_lut_LC_7_24_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1948_3_lut_LC_7_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1948_3_lut_LC_7_24_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1948_3_lut_LC_7_24_6  (
            .in0(_gnd_net_),
            .in1(N__30330),
            .in2(N__30276),
            .in3(N__30150),
            .lcout(\nx.n2889 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_67_LC_7_24_7 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_67_LC_7_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_67_LC_7_24_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_67_LC_7_24_7  (
            .in0(N__31984),
            .in1(N__34276),
            .in2(N__32089),
            .in3(N__32032),
            .lcout(\nx.n28_adj_663 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_2_lut_LC_7_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_2_lut_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_2_lut_LC_7_25_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1339_2_lut_LC_7_25_0  (
            .in0(N__30117),
            .in1(N__30116),
            .in2(N__30044),
            .in3(N__30066),
            .lcout(\nx.n2009 ),
            .ltout(),
            .carryin(bfn_7_25_0_),
            .carryout(\nx.n10642 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_3_lut_LC_7_25_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_3_lut_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_3_lut_LC_7_25_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1339_3_lut_LC_7_25_1  (
            .in0(N__30063),
            .in1(N__30062),
            .in2(N__30045),
            .in3(N__30027),
            .lcout(\nx.n2008 ),
            .ltout(),
            .carryin(\nx.n10642 ),
            .carryout(\nx.n10643 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_4_lut_LC_7_25_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_4_lut_LC_7_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_4_lut_LC_7_25_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_4_lut_LC_7_25_2  (
            .in0(N__30024),
            .in1(N__30023),
            .in2(N__30773),
            .in3(N__30012),
            .lcout(\nx.n2007 ),
            .ltout(),
            .carryin(\nx.n10643 ),
            .carryout(\nx.n10644 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_5_lut_LC_7_25_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_5_lut_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_5_lut_LC_7_25_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_5_lut_LC_7_25_3  (
            .in0(N__30009),
            .in1(N__30008),
            .in2(N__30776),
            .in3(N__29991),
            .lcout(\nx.n2006 ),
            .ltout(),
            .carryin(\nx.n10644 ),
            .carryout(\nx.n10645 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_6_lut_LC_7_25_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_6_lut_LC_7_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_6_lut_LC_7_25_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_6_lut_LC_7_25_4  (
            .in0(N__30591),
            .in1(N__30590),
            .in2(N__30774),
            .in3(N__30579),
            .lcout(\nx.n2005 ),
            .ltout(),
            .carryin(\nx.n10645 ),
            .carryout(\nx.n10646 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_7_lut_LC_7_25_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_7_lut_LC_7_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_7_lut_LC_7_25_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_7_lut_LC_7_25_5  (
            .in0(N__32430),
            .in1(N__32429),
            .in2(N__30777),
            .in3(N__30576),
            .lcout(\nx.n2004 ),
            .ltout(),
            .carryin(\nx.n10646 ),
            .carryout(\nx.n10647 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_8_lut_LC_7_25_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_8_lut_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_8_lut_LC_7_25_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_8_lut_LC_7_25_6  (
            .in0(N__30572),
            .in1(N__30571),
            .in2(N__30775),
            .in3(N__30552),
            .lcout(\nx.n2003 ),
            .ltout(),
            .carryin(\nx.n10647 ),
            .carryout(\nx.n10648 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_9_lut_LC_7_25_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_9_lut_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_9_lut_LC_7_25_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_9_lut_LC_7_25_7  (
            .in0(N__30549),
            .in1(N__30548),
            .in2(N__30778),
            .in3(N__30531),
            .lcout(\nx.n2002 ),
            .ltout(),
            .carryin(\nx.n10648 ),
            .carryout(\nx.n10649 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_10_lut_LC_7_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_10_lut_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_10_lut_LC_7_26_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_10_lut_LC_7_26_0  (
            .in0(N__30666),
            .in1(N__30665),
            .in2(N__30779),
            .in3(N__30528),
            .lcout(\nx.n2001 ),
            .ltout(),
            .carryin(bfn_7_26_0_),
            .carryout(\nx.n10650 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_11_lut_LC_7_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_11_lut_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_11_lut_LC_7_26_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_11_lut_LC_7_26_1  (
            .in0(N__32457),
            .in1(N__32456),
            .in2(N__30783),
            .in3(N__30525),
            .lcout(\nx.n2000 ),
            .ltout(),
            .carryin(\nx.n10650 ),
            .carryout(\nx.n10651 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_12_lut_LC_7_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_12_lut_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_12_lut_LC_7_26_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_12_lut_LC_7_26_2  (
            .in0(N__32388),
            .in1(N__32387),
            .in2(N__30780),
            .in3(N__30522),
            .lcout(\nx.n1999 ),
            .ltout(),
            .carryin(\nx.n10651 ),
            .carryout(\nx.n10652 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_13_lut_LC_7_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_13_lut_LC_7_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_13_lut_LC_7_26_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_13_lut_LC_7_26_3  (
            .in0(N__30518),
            .in1(N__30517),
            .in2(N__30784),
            .in3(N__30498),
            .lcout(\nx.n1998 ),
            .ltout(),
            .carryin(\nx.n10652 ),
            .carryout(\nx.n10653 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_14_lut_LC_7_26_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_14_lut_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_14_lut_LC_7_26_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_14_lut_LC_7_26_4  (
            .in0(N__32364),
            .in1(N__32363),
            .in2(N__30781),
            .in3(N__30795),
            .lcout(\nx.n1997 ),
            .ltout(),
            .carryin(\nx.n10653 ),
            .carryout(\nx.n10654 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_15_lut_LC_7_26_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_15_lut_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_15_lut_LC_7_26_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_15_lut_LC_7_26_5  (
            .in0(N__30686),
            .in1(N__30685),
            .in2(N__30785),
            .in3(N__30792),
            .lcout(\nx.n1996 ),
            .ltout(),
            .carryin(\nx.n10654 ),
            .carryout(\nx.n10655 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_16_lut_LC_7_26_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_16_lut_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_16_lut_LC_7_26_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_16_lut_LC_7_26_6  (
            .in0(N__32793),
            .in1(N__32792),
            .in2(N__30782),
            .in3(N__30789),
            .lcout(\nx.n1995 ),
            .ltout(),
            .carryin(\nx.n10655 ),
            .carryout(\nx.n10656 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_17_lut_LC_7_26_7 .C_ON=1'b0;
    defparam \nx.mod_5_add_1339_17_lut_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_17_lut_LC_7_26_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1339_17_lut_LC_7_26_7  (
            .in0(N__32819),
            .in1(N__32820),
            .in2(N__30786),
            .in3(N__30690),
            .lcout(\nx.n1994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1220_3_lut_LC_7_27_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1220_3_lut_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1220_3_lut_LC_7_27_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1220_3_lut_LC_7_27_0  (
            .in0(N__34932),
            .in1(N__34976),
            .in2(_gnd_net_),
            .in3(N__35149),
            .lcout(\nx.n1809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_3_lut_LC_7_27_1 .C_ON=1'b0;
    defparam \nx.i4_3_lut_LC_7_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.i4_3_lut_LC_7_27_1 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \nx.i4_3_lut_LC_7_27_1  (
            .in0(_gnd_net_),
            .in1(N__41279),
            .in2(N__41208),
            .in3(N__41883),
            .lcout(\nx.n24_adj_654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1216_3_lut_LC_7_27_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1216_3_lut_LC_7_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1216_3_lut_LC_7_27_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1216_3_lut_LC_7_27_2  (
            .in0(N__34764),
            .in1(N__34780),
            .in2(_gnd_net_),
            .in3(N__35150),
            .lcout(\nx.n1805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1276_3_lut_LC_7_27_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1276_3_lut_LC_7_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1276_3_lut_LC_7_27_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1276_3_lut_LC_7_27_4  (
            .in0(_gnd_net_),
            .in1(N__34578),
            .in2(N__32901),
            .in3(N__32955),
            .lcout(\nx.n1897 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1281_3_lut_LC_7_27_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1281_3_lut_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1281_3_lut_LC_7_27_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.mod_5_i1281_3_lut_LC_7_27_6  (
            .in0(N__32883),
            .in1(N__33087),
            .in2(N__34617),
            .in3(_gnd_net_),
            .lcout(\nx.n1902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9576_1_lut_LC_7_28_0 .C_ON=1'b0;
    defparam \nx.i9576_1_lut_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.i9576_1_lut_LC_7_28_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.i9576_1_lut_LC_7_28_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30644),
            .lcout(\nx.n13425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1144_3_lut_LC_7_28_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1144_3_lut_LC_7_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1144_3_lut_LC_7_28_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1144_3_lut_LC_7_28_1  (
            .in0(_gnd_net_),
            .in1(N__34482),
            .in2(N__31160),
            .in3(N__31131),
            .lcout(\nx.n1701 ),
            .ltout(\nx.n1701_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1211_3_lut_LC_7_28_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1211_3_lut_LC_7_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1211_3_lut_LC_7_28_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1211_3_lut_LC_7_28_2  (
            .in0(N__35298),
            .in1(_gnd_net_),
            .in2(N__30867),
            .in3(N__35146),
            .lcout(\nx.n1800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1212_3_lut_LC_7_28_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1212_3_lut_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1212_3_lut_LC_7_28_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1212_3_lut_LC_7_28_4  (
            .in0(_gnd_net_),
            .in1(N__35357),
            .in2(N__35343),
            .in3(N__35147),
            .lcout(\nx.n1801 ),
            .ltout(\nx.n1801_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_133_LC_7_28_5 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_133_LC_7_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_133_LC_7_28_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_adj_133_LC_7_28_5  (
            .in0(N__33016),
            .in1(N__35006),
            .in2(N__30864),
            .in3(N__34434),
            .lcout(\nx.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_3_lut_adj_82_LC_7_28_6 .C_ON=1'b0;
    defparam \nx.i3_3_lut_adj_82_LC_7_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.i3_3_lut_adj_82_LC_7_28_6 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \nx.i3_3_lut_adj_82_LC_7_28_6  (
            .in0(_gnd_net_),
            .in1(N__34965),
            .in2(N__34912),
            .in3(N__35356),
            .lcout(\nx.n16_adj_672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1149_3_lut_LC_7_28_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1149_3_lut_LC_7_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1149_3_lut_LC_7_28_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1149_3_lut_LC_7_28_7  (
            .in0(_gnd_net_),
            .in1(N__30891),
            .in2(N__30915),
            .in3(N__34481),
            .lcout(\nx.n1706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i7_LC_7_29_0.C_ON=1'b0;
    defparam neopxl_color_i7_LC_7_29_0.SEQ_MODE=4'b1001;
    defparam neopxl_color_i7_LC_7_29_0.LUT_INIT=16'b0000111100001000;
    LogicCell40 neopxl_color_i7_LC_7_29_0 (
            .in0(N__50076),
            .in1(N__49850),
            .in2(N__49601),
            .in3(N__37395),
            .lcout(neopxl_color_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48443),
            .ce(),
            .sr(N__37371));
    defparam \nx.mod_5_i1084_3_lut_LC_7_29_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1084_3_lut_LC_7_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1084_3_lut_LC_7_29_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1084_3_lut_LC_7_29_1  (
            .in0(_gnd_net_),
            .in1(N__30855),
            .in2(N__33273),
            .in3(N__30844),
            .lcout(\nx.n1609 ),
            .ltout(\nx.n1609_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_3_lut_adj_89_LC_7_29_2 .C_ON=1'b0;
    defparam \nx.i4_3_lut_adj_89_LC_7_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.i4_3_lut_adj_89_LC_7_29_2 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \nx.i4_3_lut_adj_89_LC_7_29_2  (
            .in0(_gnd_net_),
            .in1(N__31186),
            .in2(N__30804),
            .in3(N__30999),
            .lcout(\nx.n16_adj_646 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1151_3_lut_LC_7_29_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1151_3_lut_LC_7_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1151_3_lut_LC_7_29_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1151_3_lut_LC_7_29_4  (
            .in0(N__30927),
            .in1(_gnd_net_),
            .in2(N__34500),
            .in3(N__30941),
            .lcout(\nx.n1708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1145_3_lut_LC_7_29_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1145_3_lut_LC_7_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1145_3_lut_LC_7_29_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1145_3_lut_LC_7_29_5  (
            .in0(N__31187),
            .in1(_gnd_net_),
            .in2(N__31173),
            .in3(N__34476),
            .lcout(\nx.n1702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1077_3_lut_LC_7_29_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1077_3_lut_LC_7_29_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1077_3_lut_LC_7_29_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1077_3_lut_LC_7_29_7  (
            .in0(_gnd_net_),
            .in1(N__31041),
            .in2(N__33274),
            .in3(N__31031),
            .lcout(\nx.n1602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_2_lut_LC_7_30_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_2_lut_LC_7_30_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_2_lut_LC_7_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_2_lut_LC_7_30_0  (
            .in0(_gnd_net_),
            .in1(N__31004),
            .in2(_gnd_net_),
            .in3(N__30945),
            .lcout(\nx.n1677 ),
            .ltout(),
            .carryin(bfn_7_30_0_),
            .carryout(\nx.n10603 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_3_lut_LC_7_30_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_3_lut_LC_7_30_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_3_lut_LC_7_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_3_lut_LC_7_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30942),
            .in3(N__30921),
            .lcout(\nx.n1676 ),
            .ltout(),
            .carryin(\nx.n10603 ),
            .carryout(\nx.n10604 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_4_lut_LC_7_30_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_4_lut_LC_7_30_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_4_lut_LC_7_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_4_lut_LC_7_30_2  (
            .in0(_gnd_net_),
            .in1(N__44932),
            .in2(N__34554),
            .in3(N__30918),
            .lcout(\nx.n1675 ),
            .ltout(),
            .carryin(\nx.n10604 ),
            .carryout(\nx.n10605 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_5_lut_LC_7_30_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_5_lut_LC_7_30_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_5_lut_LC_7_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_5_lut_LC_7_30_3  (
            .in0(_gnd_net_),
            .in1(N__44935),
            .in2(N__30914),
            .in3(N__30882),
            .lcout(\nx.n1674 ),
            .ltout(),
            .carryin(\nx.n10605 ),
            .carryout(\nx.n10606 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_6_lut_LC_7_30_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_6_lut_LC_7_30_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_6_lut_LC_7_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_6_lut_LC_7_30_4  (
            .in0(_gnd_net_),
            .in1(N__44933),
            .in2(N__33137),
            .in3(N__30879),
            .lcout(\nx.n1673 ),
            .ltout(),
            .carryin(\nx.n10606 ),
            .carryout(\nx.n10607 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_7_lut_LC_7_30_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_7_lut_LC_7_30_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_7_lut_LC_7_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_7_lut_LC_7_30_5  (
            .in0(_gnd_net_),
            .in1(N__44936),
            .in2(N__33207),
            .in3(N__30870),
            .lcout(\nx.n1672 ),
            .ltout(),
            .carryin(\nx.n10607 ),
            .carryout(\nx.n10608 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_8_lut_LC_7_30_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_8_lut_LC_7_30_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_8_lut_LC_7_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_8_lut_LC_7_30_6  (
            .in0(_gnd_net_),
            .in1(N__44934),
            .in2(N__33176),
            .in3(N__31194),
            .lcout(\nx.n1671 ),
            .ltout(),
            .carryin(\nx.n10608 ),
            .carryout(\nx.n10609 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_9_lut_LC_7_30_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_9_lut_LC_7_30_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_9_lut_LC_7_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_9_lut_LC_7_30_7  (
            .in0(_gnd_net_),
            .in1(N__44937),
            .in2(N__31191),
            .in3(N__31164),
            .lcout(\nx.n1670 ),
            .ltout(),
            .carryin(\nx.n10609 ),
            .carryout(\nx.n10610 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_10_lut_LC_7_31_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_10_lut_LC_7_31_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_10_lut_LC_7_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_10_lut_LC_7_31_0  (
            .in0(_gnd_net_),
            .in1(N__44518),
            .in2(N__31161),
            .in3(N__31122),
            .lcout(\nx.n1669 ),
            .ltout(),
            .carryin(bfn_7_31_0_),
            .carryout(\nx.n10611 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_11_lut_LC_7_31_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_11_lut_LC_7_31_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_11_lut_LC_7_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_11_lut_LC_7_31_1  (
            .in0(_gnd_net_),
            .in1(N__44520),
            .in2(N__33392),
            .in3(N__31119),
            .lcout(\nx.n1668 ),
            .ltout(),
            .carryin(\nx.n10611 ),
            .carryout(\nx.n10612 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_12_lut_LC_7_31_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_12_lut_LC_7_31_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_12_lut_LC_7_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_12_lut_LC_7_31_2  (
            .in0(_gnd_net_),
            .in1(N__44519),
            .in2(N__31071),
            .in3(N__31116),
            .lcout(\nx.n1667 ),
            .ltout(),
            .carryin(\nx.n10612 ),
            .carryout(\nx.n10613 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_13_lut_LC_7_31_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_13_lut_LC_7_31_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_13_lut_LC_7_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1138_13_lut_LC_7_31_3  (
            .in0(_gnd_net_),
            .in1(N__44521),
            .in2(N__31113),
            .in3(N__31092),
            .lcout(\nx.n1666 ),
            .ltout(),
            .carryin(\nx.n10613 ),
            .carryout(\nx.n10614 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_14_lut_LC_7_31_4 .C_ON=1'b0;
    defparam \nx.mod_5_add_1138_14_lut_LC_7_31_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_14_lut_LC_7_31_4 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1138_14_lut_LC_7_31_4  (
            .in0(N__44522),
            .in1(N__31088),
            .in2(N__34515),
            .in3(N__31074),
            .lcout(\nx.n1697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1142_3_lut_LC_7_31_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1142_3_lut_LC_7_31_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1142_3_lut_LC_7_31_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1142_3_lut_LC_7_31_5  (
            .in0(_gnd_net_),
            .in1(N__31069),
            .in2(N__31050),
            .in3(N__34504),
            .lcout(\nx.n1699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_210_LC_9_15_5.C_ON=1'b0;
    defparam i1_4_lut_adj_210_LC_9_15_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_210_LC_9_15_5.LUT_INIT=16'b0000101000101010;
    LogicCell40 i1_4_lut_adj_210_LC_9_15_5 (
            .in0(N__47504),
            .in1(N__47995),
            .in2(N__37584),
            .in3(N__35502),
            .lcout(),
            .ltout(n7258_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i2_LC_9_15_6.C_ON=1'b0;
    defparam pin_output_i0_i2_LC_9_15_6.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i2_LC_9_15_6.LUT_INIT=16'b0000110010101100;
    LogicCell40 pin_output_i0_i2_LC_9_15_6 (
            .in0(N__37583),
            .in1(N__31360),
            .in2(N__31257),
            .in3(N__46534),
            .lcout(pin_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48417),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_202_LC_9_16_0.C_ON=1'b0;
    defparam i1_4_lut_adj_202_LC_9_16_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_202_LC_9_16_0.LUT_INIT=16'b0010001000101010;
    LogicCell40 i1_4_lut_adj_202_LC_9_16_0 (
            .in0(N__47502),
            .in1(N__35471),
            .in2(N__42645),
            .in3(N__35504),
            .lcout(n7236),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_159_LC_9_16_5.C_ON=1'b0;
    defparam i1_4_lut_adj_159_LC_9_16_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_159_LC_9_16_5.LUT_INIT=16'b0100010001001100;
    LogicCell40 i1_4_lut_adj_159_LC_9_16_5 (
            .in0(N__35525),
            .in1(N__47503),
            .in2(N__42702),
            .in3(N__37493),
            .lcout(),
            .ltout(n7270_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i5_LC_9_16_6.C_ON=1'b0;
    defparam pin_output_i0_i5_LC_9_16_6.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i5_LC_9_16_6.LUT_INIT=16'b0000110010101100;
    LogicCell40 pin_output_i0_i5_LC_9_16_6 (
            .in0(N__35526),
            .in1(N__31214),
            .in2(N__31245),
            .in3(N__46519),
            .lcout(pin_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48412),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_206_LC_9_16_7.C_ON=1'b0;
    defparam i1_4_lut_adj_206_LC_9_16_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_206_LC_9_16_7.LUT_INIT=16'b0000010011001100;
    LogicCell40 i1_4_lut_adj_206_LC_9_16_7 (
            .in0(N__35503),
            .in1(N__47501),
            .in2(N__42701),
            .in3(N__33098),
            .lcout(n7254),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_232_LC_9_17_0.C_ON=1'b0;
    defparam i1_2_lut_adj_232_LC_9_17_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_232_LC_9_17_0.LUT_INIT=16'b1010111110101111;
    LogicCell40 i1_2_lut_adj_232_LC_9_17_0 (
            .in0(N__50328),
            .in1(_gnd_net_),
            .in2(N__49050),
            .in3(_gnd_net_),
            .lcout(n6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9305_3_lut_LC_9_17_2.C_ON=1'b0;
    defparam i9305_3_lut_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam i9305_3_lut_LC_9_17_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 i9305_3_lut_LC_9_17_2 (
            .in0(N__49043),
            .in1(N__31213),
            .in2(_gnd_net_),
            .in3(N__35951),
            .lcout(),
            .ltout(n13152_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_1__bdd_4_lut_9614_LC_9_17_3.C_ON=1'b0;
    defparam current_pin_1__bdd_4_lut_9614_LC_9_17_3.SEQ_MODE=4'b0000;
    defparam current_pin_1__bdd_4_lut_9614_LC_9_17_3.LUT_INIT=16'b1110110001100100;
    LogicCell40 current_pin_1__bdd_4_lut_9614_LC_9_17_3 (
            .in0(N__50562),
            .in1(N__50327),
            .in2(N__31197),
            .in3(N__31407),
            .lcout(),
            .ltout(n13462_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13462_bdd_4_lut_LC_9_17_4.C_ON=1'b0;
    defparam n13462_bdd_4_lut_LC_9_17_4.SEQ_MODE=4'b0000;
    defparam n13462_bdd_4_lut_LC_9_17_4.LUT_INIT=16'b1111001011000010;
    LogicCell40 n13462_bdd_4_lut_LC_9_17_4 (
            .in0(N__31422),
            .in1(N__50563),
            .in2(N__31410),
            .in3(N__31341),
            .lcout(n13465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9321_3_lut_LC_9_17_5.C_ON=1'b0;
    defparam i9321_3_lut_LC_9_17_5.SEQ_MODE=4'b0000;
    defparam i9321_3_lut_LC_9_17_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 i9321_3_lut_LC_9_17_5 (
            .in0(N__40478),
            .in1(N__49044),
            .in2(_gnd_net_),
            .in3(N__40544),
            .lcout(n13168),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9306_3_lut_LC_9_17_6.C_ON=1'b0;
    defparam i9306_3_lut_LC_9_17_6.SEQ_MODE=4'b0000;
    defparam i9306_3_lut_LC_9_17_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 i9306_3_lut_LC_9_17_6 (
            .in0(N__49042),
            .in1(N__33502),
            .in2(_gnd_net_),
            .in3(N__33541),
            .lcout(n13153),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i3_LC_9_18_0.C_ON=1'b0;
    defparam pin_output_i0_i3_LC_9_18_0.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i3_LC_9_18_0.LUT_INIT=16'b0100010011100100;
    LogicCell40 pin_output_i0_i3_LC_9_18_0 (
            .in0(N__33525),
            .in1(N__31388),
            .in2(N__37521),
            .in3(N__46530),
            .lcout(pin_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48413),
            .ce(),
            .sr(_gnd_net_));
    defparam i9300_3_lut_LC_9_18_3.C_ON=1'b0;
    defparam i9300_3_lut_LC_9_18_3.SEQ_MODE=4'b0000;
    defparam i9300_3_lut_LC_9_18_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i9300_3_lut_LC_9_18_3 (
            .in0(N__31387),
            .in1(N__31361),
            .in2(_gnd_net_),
            .in3(N__49030),
            .lcout(n13147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9320_3_lut_LC_9_18_5.C_ON=1'b0;
    defparam i9320_3_lut_LC_9_18_5.SEQ_MODE=4'b0000;
    defparam i9320_3_lut_LC_9_18_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 i9320_3_lut_LC_9_18_5 (
            .in0(N__40517),
            .in1(N__39221),
            .in2(_gnd_net_),
            .in3(N__49031),
            .lcout(),
            .ltout(n13167_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13450_bdd_4_lut_LC_9_18_6.C_ON=1'b0;
    defparam n13450_bdd_4_lut_LC_9_18_6.SEQ_MODE=4'b0000;
    defparam n13450_bdd_4_lut_LC_9_18_6.LUT_INIT=16'b1110111000110000;
    LogicCell40 n13450_bdd_4_lut_LC_9_18_6 (
            .in0(N__31335),
            .in1(N__50568),
            .in2(N__31329),
            .in3(N__31326),
            .lcout(n13453),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1817_3_lut_LC_9_19_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1817_3_lut_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1817_3_lut_LC_9_19_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1817_3_lut_LC_9_19_0  (
            .in0(N__33699),
            .in1(_gnd_net_),
            .in2(N__36194),
            .in3(N__33719),
            .lcout(\nx.n2694 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1820_3_lut_LC_9_19_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1820_3_lut_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1820_3_lut_LC_9_19_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1820_3_lut_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__36306),
            .in2(N__33765),
            .in3(N__36158),
            .lcout(\nx.n2697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1827_3_lut_LC_9_19_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1827_3_lut_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1827_3_lut_LC_9_19_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1827_3_lut_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__37928),
            .in2(N__36191),
            .in3(N__33639),
            .lcout(\nx.n2704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1818_3_lut_LC_9_19_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1818_3_lut_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1818_3_lut_LC_9_19_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1818_3_lut_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__36387),
            .in2(N__33735),
            .in3(N__36151),
            .lcout(\nx.n2695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1821_3_lut_LC_9_19_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1821_3_lut_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1821_3_lut_LC_9_19_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1821_3_lut_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__36369),
            .in2(N__36193),
            .in3(N__33570),
            .lcout(\nx.n2698 ),
            .ltout(\nx.n2698_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_23_LC_9_19_5 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_23_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_23_LC_9_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_23_LC_9_19_5  (
            .in0(N__31585),
            .in1(N__36080),
            .in2(N__31494),
            .in3(N__31474),
            .lcout(\nx.n39_adj_610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1826_3_lut_LC_9_19_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1826_3_lut_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1826_3_lut_LC_9_19_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1826_3_lut_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__33627),
            .in2(N__36192),
            .in3(N__36339),
            .lcout(\nx.n2703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1832_3_lut_LC_9_19_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1832_3_lut_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1832_3_lut_LC_9_19_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i1832_3_lut_LC_9_19_7  (
            .in0(N__35907),
            .in1(N__33471),
            .in2(_gnd_net_),
            .in3(N__36144),
            .lcout(\nx.n2709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1696_3_lut_LC_9_20_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1696_3_lut_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1696_3_lut_LC_9_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1696_3_lut_LC_9_20_0  (
            .in0(N__41226),
            .in1(N__41275),
            .in2(_gnd_net_),
            .in3(N__41593),
            .lcout(\nx.n2509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1813_3_lut_LC_9_20_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1813_3_lut_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1813_3_lut_LC_9_20_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1813_3_lut_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__36411),
            .in2(N__36197),
            .in3(N__33660),
            .lcout(\nx.n2690 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1747_3_lut_LC_9_20_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1747_3_lut_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1747_3_lut_LC_9_20_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1747_3_lut_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__38295),
            .in2(N__39548),
            .in3(N__38271),
            .lcout(\nx.n2592 ),
            .ltout(\nx.n2592_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1814_3_lut_LC_9_20_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1814_3_lut_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1814_3_lut_LC_9_20_4 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.mod_5_i1814_3_lut_LC_9_20_4  (
            .in0(N__36166),
            .in1(N__33669),
            .in2(N__31425),
            .in3(_gnd_net_),
            .lcout(\nx.n2691 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1812_rep_23_3_lut_LC_9_20_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1812_rep_23_3_lut_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1812_rep_23_3_lut_LC_9_20_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1812_rep_23_3_lut_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__36170),
            .in2(N__36438),
            .in3(N__33651),
            .lcout(\nx.n2689 ),
            .ltout(\nx.n2689_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_20_LC_9_20_6 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_20_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_20_LC_9_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_20_LC_9_20_6  (
            .in0(N__31648),
            .in1(N__33884),
            .in2(N__31632),
            .in3(N__31610),
            .lcout(\nx.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1824_3_lut_LC_9_20_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1824_3_lut_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1824_3_lut_LC_9_20_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1824_3_lut_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__33600),
            .in2(N__36270),
            .in3(N__36171),
            .lcout(\nx.n2701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1419_3_lut_LC_9_21_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1419_3_lut_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1419_3_lut_LC_9_21_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1419_3_lut_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__32013),
            .in2(N__32049),
            .in3(N__34160),
            .lcout(\nx.n2104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1420_3_lut_LC_9_21_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1420_3_lut_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1420_3_lut_LC_9_21_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1420_3_lut_LC_9_21_1  (
            .in0(N__32061),
            .in1(_gnd_net_),
            .in2(N__34190),
            .in3(N__32097),
            .lcout(\nx.n2105 ),
            .ltout(\nx.n2105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_3_lut_LC_9_21_2 .C_ON=1'b0;
    defparam \nx.i9_3_lut_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9_3_lut_LC_9_21_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \nx.i9_3_lut_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__36737),
            .in2(N__31572),
            .in3(N__37316),
            .lcout(\nx.n26_adj_667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1410_3_lut_LC_9_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1410_3_lut_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1410_3_lut_LC_9_21_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1410_3_lut_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__32196),
            .in2(N__32157),
            .in3(N__34159),
            .lcout(\nx.n2095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1686_3_lut_LC_9_21_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1686_3_lut_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1686_3_lut_LC_9_21_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1686_3_lut_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__41385),
            .in2(N__43698),
            .in3(N__41612),
            .lcout(\nx.n2499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1750_3_lut_LC_9_21_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1750_3_lut_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1750_3_lut_LC_9_21_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1750_3_lut_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__37972),
            .in2(N__37947),
            .in3(N__39544),
            .lcout(\nx.n2595 ),
            .ltout(\nx.n2595_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_LC_9_21_7 .C_ON=1'b0;
    defparam \nx.i13_4_lut_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_LC_9_21_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_LC_9_21_7  (
            .in0(N__36009),
            .in1(N__36713),
            .in2(N__31950),
            .in3(N__33680),
            .lcout(\nx.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1418_3_lut_LC_9_22_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1418_3_lut_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1418_3_lut_LC_9_22_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1418_3_lut_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__31965),
            .in2(N__32001),
            .in3(N__34164),
            .lcout(\nx.n2103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_68_LC_9_22_1 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_68_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_68_LC_9_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_68_LC_9_22_1  (
            .in0(N__32332),
            .in1(N__32287),
            .in2(N__32247),
            .in3(N__34233),
            .lcout(),
            .ltout(\nx.n26_adj_664_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_71_LC_9_22_2 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_71_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_71_LC_9_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_71_LC_9_22_2  (
            .in0(N__31947),
            .in1(N__33990),
            .in2(N__31935),
            .in3(N__31932),
            .lcout(\nx.n2027 ),
            .ltout(\nx.n2027_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1413_3_lut_LC_9_22_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1413_3_lut_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1413_3_lut_LC_9_22_3 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \nx.mod_5_i1413_3_lut_LC_9_22_3  (
            .in0(N__32245),
            .in1(N__32214),
            .in2(N__31923),
            .in3(_gnd_net_),
            .lcout(\nx.n2098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1414_3_lut_LC_9_22_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1414_3_lut_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1414_3_lut_LC_9_22_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1414_3_lut_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__32259),
            .in2(N__32292),
            .in3(N__34168),
            .lcout(\nx.n2099 ),
            .ltout(\nx.n2099_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_73_LC_9_22_5 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_73_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_73_LC_9_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_73_LC_9_22_5  (
            .in0(N__37097),
            .in1(N__36976),
            .in2(N__31920),
            .in3(N__37027),
            .lcout(\nx.n28_adj_669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2030_3_lut_LC_9_22_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2030_3_lut_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2030_3_lut_LC_9_22_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2030_3_lut_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__31917),
            .in2(N__31890),
            .in3(N__31878),
            .lcout(\nx.n3003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1415_3_lut_LC_9_22_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1415_3_lut_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1415_3_lut_LC_9_22_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1415_3_lut_LC_9_22_7  (
            .in0(N__32333),
            .in1(_gnd_net_),
            .in2(N__34191),
            .in3(N__32304),
            .lcout(\nx.n2100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_2_lut_LC_9_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_2_lut_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_2_lut_LC_9_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_2_lut_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__34075),
            .in2(_gnd_net_),
            .in3(N__32109),
            .lcout(\nx.n2077 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\nx.n10657 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_3_lut_LC_9_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_3_lut_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_3_lut_LC_9_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_3_lut_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34016),
            .in3(N__32106),
            .lcout(\nx.n2076 ),
            .ltout(),
            .carryin(\nx.n10657 ),
            .carryout(\nx.n10658 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_4_lut_LC_9_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_4_lut_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_4_lut_LC_9_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_4_lut_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__44631),
            .in2(N__34290),
            .in3(N__32103),
            .lcout(\nx.n2075 ),
            .ltout(),
            .carryin(\nx.n10658 ),
            .carryout(\nx.n10659 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_5_lut_LC_9_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_5_lut_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_5_lut_LC_9_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_5_lut_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__44634),
            .in2(N__34691),
            .in3(N__32100),
            .lcout(\nx.n2074 ),
            .ltout(),
            .carryin(\nx.n10659 ),
            .carryout(\nx.n10660 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_6_lut_LC_9_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_6_lut_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_6_lut_LC_9_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_6_lut_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__44632),
            .in2(N__32096),
            .in3(N__32052),
            .lcout(\nx.n2073 ),
            .ltout(),
            .carryin(\nx.n10660 ),
            .carryout(\nx.n10661 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_7_lut_LC_9_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_7_lut_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_7_lut_LC_9_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_7_lut_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__44635),
            .in2(N__32048),
            .in3(N__32004),
            .lcout(\nx.n2072 ),
            .ltout(),
            .carryin(\nx.n10661 ),
            .carryout(\nx.n10662 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_8_lut_LC_9_23_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_8_lut_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_8_lut_LC_9_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_8_lut_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__44633),
            .in2(N__32000),
            .in3(N__31959),
            .lcout(\nx.n2071 ),
            .ltout(),
            .carryin(\nx.n10662 ),
            .carryout(\nx.n10663 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_9_lut_LC_9_23_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_9_lut_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_9_lut_LC_9_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_9_lut_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__44636),
            .in2(N__34041),
            .in3(N__31956),
            .lcout(\nx.n2070 ),
            .ltout(),
            .carryin(\nx.n10663 ),
            .carryout(\nx.n10664 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_10_lut_LC_9_24_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_10_lut_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_10_lut_LC_9_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_10_lut_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__45134),
            .in2(N__34658),
            .in3(N__31953),
            .lcout(\nx.n2069 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\nx.n10665 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_11_lut_LC_9_24_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_11_lut_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_11_lut_LC_9_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_11_lut_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__45138),
            .in2(N__32334),
            .in3(N__32295),
            .lcout(\nx.n2068 ),
            .ltout(),
            .carryin(\nx.n10665 ),
            .carryout(\nx.n10666 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_12_lut_LC_9_24_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_12_lut_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_12_lut_LC_9_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_12_lut_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__45135),
            .in2(N__32291),
            .in3(N__32250),
            .lcout(\nx.n2067 ),
            .ltout(),
            .carryin(\nx.n10666 ),
            .carryout(\nx.n10667 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_13_lut_LC_9_24_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_13_lut_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_13_lut_LC_9_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_13_lut_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__45139),
            .in2(N__32246),
            .in3(N__32205),
            .lcout(\nx.n2066 ),
            .ltout(),
            .carryin(\nx.n10667 ),
            .carryout(\nx.n10668 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_14_lut_LC_9_24_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_14_lut_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_14_lut_LC_9_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_14_lut_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(N__45136),
            .in2(N__34231),
            .in3(N__32202),
            .lcout(\nx.n2065 ),
            .ltout(),
            .carryin(\nx.n10668 ),
            .carryout(\nx.n10669 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_15_lut_LC_9_24_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_15_lut_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_15_lut_LC_9_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_15_lut_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(N__45140),
            .in2(N__34388),
            .in3(N__32199),
            .lcout(\nx.n2064 ),
            .ltout(),
            .carryin(\nx.n10669 ),
            .carryout(\nx.n10670 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_16_lut_LC_9_24_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_16_lut_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_16_lut_LC_9_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_16_lut_LC_9_24_6  (
            .in0(_gnd_net_),
            .in1(N__45137),
            .in2(N__32195),
            .in3(N__32142),
            .lcout(\nx.n2063 ),
            .ltout(),
            .carryin(\nx.n10670 ),
            .carryout(\nx.n10671 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_17_lut_LC_9_24_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_17_lut_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_17_lut_LC_9_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_17_lut_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(N__45141),
            .in2(N__34346),
            .in3(N__32139),
            .lcout(\nx.n2062 ),
            .ltout(),
            .carryin(\nx.n10671 ),
            .carryout(\nx.n10672 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_18_lut_LC_9_25_0 .C_ON=1'b0;
    defparam \nx.mod_5_add_1406_18_lut_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_18_lut_LC_9_25_0 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_1406_18_lut_LC_9_25_0  (
            .in0(N__44630),
            .in1(N__34192),
            .in2(N__32136),
            .in3(N__32112),
            .lcout(\nx.n2093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1280_3_lut_LC_9_25_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1280_3_lut_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1280_3_lut_LC_9_25_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1280_3_lut_LC_9_25_2  (
            .in0(N__33075),
            .in1(_gnd_net_),
            .in2(N__35007),
            .in3(N__32903),
            .lcout(\nx.n1901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9518_3_lut_LC_9_25_4 .C_ON=1'b0;
    defparam \nx.i9518_3_lut_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.i9518_3_lut_LC_9_25_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.i9518_3_lut_LC_9_25_4  (
            .in0(_gnd_net_),
            .in1(N__34433),
            .in2(N__32553),
            .in3(N__32902),
            .lcout(\nx.n1905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_LC_9_25_5 .C_ON=1'b0;
    defparam \nx.i10_4_lut_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_LC_9_25_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_LC_9_25_5  (
            .in0(N__32422),
            .in1(N__32380),
            .in2(N__32791),
            .in3(N__32812),
            .lcout(\nx.n25_adj_606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8_4_lut_adj_155_LC_9_26_0 .C_ON=1'b0;
    defparam \nx.i8_4_lut_adj_155_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.i8_4_lut_adj_155_LC_9_26_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i8_4_lut_adj_155_LC_9_26_0  (
            .in0(N__32978),
            .in1(N__34570),
            .in2(N__35049),
            .in3(N__32933),
            .lcout(\nx.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1279_3_lut_LC_9_26_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1279_3_lut_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1279_3_lut_LC_9_26_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1279_3_lut_LC_9_26_1  (
            .in0(_gnd_net_),
            .in1(N__33063),
            .in2(N__33039),
            .in3(N__32896),
            .lcout(\nx.n1900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1210_3_lut_LC_9_26_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1210_3_lut_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1210_3_lut_LC_9_26_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1210_3_lut_LC_9_26_2  (
            .in0(N__35262),
            .in1(N__35283),
            .in2(_gnd_net_),
            .in3(N__35125),
            .lcout(\nx.n1799 ),
            .ltout(\nx.n1799_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1277_3_lut_LC_9_26_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1277_3_lut_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1277_3_lut_LC_9_26_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1277_3_lut_LC_9_26_3  (
            .in0(_gnd_net_),
            .in1(N__32967),
            .in2(N__32367),
            .in3(N__32898),
            .lcout(\nx.n1898 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1218_3_lut_LC_9_26_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1218_3_lut_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1218_3_lut_LC_9_26_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i1218_3_lut_LC_9_26_5  (
            .in0(N__35127),
            .in1(_gnd_net_),
            .in2(N__34869),
            .in3(N__34830),
            .lcout(\nx.n1807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1208_3_lut_LC_9_26_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1208_3_lut_LC_9_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1208_3_lut_LC_9_26_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1208_3_lut_LC_9_26_6  (
            .in0(_gnd_net_),
            .in1(N__35205),
            .in2(N__35169),
            .in3(N__35126),
            .lcout(\nx.n1797 ),
            .ltout(\nx.n1797_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1275_3_lut_LC_9_26_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1275_3_lut_LC_9_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1275_3_lut_LC_9_26_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1275_3_lut_LC_9_26_7  (
            .in0(_gnd_net_),
            .in1(N__32897),
            .in2(N__32337),
            .in3(N__32922),
            .lcout(\nx.n1896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2_2_lut_adj_134_LC_9_27_0 .C_ON=1'b1;
    defparam \nx.i2_2_lut_adj_134_LC_9_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.i2_2_lut_adj_134_LC_9_27_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \nx.i2_2_lut_adj_134_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__32765),
            .in2(_gnd_net_),
            .in3(N__32721),
            .lcout(\nx.n30_adj_703 ),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\nx.n10628 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_3_lut_LC_9_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_3_lut_LC_9_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_3_lut_LC_9_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_3_lut_LC_9_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32667),
            .in3(N__32631),
            .lcout(\nx.n1876 ),
            .ltout(),
            .carryin(\nx.n10628 ),
            .carryout(\nx.n10629 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_4_lut_LC_9_27_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_4_lut_LC_9_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_4_lut_LC_9_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_4_lut_LC_9_27_2  (
            .in0(_gnd_net_),
            .in1(N__44956),
            .in2(N__32628),
            .in3(N__32595),
            .lcout(\nx.n1875 ),
            .ltout(),
            .carryin(\nx.n10629 ),
            .carryout(\nx.n10630 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_5_lut_LC_9_27_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_5_lut_LC_9_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_5_lut_LC_9_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_5_lut_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(N__45296),
            .in2(N__32587),
            .in3(N__32556),
            .lcout(\nx.n1874 ),
            .ltout(),
            .carryin(\nx.n10630 ),
            .carryout(\nx.n10631 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_6_lut_LC_9_27_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_6_lut_LC_9_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_6_lut_LC_9_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_6_lut_LC_9_27_4  (
            .in0(_gnd_net_),
            .in1(N__44957),
            .in2(N__34432),
            .in3(N__32541),
            .lcout(\nx.n1873 ),
            .ltout(),
            .carryin(\nx.n10631 ),
            .carryout(\nx.n10632 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_7_lut_LC_9_27_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_7_lut_LC_9_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_7_lut_LC_9_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_7_lut_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(N__45297),
            .in2(N__32537),
            .in3(N__32493),
            .lcout(\nx.n1872 ),
            .ltout(),
            .carryin(\nx.n10632 ),
            .carryout(\nx.n10633 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_8_lut_LC_9_27_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_8_lut_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_8_lut_LC_9_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_8_lut_LC_9_27_6  (
            .in0(_gnd_net_),
            .in1(N__44958),
            .in2(N__32490),
            .in3(N__32460),
            .lcout(\nx.n1871 ),
            .ltout(),
            .carryin(\nx.n10633 ),
            .carryout(\nx.n10634 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_9_lut_LC_9_27_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_9_lut_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_9_lut_LC_9_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_9_lut_LC_9_27_7  (
            .in0(_gnd_net_),
            .in1(N__34612),
            .in2(N__45391),
            .in3(N__33078),
            .lcout(\nx.n1870 ),
            .ltout(),
            .carryin(\nx.n10634 ),
            .carryout(\nx.n10635 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_10_lut_LC_9_28_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_10_lut_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_10_lut_LC_9_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_10_lut_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(N__44717),
            .in2(N__35005),
            .in3(N__33066),
            .lcout(\nx.n1869 ),
            .ltout(),
            .carryin(bfn_9_28_0_),
            .carryout(\nx.n10636 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_11_lut_LC_9_28_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_11_lut_LC_9_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_11_lut_LC_9_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_11_lut_LC_9_28_1  (
            .in0(_gnd_net_),
            .in1(N__45096),
            .in2(N__33062),
            .in3(N__33027),
            .lcout(\nx.n1868 ),
            .ltout(),
            .carryin(\nx.n10636 ),
            .carryout(\nx.n10637 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_12_lut_LC_9_28_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_12_lut_LC_9_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_12_lut_LC_9_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_12_lut_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(N__44718),
            .in2(N__33024),
            .in3(N__32985),
            .lcout(\nx.n1867 ),
            .ltout(),
            .carryin(\nx.n10637 ),
            .carryout(\nx.n10638 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_13_lut_LC_9_28_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_13_lut_LC_9_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_13_lut_LC_9_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_13_lut_LC_9_28_3  (
            .in0(_gnd_net_),
            .in1(N__32982),
            .in2(N__45095),
            .in3(N__32958),
            .lcout(\nx.n1866 ),
            .ltout(),
            .carryin(\nx.n10638 ),
            .carryout(\nx.n10639 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_14_lut_LC_9_28_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_14_lut_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_14_lut_LC_9_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_14_lut_LC_9_28_4  (
            .in0(_gnd_net_),
            .in1(N__44722),
            .in2(N__34577),
            .in3(N__32943),
            .lcout(\nx.n1865 ),
            .ltout(),
            .carryin(\nx.n10639 ),
            .carryout(\nx.n10640 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_15_lut_LC_9_28_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_15_lut_LC_9_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_15_lut_LC_9_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1272_15_lut_LC_9_28_5  (
            .in0(_gnd_net_),
            .in1(N__45097),
            .in2(N__32940),
            .in3(N__32913),
            .lcout(\nx.n1864 ),
            .ltout(),
            .carryin(\nx.n10640 ),
            .carryout(\nx.n10641 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_16_lut_LC_9_28_6 .C_ON=1'b0;
    defparam \nx.mod_5_add_1272_16_lut_LC_9_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_16_lut_LC_9_28_6 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1272_16_lut_LC_9_28_6  (
            .in0(N__45098),
            .in1(N__35045),
            .in2(N__32910),
            .in3(N__32823),
            .lcout(\nx.n1895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1143_3_lut_LC_9_28_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1143_3_lut_LC_9_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1143_3_lut_LC_9_28_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1143_3_lut_LC_9_28_7  (
            .in0(_gnd_net_),
            .in1(N__33411),
            .in2(N__33399),
            .in3(N__34518),
            .lcout(\nx.n1700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i4_LC_9_29_0.C_ON=1'b0;
    defparam neopxl_color_i4_LC_9_29_0.SEQ_MODE=4'b1001;
    defparam neopxl_color_i4_LC_9_29_0.LUT_INIT=16'b0000111100001000;
    LogicCell40 neopxl_color_i4_LC_9_29_0 (
            .in0(N__49829),
            .in1(N__50078),
            .in2(N__49602),
            .in3(N__40864),
            .lcout(neopxl_color_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48446),
            .ce(),
            .sr(N__40842));
    defparam \nx.mod_5_i1083_3_lut_LC_9_29_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1083_3_lut_LC_9_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1083_3_lut_LC_9_29_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1083_3_lut_LC_9_29_2  (
            .in0(_gnd_net_),
            .in1(N__33369),
            .in2(N__33339),
            .in3(N__33270),
            .lcout(\nx.n1608 ),
            .ltout(\nx.n1608_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_2_lut_LC_9_29_3 .C_ON=1'b0;
    defparam \nx.i6_2_lut_LC_9_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.i6_2_lut_LC_9_29_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i6_2_lut_LC_9_29_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33324),
            .in3(N__33196),
            .lcout(\nx.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1080_3_lut_LC_9_29_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1080_3_lut_LC_9_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1080_3_lut_LC_9_29_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1080_3_lut_LC_9_29_4  (
            .in0(_gnd_net_),
            .in1(N__33312),
            .in2(N__33291),
            .in3(N__33271),
            .lcout(\nx.n1605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1146_3_lut_LC_9_29_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1146_3_lut_LC_9_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1146_3_lut_LC_9_29_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1146_3_lut_LC_9_29_5  (
            .in0(_gnd_net_),
            .in1(N__33177),
            .in2(N__33153),
            .in3(N__34511),
            .lcout(\nx.n1703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1148_3_lut_LC_9_29_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1148_3_lut_LC_9_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1148_3_lut_LC_9_29_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1148_3_lut_LC_9_29_6  (
            .in0(N__33138),
            .in1(_gnd_net_),
            .in2(N__34517),
            .in3(N__33120),
            .lcout(\nx.n1705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_1096_i21_2_lut_LC_10_15_0.C_ON=1'b0;
    defparam equal_1096_i21_2_lut_LC_10_15_0.SEQ_MODE=4'b0000;
    defparam equal_1096_i21_2_lut_LC_10_15_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 equal_1096_i21_2_lut_LC_10_15_0 (
            .in0(_gnd_net_),
            .in1(N__50554),
            .in2(_gnd_net_),
            .in3(N__50357),
            .lcout(n21),
            .ltout(n21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2930_3_lut_4_lut_LC_10_15_1.C_ON=1'b0;
    defparam i2930_3_lut_4_lut_LC_10_15_1.SEQ_MODE=4'b0000;
    defparam i2930_3_lut_4_lut_LC_10_15_1.LUT_INIT=16'b1100110011001000;
    LogicCell40 i2930_3_lut_4_lut_LC_10_15_1 (
            .in0(N__40441),
            .in1(N__46965),
            .in2(N__33108),
            .in3(N__40352),
            .lcout(n6150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i6_LC_10_16_0.C_ON=1'b0;
    defparam pin_output_i0_i6_LC_10_16_0.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i6_LC_10_16_0.LUT_INIT=16'b0111001001010000;
    LogicCell40 pin_output_i0_i6_LC_10_16_0 (
            .in0(N__33477),
            .in1(N__46523),
            .in2(N__33548),
            .in3(N__33486),
            .lcout(pin_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48415),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_213_LC_10_16_2.C_ON=1'b0;
    defparam i1_4_lut_adj_213_LC_10_16_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_213_LC_10_16_2.LUT_INIT=16'b0100110001000100;
    LogicCell40 i1_4_lut_adj_213_LC_10_16_2 (
            .in0(N__37517),
            .in1(N__47495),
            .in2(N__35508),
            .in3(N__43293),
            .lcout(n7262),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i7_LC_10_16_4.C_ON=1'b0;
    defparam pin_output_i0_i7_LC_10_16_4.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i7_LC_10_16_4.LUT_INIT=16'b0101000011011000;
    LogicCell40 pin_output_i0_i7_LC_10_16_4 (
            .in0(N__35445),
            .in1(N__35454),
            .in2(N__33509),
            .in3(N__46524),
            .lcout(pin_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48415),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_10_16_6.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_10_16_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_10_16_6.LUT_INIT=16'b1111000011010000;
    LogicCell40 i1_3_lut_4_lut_LC_10_16_6 (
            .in0(N__50126),
            .in1(N__40444),
            .in2(N__46959),
            .in3(N__46683),
            .lcout(n8_adj_780),
            .ltout(n8_adj_780_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_161_LC_10_16_7.C_ON=1'b0;
    defparam i1_4_lut_adj_161_LC_10_16_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_161_LC_10_16_7.LUT_INIT=16'b0000101000101010;
    LogicCell40 i1_4_lut_adj_161_LC_10_16_7 (
            .in0(N__47496),
            .in1(N__37494),
            .in2(N__33480),
            .in3(N__47981),
            .lcout(n7274),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_2_lut_LC_10_17_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_2_lut_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_2_lut_LC_10_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_2_lut_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__35906),
            .in2(_gnd_net_),
            .in3(N__33462),
            .lcout(\nx.n2677 ),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\nx.n10768 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_3_lut_LC_10_17_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_3_lut_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_3_lut_LC_10_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_3_lut_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35924),
            .in3(N__33444),
            .lcout(\nx.n2676 ),
            .ltout(),
            .carryin(\nx.n10768 ),
            .carryout(\nx.n10769 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_4_lut_LC_10_17_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_4_lut_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_4_lut_LC_10_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_4_lut_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__45685),
            .in2(N__35825),
            .in3(N__33429),
            .lcout(\nx.n2675 ),
            .ltout(),
            .carryin(\nx.n10769 ),
            .carryout(\nx.n10770 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_5_lut_LC_10_17_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_5_lut_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_5_lut_LC_10_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_5_lut_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__45688),
            .in2(N__39422),
            .in3(N__33414),
            .lcout(\nx.n2674 ),
            .ltout(),
            .carryin(\nx.n10770 ),
            .carryout(\nx.n10771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_6_lut_LC_10_17_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_6_lut_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_6_lut_LC_10_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_6_lut_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__45686),
            .in2(N__36240),
            .in3(N__33642),
            .lcout(\nx.n2673 ),
            .ltout(),
            .carryin(\nx.n10771 ),
            .carryout(\nx.n10772 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_7_lut_LC_10_17_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_7_lut_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_7_lut_LC_10_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_7_lut_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__45689),
            .in2(N__37932),
            .in3(N__33630),
            .lcout(\nx.n2672 ),
            .ltout(),
            .carryin(\nx.n10772 ),
            .carryout(\nx.n10773 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_8_lut_LC_10_17_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_8_lut_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_8_lut_LC_10_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_8_lut_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__45687),
            .in2(N__36335),
            .in3(N__33618),
            .lcout(\nx.n2671 ),
            .ltout(),
            .carryin(\nx.n10773 ),
            .carryout(\nx.n10774 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_9_lut_LC_10_17_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_9_lut_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_9_lut_LC_10_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_9_lut_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__45690),
            .in2(N__36686),
            .in3(N__33603),
            .lcout(\nx.n2670 ),
            .ltout(),
            .carryin(\nx.n10774 ),
            .carryout(\nx.n10775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_10_lut_LC_10_18_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_10_lut_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_10_lut_LC_10_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_10_lut_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__45742),
            .in2(N__36263),
            .in3(N__33591),
            .lcout(\nx.n2669 ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\nx.n10776 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_11_lut_LC_10_18_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_11_lut_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_11_lut_LC_10_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_11_lut_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__45746),
            .in2(N__37667),
            .in3(N__33576),
            .lcout(\nx.n2668 ),
            .ltout(),
            .carryin(\nx.n10776 ),
            .carryout(\nx.n10777 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_12_lut_LC_10_18_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_12_lut_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_12_lut_LC_10_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_12_lut_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__45743),
            .in2(N__37617),
            .in3(N__33573),
            .lcout(\nx.n2667 ),
            .ltout(),
            .carryin(\nx.n10777 ),
            .carryout(\nx.n10778 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_13_lut_LC_10_18_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_13_lut_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_13_lut_LC_10_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_13_lut_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__45747),
            .in2(N__36365),
            .in3(N__33564),
            .lcout(\nx.n2666 ),
            .ltout(),
            .carryin(\nx.n10778 ),
            .carryout(\nx.n10779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_14_lut_LC_10_18_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_14_lut_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_14_lut_LC_10_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_14_lut_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(N__45744),
            .in2(N__36301),
            .in3(N__33756),
            .lcout(\nx.n2665 ),
            .ltout(),
            .carryin(\nx.n10779 ),
            .carryout(\nx.n10780 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_15_lut_LC_10_18_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_15_lut_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_15_lut_LC_10_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_15_lut_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__45748),
            .in2(N__37694),
            .in3(N__33738),
            .lcout(\nx.n2664 ),
            .ltout(),
            .carryin(\nx.n10780 ),
            .carryout(\nx.n10781 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_16_lut_LC_10_18_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_16_lut_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_16_lut_LC_10_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_16_lut_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__45745),
            .in2(N__36386),
            .in3(N__33726),
            .lcout(\nx.n2663 ),
            .ltout(),
            .carryin(\nx.n10781 ),
            .carryout(\nx.n10782 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_17_lut_LC_10_18_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_17_lut_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_17_lut_LC_10_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_17_lut_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__45749),
            .in2(N__33723),
            .in3(N__33693),
            .lcout(\nx.n2662 ),
            .ltout(),
            .carryin(\nx.n10782 ),
            .carryout(\nx.n10783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_18_lut_LC_10_19_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_18_lut_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_18_lut_LC_10_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_18_lut_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__45733),
            .in2(N__36008),
            .in3(N__33690),
            .lcout(\nx.n2661 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\nx.n10784 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_19_lut_LC_10_19_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_19_lut_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_19_lut_LC_10_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_19_lut_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__36714),
            .in2(N__45765),
            .in3(N__33687),
            .lcout(\nx.n2660 ),
            .ltout(),
            .carryin(\nx.n10784 ),
            .carryout(\nx.n10785 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_20_lut_LC_10_19_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_20_lut_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_20_lut_LC_10_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_20_lut_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__45737),
            .in2(N__33684),
            .in3(N__33663),
            .lcout(\nx.n2659 ),
            .ltout(),
            .carryin(\nx.n10785 ),
            .carryout(\nx.n10786 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_21_lut_LC_10_19_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_21_lut_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_21_lut_LC_10_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_21_lut_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__45739),
            .in2(N__36410),
            .in3(N__33654),
            .lcout(\nx.n2658 ),
            .ltout(),
            .carryin(\nx.n10786 ),
            .carryout(\nx.n10787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_22_lut_LC_10_19_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_22_lut_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_22_lut_LC_10_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_22_lut_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__45738),
            .in2(N__36434),
            .in3(N__33645),
            .lcout(\nx.n2657 ),
            .ltout(),
            .carryin(\nx.n10787 ),
            .carryout(\nx.n10788 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_23_lut_LC_10_19_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_23_lut_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_23_lut_LC_10_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_23_lut_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__45740),
            .in2(N__36657),
            .in3(N__33921),
            .lcout(\nx.n2656 ),
            .ltout(),
            .carryin(\nx.n10788 ),
            .carryout(\nx.n10789 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_24_lut_LC_10_19_6 .C_ON=1'b0;
    defparam \nx.mod_5_add_1808_24_lut_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_24_lut_LC_10_19_6 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1808_24_lut_LC_10_19_6  (
            .in0(N__45741),
            .in1(N__38169),
            .in2(N__36198),
            .in3(N__33918),
            .lcout(\nx.n2687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1815_3_lut_LC_10_20_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1815_3_lut_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1815_3_lut_LC_10_20_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1815_3_lut_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__36712),
            .in2(N__33915),
            .in3(N__36159),
            .lcout(\nx.n2692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_17_LC_10_20_1 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_17_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_17_LC_10_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_17_LC_10_20_1  (
            .in0(N__36427),
            .in1(N__36403),
            .in2(N__36656),
            .in3(N__38168),
            .lcout(),
            .ltout(\nx.n34_adj_603_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_3_lut_LC_10_20_2 .C_ON=1'b0;
    defparam \nx.i17_3_lut_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.i17_3_lut_LC_10_20_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \nx.i17_3_lut_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__37615),
            .in2(N__33873),
            .in3(N__36676),
            .lcout(),
            .ltout(\nx.n39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i21_4_lut_LC_10_20_3 .C_ON=1'b0;
    defparam \nx.i21_4_lut_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.i21_4_lut_LC_10_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i21_4_lut_LC_10_20_3  (
            .in0(N__36312),
            .in1(N__36276),
            .in2(N__33870),
            .in3(N__35835),
            .lcout(\nx.n2621 ),
            .ltout(\nx.n2621_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1816_3_lut_LC_10_20_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1816_3_lut_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1816_3_lut_LC_10_20_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1816_3_lut_LC_10_20_4  (
            .in0(N__36004),
            .in1(_gnd_net_),
            .in2(N__33867),
            .in3(N__33864),
            .lcout(\nx.n2693 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1822_3_lut_LC_10_20_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1822_3_lut_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1822_3_lut_LC_10_20_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1822_3_lut_LC_10_20_5  (
            .in0(N__37616),
            .in1(_gnd_net_),
            .in2(N__36196),
            .in3(N__33822),
            .lcout(\nx.n2699 ),
            .ltout(\nx.n2699_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_22_LC_10_20_6 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_22_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_22_LC_10_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_22_LC_10_20_6  (
            .in0(N__33779),
            .in1(N__36625),
            .in2(N__33768),
            .in3(N__33984),
            .lcout(\nx.n41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1811_3_lut_LC_10_20_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1811_3_lut_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1811_3_lut_LC_10_20_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1811_3_lut_LC_10_20_7  (
            .in0(N__36652),
            .in1(_gnd_net_),
            .in2(N__36195),
            .in3(N__33966),
            .lcout(\nx.n2688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1683_3_lut_LC_10_21_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1683_3_lut_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1683_3_lut_LC_10_21_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1683_3_lut_LC_10_21_0  (
            .in0(N__41316),
            .in1(_gnd_net_),
            .in2(N__41661),
            .in3(N__43200),
            .lcout(\nx.n2496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_59_LC_10_21_1 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_59_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_59_LC_10_21_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_59_LC_10_21_1  (
            .in0(N__41722),
            .in1(N__44010),
            .in2(N__41478),
            .in3(N__41764),
            .lcout(),
            .ltout(\nx.n31_adj_655_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_60_LC_10_21_2 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_60_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_60_LC_10_21_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_60_LC_10_21_2  (
            .in0(N__41804),
            .in1(N__41843),
            .in2(N__33960),
            .in3(N__33957),
            .lcout(),
            .ltout(\nx.n36_adj_656_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_65_LC_10_21_3 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_65_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_65_LC_10_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_65_LC_10_21_3  (
            .in0(N__43641),
            .in1(N__39702),
            .in2(N__33942),
            .in3(N__33939),
            .lcout(\nx.n2423 ),
            .ltout(\nx.n2423_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1677_3_lut_LC_10_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1677_3_lut_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1677_3_lut_LC_10_21_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1677_3_lut_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__41477),
            .in2(N__33927),
            .in3(N__41685),
            .lcout(\nx.n2490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1678_3_lut_LC_10_21_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1678_3_lut_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1678_3_lut_LC_10_21_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1678_3_lut_LC_10_21_5  (
            .in0(N__41723),
            .in1(_gnd_net_),
            .in2(N__41703),
            .in3(N__41636),
            .lcout(\nx.n2491 ),
            .ltout(\nx.n2491_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_56_LC_10_21_6 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_56_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_56_LC_10_21_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_56_LC_10_21_6  (
            .in0(N__38248),
            .in1(N__38315),
            .in2(N__33924),
            .in3(N__38284),
            .lcout(\nx.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1679_3_lut_LC_10_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1679_3_lut_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1679_3_lut_LC_10_21_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1679_3_lut_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__41765),
            .in2(N__41748),
            .in3(N__41635),
            .lcout(\nx.n2492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1611_3_lut_LC_10_22_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1611_3_lut_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1611_3_lut_LC_10_22_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1611_3_lut_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__45828),
            .in2(N__45848),
            .in3(N__44122),
            .lcout(\nx.n2392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1612_3_lut_LC_10_22_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1612_3_lut_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1612_3_lut_LC_10_22_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1612_3_lut_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__45890),
            .in2(N__44129),
            .in3(N__45870),
            .lcout(\nx.n2393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1613_3_lut_LC_10_22_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1613_3_lut_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1613_3_lut_LC_10_22_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1613_3_lut_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__45938),
            .in2(N__45918),
            .in3(N__44118),
            .lcout(\nx.n2394 ),
            .ltout(\nx.n2394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1680_3_lut_LC_10_22_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1680_3_lut_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1680_3_lut_LC_10_22_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1680_3_lut_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__41611),
            .in2(N__34113),
            .in3(N__41790),
            .lcout(\nx.n2493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1424_3_lut_LC_10_22_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1424_3_lut_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1424_3_lut_LC_10_22_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1424_3_lut_LC_10_22_7  (
            .in0(N__34110),
            .in1(N__34083),
            .in2(_gnd_net_),
            .in3(N__34189),
            .lcout(\nx.n2109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1417_3_lut_LC_10_23_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1417_3_lut_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1417_3_lut_LC_10_23_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1417_3_lut_LC_10_23_0  (
            .in0(N__34040),
            .in1(_gnd_net_),
            .in2(N__34197),
            .in3(N__34104),
            .lcout(\nx.n2102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1416_3_lut_LC_10_23_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1416_3_lut_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1416_3_lut_LC_10_23_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1416_3_lut_LC_10_23_1  (
            .in0(N__34659),
            .in1(_gnd_net_),
            .in2(N__34098),
            .in3(N__34183),
            .lcout(\nx.n2101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1423_3_lut_LC_10_23_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1423_3_lut_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1423_3_lut_LC_10_23_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1423_3_lut_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__34089),
            .in2(N__34195),
            .in3(N__34015),
            .lcout(\nx.n2108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_69_LC_10_23_3 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_69_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_69_LC_10_23_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \nx.i11_4_lut_adj_69_LC_10_23_3  (
            .in0(N__34076),
            .in1(N__34039),
            .in2(N__34017),
            .in3(N__34626),
            .lcout(\nx.n27_adj_665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1421_3_lut_LC_10_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1421_3_lut_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1421_3_lut_LC_10_23_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1421_3_lut_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__34404),
            .in2(N__34196),
            .in3(N__34687),
            .lcout(\nx.n2106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1411_3_lut_LC_10_23_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1411_3_lut_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1411_3_lut_LC_10_23_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1411_3_lut_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(N__34398),
            .in2(N__34392),
            .in3(N__34184),
            .lcout(\nx.n2096 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1409_3_lut_LC_10_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1409_3_lut_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1409_3_lut_LC_10_23_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1409_3_lut_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(N__34356),
            .in2(N__34350),
            .in3(N__34185),
            .lcout(\nx.n2094 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_72_LC_10_24_0 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_72_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_72_LC_10_24_0 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \nx.i13_4_lut_adj_72_LC_10_24_0  (
            .in0(N__37081),
            .in1(N__36910),
            .in2(N__36873),
            .in3(N__34311),
            .lcout(),
            .ltout(\nx.n30_adj_668_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_76_LC_10_24_1 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_76_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_76_LC_10_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_76_LC_10_24_1  (
            .in0(N__34245),
            .in1(N__34698),
            .in2(N__34302),
            .in3(N__34299),
            .lcout(\nx.n2126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1422_3_lut_LC_10_24_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1422_3_lut_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1422_3_lut_LC_10_24_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1422_3_lut_LC_10_24_2  (
            .in0(_gnd_net_),
            .in1(N__34289),
            .in2(N__34257),
            .in3(N__34193),
            .lcout(\nx.n2107 ),
            .ltout(\nx.n2107_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_74_LC_10_24_3 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_74_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_74_LC_10_24_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_74_LC_10_24_3  (
            .in0(N__36826),
            .in1(N__36790),
            .in2(N__34248),
            .in3(N__37294),
            .lcout(\nx.n29_adj_670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1412_3_lut_LC_10_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1412_3_lut_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1412_3_lut_LC_10_24_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1412_3_lut_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(N__34239),
            .in2(N__34232),
            .in3(N__34194),
            .lcout(\nx.n2097 ),
            .ltout(\nx.n2097_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_75_LC_10_24_5 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_75_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_75_LC_10_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_75_LC_10_24_5  (
            .in0(N__37060),
            .in1(N__36940),
            .in2(N__34701),
            .in3(N__37270),
            .lcout(\nx.n27_adj_671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9587_1_lut_LC_10_24_6 .C_ON=1'b0;
    defparam \nx.i9587_1_lut_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9587_1_lut_LC_10_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.i9587_1_lut_LC_10_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37193),
            .lcout(\nx.n13436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_2_lut_adj_66_LC_10_25_2 .C_ON=1'b0;
    defparam \nx.i6_2_lut_adj_66_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.i6_2_lut_adj_66_LC_10_25_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i6_2_lut_adj_66_LC_10_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34692),
            .in3(N__34645),
            .lcout(\nx.n22_adj_662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1214_3_lut_LC_10_27_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1214_3_lut_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1214_3_lut_LC_10_27_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1214_3_lut_LC_10_27_0  (
            .in0(_gnd_net_),
            .in1(N__35439),
            .in2(N__35128),
            .in3(N__35403),
            .lcout(\nx.n1803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_83_LC_10_27_1 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_83_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_83_LC_10_27_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_adj_83_LC_10_27_1  (
            .in0(N__34787),
            .in1(N__34741),
            .in2(N__34818),
            .in3(N__35318),
            .lcout(),
            .ltout(\nx.n22_adj_673_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_99_LC_10_27_2 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_99_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_99_LC_10_27_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_99_LC_10_27_2  (
            .in0(N__35278),
            .in1(N__35242),
            .in2(N__34593),
            .in3(N__34590),
            .lcout(\nx.n24_adj_685 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1209_3_lut_LC_10_27_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1209_3_lut_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1209_3_lut_LC_10_27_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1209_3_lut_LC_10_27_3  (
            .in0(_gnd_net_),
            .in1(N__35217),
            .in2(N__35249),
            .in3(N__35108),
            .lcout(\nx.n1798 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1150_rep_76_3_lut_LC_10_27_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1150_rep_76_3_lut_LC_10_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1150_rep_76_3_lut_LC_10_27_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1150_rep_76_3_lut_LC_10_27_4  (
            .in0(_gnd_net_),
            .in1(N__34550),
            .in2(N__34533),
            .in3(N__34516),
            .lcout(\nx.n1707 ),
            .ltout(\nx.n1707_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9517_3_lut_LC_10_27_5 .C_ON=1'b0;
    defparam \nx.i9517_3_lut_LC_10_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9517_3_lut_LC_10_27_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.i9517_3_lut_LC_10_27_5  (
            .in0(_gnd_net_),
            .in1(N__34803),
            .in2(N__34437),
            .in3(N__35107),
            .lcout(\nx.n1806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_110_LC_10_27_6 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_110_LC_10_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_110_LC_10_27_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_110_LC_10_27_6  (
            .in0(N__35393),
            .in1(N__34868),
            .in2(N__35031),
            .in3(N__35016),
            .lcout(\nx.n1730 ),
            .ltout(\nx.n1730_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1213_3_lut_LC_10_27_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1213_3_lut_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1213_3_lut_LC_10_27_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1213_3_lut_LC_10_27_7  (
            .in0(N__35373),
            .in1(_gnd_net_),
            .in2(N__35010),
            .in3(N__35394),
            .lcout(\nx.n1802 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_2_lut_LC_10_28_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_2_lut_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_2_lut_LC_10_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_2_lut_LC_10_28_0  (
            .in0(_gnd_net_),
            .in1(N__34975),
            .in2(_gnd_net_),
            .in3(N__34920),
            .lcout(\nx.n1777 ),
            .ltout(),
            .carryin(bfn_10_28_0_),
            .carryout(\nx.n10615 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_3_lut_LC_10_28_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_3_lut_LC_10_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_3_lut_LC_10_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_3_lut_LC_10_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34917),
            .in3(N__34872),
            .lcout(\nx.n1776 ),
            .ltout(),
            .carryin(\nx.n10615 ),
            .carryout(\nx.n10616 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_4_lut_LC_10_28_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_4_lut_LC_10_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_4_lut_LC_10_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_4_lut_LC_10_28_2  (
            .in0(_gnd_net_),
            .in1(N__44596),
            .in2(N__34867),
            .in3(N__34821),
            .lcout(\nx.n1775 ),
            .ltout(),
            .carryin(\nx.n10616 ),
            .carryout(\nx.n10617 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_5_lut_LC_10_28_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_5_lut_LC_10_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_5_lut_LC_10_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_5_lut_LC_10_28_3  (
            .in0(_gnd_net_),
            .in1(N__34814),
            .in2(N__44955),
            .in3(N__34797),
            .lcout(\nx.n1774 ),
            .ltout(),
            .carryin(\nx.n10617 ),
            .carryout(\nx.n10618 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_6_lut_LC_10_28_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_6_lut_LC_10_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_6_lut_LC_10_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_6_lut_LC_10_28_4  (
            .in0(_gnd_net_),
            .in1(N__44600),
            .in2(N__34794),
            .in3(N__34752),
            .lcout(\nx.n1773 ),
            .ltout(),
            .carryin(\nx.n10618 ),
            .carryout(\nx.n10619 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_7_lut_LC_10_28_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_7_lut_LC_10_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_7_lut_LC_10_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_7_lut_LC_10_28_5  (
            .in0(_gnd_net_),
            .in1(N__44862),
            .in2(N__34742),
            .in3(N__34704),
            .lcout(\nx.n1772 ),
            .ltout(),
            .carryin(\nx.n10619 ),
            .carryout(\nx.n10620 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_8_lut_LC_10_28_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_8_lut_LC_10_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_8_lut_LC_10_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_8_lut_LC_10_28_6  (
            .in0(_gnd_net_),
            .in1(N__44601),
            .in2(N__35438),
            .in3(N__35397),
            .lcout(\nx.n1771 ),
            .ltout(),
            .carryin(\nx.n10620 ),
            .carryout(\nx.n10621 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_9_lut_LC_10_28_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_9_lut_LC_10_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_9_lut_LC_10_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_9_lut_LC_10_28_7  (
            .in0(_gnd_net_),
            .in1(N__44863),
            .in2(N__35392),
            .in3(N__35367),
            .lcout(\nx.n1770 ),
            .ltout(),
            .carryin(\nx.n10621 ),
            .carryout(\nx.n10622 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_10_lut_LC_10_29_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_10_lut_LC_10_29_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_10_lut_LC_10_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_10_lut_LC_10_29_0  (
            .in0(_gnd_net_),
            .in1(N__44433),
            .in2(N__35364),
            .in3(N__35325),
            .lcout(\nx.n1769 ),
            .ltout(),
            .carryin(bfn_10_29_0_),
            .carryout(\nx.n10623 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_11_lut_LC_10_29_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_11_lut_LC_10_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_11_lut_LC_10_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_11_lut_LC_10_29_1  (
            .in0(_gnd_net_),
            .in1(N__44436),
            .in2(N__35322),
            .in3(N__35286),
            .lcout(\nx.n1768 ),
            .ltout(),
            .carryin(\nx.n10623 ),
            .carryout(\nx.n10624 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_12_lut_LC_10_29_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_12_lut_LC_10_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_12_lut_LC_10_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_12_lut_LC_10_29_2  (
            .in0(_gnd_net_),
            .in1(N__35279),
            .in2(N__44716),
            .in3(N__35253),
            .lcout(\nx.n1767 ),
            .ltout(),
            .carryin(\nx.n10624 ),
            .carryout(\nx.n10625 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_13_lut_LC_10_29_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_13_lut_LC_10_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_13_lut_LC_10_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_13_lut_LC_10_29_3  (
            .in0(_gnd_net_),
            .in1(N__44440),
            .in2(N__35250),
            .in3(N__35208),
            .lcout(\nx.n1766 ),
            .ltout(),
            .carryin(\nx.n10625 ),
            .carryout(\nx.n10626 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_14_lut_LC_10_29_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_14_lut_LC_10_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_14_lut_LC_10_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1205_14_lut_LC_10_29_4  (
            .in0(_gnd_net_),
            .in1(N__44434),
            .in2(N__35204),
            .in3(N__35154),
            .lcout(\nx.n1765 ),
            .ltout(),
            .carryin(\nx.n10626 ),
            .carryout(\nx.n10627 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_15_lut_LC_10_29_5 .C_ON=1'b0;
    defparam \nx.mod_5_add_1205_15_lut_LC_10_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_15_lut_LC_10_29_5 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_1205_15_lut_LC_10_29_5  (
            .in0(N__44435),
            .in1(N__35145),
            .in2(N__35073),
            .in3(N__35052),
            .lcout(\nx.n1796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i1_LC_11_14_4.C_ON=1'b0;
    defparam pin_output_enable__i1_LC_11_14_4.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i1_LC_11_14_4.LUT_INIT=16'b0000000000100010;
    LogicCell40 pin_output_enable__i1_LC_11_14_4 (
            .in0(N__50067),
            .in1(N__49838),
            .in2(_gnd_net_),
            .in3(N__49570),
            .lcout(pin_oe_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48421),
            .ce(N__37338),
            .sr(_gnd_net_));
    defparam i2938_3_lut_4_lut_LC_11_15_0.C_ON=1'b0;
    defparam i2938_3_lut_4_lut_LC_11_15_0.SEQ_MODE=4'b0000;
    defparam i2938_3_lut_4_lut_LC_11_15_0.LUT_INIT=16'b1110111100000000;
    LogicCell40 i2938_3_lut_4_lut_LC_11_15_0 (
            .in0(N__38906),
            .in1(N__40401),
            .in2(N__49048),
            .in3(N__46964),
            .lcout(n6158),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_290_i8_2_lut_3_lut_LC_11_15_2.C_ON=1'b0;
    defparam equal_290_i8_2_lut_3_lut_LC_11_15_2.SEQ_MODE=4'b0000;
    defparam equal_290_i8_2_lut_3_lut_LC_11_15_2.LUT_INIT=16'b1111111111111010;
    LogicCell40 equal_290_i8_2_lut_3_lut_LC_11_15_2 (
            .in0(N__48701),
            .in1(_gnd_net_),
            .in2(N__50778),
            .in3(N__50555),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_1101_i22_2_lut_LC_11_15_5.C_ON=1'b0;
    defparam equal_1101_i22_2_lut_LC_11_15_5.SEQ_MODE=4'b0000;
    defparam equal_1101_i22_2_lut_LC_11_15_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 equal_1101_i22_2_lut_LC_11_15_5 (
            .in0(_gnd_net_),
            .in1(N__48700),
            .in2(_gnd_net_),
            .in3(N__50773),
            .lcout(n22_adj_740),
            .ltout(n22_adj_740_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2691_3_lut_4_lut_LC_11_15_6.C_ON=1'b0;
    defparam i2691_3_lut_4_lut_LC_11_15_6.SEQ_MODE=4'b0000;
    defparam i2691_3_lut_4_lut_LC_11_15_6.LUT_INIT=16'b1100110011001000;
    LogicCell40 i2691_3_lut_4_lut_LC_11_15_6 (
            .in0(N__46722),
            .in1(N__46963),
            .in2(N__35475),
            .in3(N__46642),
            .lcout(n5907),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2936_3_lut_4_lut_LC_11_16_0.C_ON=1'b0;
    defparam i2936_3_lut_4_lut_LC_11_16_0.SEQ_MODE=4'b0000;
    defparam i2936_3_lut_4_lut_LC_11_16_0.LUT_INIT=16'b1010101010101000;
    LogicCell40 i2936_3_lut_4_lut_LC_11_16_0 (
            .in0(N__46923),
            .in1(N__40397),
            .in2(N__49049),
            .in3(N__38910),
            .lcout(n6156),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i21_LC_11_16_2.C_ON=1'b0;
    defparam pin_output_i0_i21_LC_11_16_2.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i21_LC_11_16_2.LUT_INIT=16'b0101000011011000;
    LogicCell40 pin_output_i0_i21_LC_11_16_2 (
            .in0(N__39072),
            .in1(N__39084),
            .in2(N__42899),
            .in3(N__46529),
            .lcout(pin_out_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48418),
            .ce(),
            .sr(_gnd_net_));
    defparam i2942_3_lut_4_lut_LC_11_16_5.C_ON=1'b0;
    defparam i2942_3_lut_4_lut_LC_11_16_5.SEQ_MODE=4'b0000;
    defparam i2942_3_lut_4_lut_LC_11_16_5.LUT_INIT=16'b1111000010110000;
    LogicCell40 i2942_3_lut_4_lut_LC_11_16_5 (
            .in0(N__40443),
            .in1(N__50127),
            .in2(N__46958),
            .in3(N__40361),
            .lcout(n6162),
            .ltout(n6162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_163_LC_11_16_6.C_ON=1'b0;
    defparam i1_4_lut_adj_163_LC_11_16_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_163_LC_11_16_6.LUT_INIT=16'b0010111100000000;
    LogicCell40 i1_4_lut_adj_163_LC_11_16_6 (
            .in0(N__43294),
            .in1(N__37480),
            .in2(N__35448),
            .in3(N__47497),
            .lcout(n7278),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_11_17_0.C_ON=1'b0;
    defparam i1_4_lut_LC_11_17_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_11_17_0.LUT_INIT=16'b0000101000101010;
    LogicCell40 i1_4_lut_LC_11_17_0 (
            .in0(N__47422),
            .in1(N__42640),
            .in2(N__35982),
            .in3(N__37481),
            .lcout(),
            .ltout(n7266_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i4_LC_11_17_1.C_ON=1'b0;
    defparam pin_output_i0_i4_LC_11_17_1.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i4_LC_11_17_1.LUT_INIT=16'b0000110010101100;
    LogicCell40 pin_output_i0_i4_LC_11_17_1 (
            .in0(N__35981),
            .in1(N__35947),
            .in2(N__35967),
            .in3(N__46528),
            .lcout(pin_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48414),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_751_i10_2_lut_LC_11_17_5.C_ON=1'b0;
    defparam equal_751_i10_2_lut_LC_11_17_5.SEQ_MODE=4'b0000;
    defparam equal_751_i10_2_lut_LC_11_17_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 equal_751_i10_2_lut_LC_11_17_5 (
            .in0(_gnd_net_),
            .in1(N__50730),
            .in2(_gnd_net_),
            .in3(N__50564),
            .lcout(n10_adj_736),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1764_3_lut_LC_11_18_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1764_3_lut_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1764_3_lut_LC_11_18_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1764_3_lut_LC_11_18_0  (
            .in0(N__37833),
            .in1(N__37892),
            .in2(_gnd_net_),
            .in3(N__39509),
            .lcout(\nx.n2609 ),
            .ltout(\nx.n2609_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_3_lut_LC_11_18_1 .C_ON=1'b0;
    defparam \nx.i6_3_lut_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.i6_3_lut_LC_11_18_1 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \nx.i6_3_lut_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__35899),
            .in2(N__35853),
            .in3(N__37681),
            .lcout(),
            .ltout(\nx.n28_adj_599_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_LC_11_18_2 .C_ON=1'b0;
    defparam \nx.i18_4_lut_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_LC_11_18_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_LC_11_18_2  (
            .in0(N__35821),
            .in1(N__37660),
            .in2(N__35850),
            .in3(N__35847),
            .lcout(\nx.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1753_3_lut_LC_11_18_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1753_3_lut_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1753_3_lut_LC_11_18_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1753_3_lut_LC_11_18_4  (
            .in0(N__38034),
            .in1(_gnd_net_),
            .in2(N__38070),
            .in3(N__39517),
            .lcout(\nx.n2598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1763_3_lut_LC_11_18_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1763_3_lut_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1763_3_lut_LC_11_18_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1763_3_lut_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__37788),
            .in2(N__39538),
            .in3(N__37821),
            .lcout(\nx.n2608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9530_3_lut_LC_11_18_6 .C_ON=1'b0;
    defparam \nx.i9530_3_lut_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9530_3_lut_LC_11_18_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.i9530_3_lut_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__37754),
            .in2(N__37725),
            .in3(N__39513),
            .lcout(\nx.n2604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9520_3_lut_LC_11_18_7 .C_ON=1'b0;
    defparam \nx.i9520_3_lut_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.i9520_3_lut_LC_11_18_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.i9520_3_lut_LC_11_18_7  (
            .in0(N__39597),
            .in1(_gnd_net_),
            .in2(N__39539),
            .in3(N__38085),
            .lcout(\nx.n2599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1751_3_lut_LC_11_19_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1751_3_lut_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1751_3_lut_LC_11_19_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1751_3_lut_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__37989),
            .in2(N__39537),
            .in3(N__38003),
            .lcout(\nx.n2596 ),
            .ltout(\nx.n2596_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_LC_11_19_1 .C_ON=1'b0;
    defparam \nx.i15_4_lut_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_LC_11_19_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_LC_11_19_1  (
            .in0(N__37921),
            .in1(N__36361),
            .in2(N__36342),
            .in3(N__36331),
            .lcout(\nx.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_18_LC_11_19_2 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_18_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_18_LC_11_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_18_LC_11_19_2  (
            .in0(N__36259),
            .in1(N__39412),
            .in2(N__36302),
            .in3(N__36236),
            .lcout(\nx.n38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9526_3_lut_LC_11_19_3 .C_ON=1'b0;
    defparam \nx.i9526_3_lut_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9526_3_lut_LC_11_19_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.i9526_3_lut_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__38142),
            .in2(N__39357),
            .in3(N__39503),
            .lcout(\nx.n2602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1761_3_lut_LC_11_19_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1761_3_lut_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1761_3_lut_LC_11_19_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1761_3_lut_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__37773),
            .in2(N__39536),
            .in3(N__39637),
            .lcout(\nx.n2606 ),
            .ltout(\nx.n2606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1828_3_lut_LC_11_19_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1828_3_lut_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1828_3_lut_LC_11_19_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1828_3_lut_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__36222),
            .in2(N__36213),
            .in3(N__36172),
            .lcout(\nx.n2705 ),
            .ltout(\nx.n2705_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1895_3_lut_LC_11_19_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1895_3_lut_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1895_3_lut_LC_11_19_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1895_3_lut_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__36060),
            .in2(N__36051),
            .in3(N__36586),
            .lcout(\nx.n2804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1749_3_lut_LC_11_19_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1749_3_lut_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1749_3_lut_LC_11_19_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1749_3_lut_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__38328),
            .in2(N__39387),
            .in3(N__39499),
            .lcout(\nx.n2594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9536_3_lut_LC_11_20_0 .C_ON=1'b0;
    defparam \nx.i9536_3_lut_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.i9536_3_lut_LC_11_20_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.i9536_3_lut_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__41061),
            .in2(N__41031),
            .in3(N__41600),
            .lcout(\nx.n2504 ),
            .ltout(\nx.n2504_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9528_3_lut_LC_11_20_1 .C_ON=1'b0;
    defparam \nx.i9528_3_lut_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9528_3_lut_LC_11_20_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.i9528_3_lut_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__37710),
            .in2(N__36690),
            .in3(N__39518),
            .lcout(\nx.n2603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i6_LC_11_20_2.C_ON=1'b0;
    defparam neopxl_color_i6_LC_11_20_2.SEQ_MODE=4'b1001;
    defparam neopxl_color_i6_LC_11_20_2.LUT_INIT=16'b0101010101000000;
    LogicCell40 neopxl_color_i6_LC_11_20_2 (
            .in0(N__49581),
            .in1(N__50034),
            .in2(N__49828),
            .in3(N__40746),
            .lcout(neopxl_color_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48422),
            .ce(),
            .sr(N__40719));
    defparam \nx.mod_5_i1744_3_lut_LC_11_20_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1744_3_lut_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1744_3_lut_LC_11_20_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1744_3_lut_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__39685),
            .in2(N__38187),
            .in3(N__39523),
            .lcout(\nx.n2589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1878_3_lut_LC_11_20_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1878_3_lut_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1878_3_lut_LC_11_20_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1878_3_lut_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(N__36629),
            .in2(N__36609),
            .in3(N__36477),
            .lcout(\nx.n2787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1745_3_lut_LC_11_20_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1745_3_lut_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1745_3_lut_LC_11_20_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1745_3_lut_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__38213),
            .in2(N__39540),
            .in3(N__38199),
            .lcout(\nx.n2590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1746_3_lut_LC_11_20_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1746_3_lut_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1746_3_lut_LC_11_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1746_3_lut_LC_11_20_7  (
            .in0(N__38232),
            .in1(N__38252),
            .in2(_gnd_net_),
            .in3(N__39519),
            .lcout(\nx.n2591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i5_LC_11_21_0.C_ON=1'b0;
    defparam neopxl_color_i5_LC_11_21_0.SEQ_MODE=4'b1001;
    defparam neopxl_color_i5_LC_11_21_0.LUT_INIT=16'b0011001000100010;
    LogicCell40 neopxl_color_i5_LC_11_21_0 (
            .in0(N__39777),
            .in1(N__49580),
            .in2(N__50066),
            .in3(N__49818),
            .lcout(neopxl_color_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48425),
            .ce(),
            .sr(N__39744));
    defparam \nx.mod_5_i1547_3_lut_LC_11_21_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1547_3_lut_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1547_3_lut_LC_11_21_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1547_3_lut_LC_11_21_1  (
            .in0(N__40228),
            .in1(_gnd_net_),
            .in2(N__41988),
            .in3(N__40206),
            .lcout(\nx.n2296 ),
            .ltout(\nx.n2296_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1614_3_lut_LC_11_21_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1614_3_lut_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1614_3_lut_LC_11_21_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1614_3_lut_LC_11_21_2  (
            .in0(N__45960),
            .in1(_gnd_net_),
            .in2(N__36723),
            .in3(N__44127),
            .lcout(\nx.n2395 ),
            .ltout(\nx.n2395_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1681_3_lut_LC_11_21_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1681_3_lut_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1681_3_lut_LC_11_21_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1681_3_lut_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__41826),
            .in2(N__36720),
            .in3(N__41598),
            .lcout(\nx.n2494 ),
            .ltout(\nx.n2494_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1748_3_lut_LC_11_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1748_3_lut_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1748_3_lut_LC_11_21_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1748_3_lut_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__38304),
            .in2(N__36717),
            .in3(N__39526),
            .lcout(\nx.n2593 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9542_3_lut_LC_11_21_5 .C_ON=1'b0;
    defparam \nx.i9542_3_lut_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9542_3_lut_LC_11_21_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.i9542_3_lut_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(N__41442),
            .in2(N__43626),
            .in3(N__41599),
            .lcout(\nx.n2501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9529_3_lut_LC_11_21_6 .C_ON=1'b0;
    defparam \nx.i9529_3_lut_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9529_3_lut_LC_11_21_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.i9529_3_lut_LC_11_21_6  (
            .in0(N__41076),
            .in1(_gnd_net_),
            .in2(N__41631),
            .in3(N__43599),
            .lcout(\nx.n2505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_2_lut_LC_11_21_7 .C_ON=1'b0;
    defparam \nx.i3_2_lut_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.i3_2_lut_LC_11_21_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i3_2_lut_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40230),
            .in3(N__40189),
            .lcout(\nx.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1694_3_lut_LC_11_22_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1694_3_lut_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1694_3_lut_LC_11_22_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1694_3_lut_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__41124),
            .in2(N__41154),
            .in3(N__41594),
            .lcout(\nx.n2507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1545_3_lut_LC_11_22_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1545_3_lut_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1545_3_lut_LC_11_22_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1545_3_lut_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__40151),
            .in2(N__40125),
            .in3(N__41948),
            .lcout(\nx.n2294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1544_3_lut_LC_11_22_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1544_3_lut_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1544_3_lut_LC_11_22_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1544_3_lut_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__40077),
            .in2(N__40106),
            .in3(N__41949),
            .lcout(\nx.n2293 ),
            .ltout(\nx.n2293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_LC_11_22_5 .C_ON=1'b0;
    defparam \nx.i11_4_lut_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_LC_11_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_LC_11_22_5  (
            .in0(N__45934),
            .in1(N__45886),
            .in2(N__36921),
            .in3(N__45971),
            .lcout(\nx.n30_adj_640 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1546_3_lut_LC_11_22_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1546_3_lut_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1546_3_lut_LC_11_22_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1546_3_lut_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__40190),
            .in2(N__41974),
            .in3(N__40167),
            .lcout(\nx.n2295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_2_lut_LC_11_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_2_lut_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_2_lut_LC_11_23_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1473_2_lut_LC_11_23_0  (
            .in0(N__36918),
            .in1(N__36917),
            .in2(N__36848),
            .in3(N__36876),
            .lcout(\nx.n2209 ),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\nx.n10673 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_3_lut_LC_11_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_3_lut_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_3_lut_LC_11_23_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1473_3_lut_LC_11_23_1  (
            .in0(N__36869),
            .in1(N__36868),
            .in2(N__36849),
            .in3(N__36831),
            .lcout(\nx.n2208 ),
            .ltout(),
            .carryin(\nx.n10673 ),
            .carryout(\nx.n10674 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_4_lut_LC_11_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_4_lut_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_4_lut_LC_11_23_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_4_lut_LC_11_23_2  (
            .in0(N__36828),
            .in1(N__36827),
            .in2(N__37242),
            .in3(N__36810),
            .lcout(\nx.n2207 ),
            .ltout(),
            .carryin(\nx.n10674 ),
            .carryout(\nx.n10675 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_5_lut_LC_11_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_5_lut_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_5_lut_LC_11_23_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_5_lut_LC_11_23_3  (
            .in0(N__36807),
            .in1(N__36806),
            .in2(N__37245),
            .in3(N__36795),
            .lcout(\nx.n2206 ),
            .ltout(),
            .carryin(\nx.n10675 ),
            .carryout(\nx.n10676 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_6_lut_LC_11_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_6_lut_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_6_lut_LC_11_23_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_6_lut_LC_11_23_4  (
            .in0(N__36792),
            .in1(N__36791),
            .in2(N__37243),
            .in3(N__36774),
            .lcout(\nx.n2205 ),
            .ltout(),
            .carryin(\nx.n10676 ),
            .carryout(\nx.n10677 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_7_lut_LC_11_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_7_lut_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_7_lut_LC_11_23_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_7_lut_LC_11_23_5  (
            .in0(N__36771),
            .in1(N__36770),
            .in2(N__37246),
            .in3(N__36753),
            .lcout(\nx.n2204 ),
            .ltout(),
            .carryin(\nx.n10677 ),
            .carryout(\nx.n10678 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_8_lut_LC_11_23_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_8_lut_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_8_lut_LC_11_23_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_8_lut_LC_11_23_6  (
            .in0(N__36750),
            .in1(N__36749),
            .in2(N__37244),
            .in3(N__36726),
            .lcout(\nx.n2203 ),
            .ltout(),
            .carryin(\nx.n10678 ),
            .carryout(\nx.n10679 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_9_lut_LC_11_23_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_9_lut_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_9_lut_LC_11_23_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_9_lut_LC_11_23_7  (
            .in0(N__37110),
            .in1(N__37109),
            .in2(N__37247),
            .in3(N__37086),
            .lcout(\nx.n2202 ),
            .ltout(),
            .carryin(\nx.n10679 ),
            .carryout(\nx.n10680 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_10_lut_LC_11_24_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_10_lut_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_10_lut_LC_11_24_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_10_lut_LC_11_24_0  (
            .in0(N__37083),
            .in1(N__37082),
            .in2(N__37248),
            .in3(N__37065),
            .lcout(\nx.n2201 ),
            .ltout(),
            .carryin(bfn_11_24_0_),
            .carryout(\nx.n10681 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_11_lut_LC_11_24_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_11_lut_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_11_lut_LC_11_24_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_11_lut_LC_11_24_1  (
            .in0(N__37062),
            .in1(N__37061),
            .in2(N__37252),
            .in3(N__37044),
            .lcout(\nx.n2200 ),
            .ltout(),
            .carryin(\nx.n10681 ),
            .carryout(\nx.n10682 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_12_lut_LC_11_24_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_12_lut_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_12_lut_LC_11_24_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_12_lut_LC_11_24_2  (
            .in0(N__37041),
            .in1(N__37040),
            .in2(N__37249),
            .in3(N__37014),
            .lcout(\nx.n2199 ),
            .ltout(),
            .carryin(\nx.n10682 ),
            .carryout(\nx.n10683 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_13_lut_LC_11_24_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_13_lut_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_13_lut_LC_11_24_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_13_lut_LC_11_24_3  (
            .in0(N__37011),
            .in1(N__37010),
            .in2(N__37253),
            .in3(N__36993),
            .lcout(\nx.n2198 ),
            .ltout(),
            .carryin(\nx.n10683 ),
            .carryout(\nx.n10684 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_14_lut_LC_11_24_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_14_lut_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_14_lut_LC_11_24_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_14_lut_LC_11_24_4  (
            .in0(N__36990),
            .in1(N__36989),
            .in2(N__37250),
            .in3(N__36963),
            .lcout(\nx.n2197 ),
            .ltout(),
            .carryin(\nx.n10684 ),
            .carryout(\nx.n10685 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_15_lut_LC_11_24_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_15_lut_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_15_lut_LC_11_24_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_15_lut_LC_11_24_5  (
            .in0(N__36960),
            .in1(N__36956),
            .in2(N__37254),
            .in3(N__36945),
            .lcout(\nx.n2196 ),
            .ltout(),
            .carryin(\nx.n10685 ),
            .carryout(\nx.n10686 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_16_lut_LC_11_24_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_16_lut_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_16_lut_LC_11_24_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_16_lut_LC_11_24_6  (
            .in0(N__36942),
            .in1(N__36941),
            .in2(N__37251),
            .in3(N__36924),
            .lcout(\nx.n2195 ),
            .ltout(),
            .carryin(\nx.n10686 ),
            .carryout(\nx.n10687 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_17_lut_LC_11_24_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_17_lut_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_17_lut_LC_11_24_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_17_lut_LC_11_24_7  (
            .in0(N__37329),
            .in1(N__37328),
            .in2(N__37255),
            .in3(N__37305),
            .lcout(\nx.n2194 ),
            .ltout(),
            .carryin(\nx.n10687 ),
            .carryout(\nx.n10688 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_18_lut_LC_11_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_18_lut_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_18_lut_LC_11_25_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_18_lut_LC_11_25_0  (
            .in0(N__37302),
            .in1(N__37301),
            .in2(N__37256),
            .in3(N__37281),
            .lcout(\nx.n2193 ),
            .ltout(),
            .carryin(bfn_11_25_0_),
            .carryout(\nx.n10689 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_19_lut_LC_11_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_add_1473_19_lut_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_19_lut_LC_11_25_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1473_19_lut_LC_11_25_1  (
            .in0(N__37277),
            .in1(N__37278),
            .in2(N__37257),
            .in3(N__37137),
            .lcout(\nx.n2192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7849_4_lut_LC_11_25_3.C_ON=1'b0;
    defparam i7849_4_lut_LC_11_25_3.SEQ_MODE=4'b0000;
    defparam i7849_4_lut_LC_11_25_3.LUT_INIT=16'b1110101010101010;
    LogicCell40 i7849_4_lut_LC_11_25_3 (
            .in0(N__37347),
            .in1(N__38631),
            .in2(N__37134),
            .in3(N__38889),
            .lcout(n11612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_229_LC_11_25_6.C_ON=1'b0;
    defparam i4_4_lut_adj_229_LC_11_25_6.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_229_LC_11_25_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i4_4_lut_adj_229_LC_11_25_6 (
            .in0(N__38673),
            .in1(N__37125),
            .in2(N__38715),
            .in3(N__37443),
            .lcout(n12171),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_11_25_7.C_ON=1'b0;
    defparam i1_2_lut_LC_11_25_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_11_25_7.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_LC_11_25_7 (
            .in0(N__38691),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38652),
            .lcout(n6_adj_761),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_11_26_0.C_ON=1'b0;
    defparam i6_4_lut_LC_11_26_0.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_11_26_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_LC_11_26_0 (
            .in0(N__38378),
            .in1(N__38552),
            .in2(N__38397),
            .in3(N__38537),
            .lcout(),
            .ltout(n15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_LC_11_26_1.C_ON=1'b0;
    defparam i8_4_lut_LC_11_26_1.SEQ_MODE=4'b0000;
    defparam i8_4_lut_LC_11_26_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i8_4_lut_LC_11_26_1 (
            .in0(N__38567),
            .in1(N__38363),
            .in2(N__37119),
            .in3(N__37116),
            .lcout(n12091),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_3_lut_LC_11_26_4.C_ON=1'b0;
    defparam i5_3_lut_LC_11_26_4.SEQ_MODE=4'b0000;
    defparam i5_3_lut_LC_11_26_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 i5_3_lut_LC_11_26_4 (
            .in0(N__38597),
            .in1(N__38582),
            .in2(_gnd_net_),
            .in3(N__38612),
            .lcout(n14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1390_4_lut_LC_11_27_0.C_ON=1'b0;
    defparam i1390_4_lut_LC_11_27_0.SEQ_MODE=4'b0000;
    defparam i1390_4_lut_LC_11_27_0.LUT_INIT=16'b1110101000000000;
    LogicCell40 i1390_4_lut_LC_11_27_0 (
            .in0(N__38504),
            .in1(N__37452),
            .in2(N__38523),
            .in3(N__38489),
            .lcout(),
            .ltout(n24_adj_720_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_226_LC_11_27_1.C_ON=1'b0;
    defparam i2_4_lut_adj_226_LC_11_27_1.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_226_LC_11_27_1.LUT_INIT=16'b1010100000000000;
    LogicCell40 i2_4_lut_adj_226_LC_11_27_1 (
            .in0(N__38744),
            .in1(N__38759),
            .in2(N__37446),
            .in3(N__38729),
            .lcout(n11898),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_228_LC_11_28_0.C_ON=1'b0;
    defparam i7_4_lut_adj_228_LC_11_28_0.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_228_LC_11_28_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i7_4_lut_adj_228_LC_11_28_0 (
            .in0(N__38792),
            .in1(N__39041),
            .in2(N__38856),
            .in3(N__38837),
            .lcout(n17_adj_765),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_195_LC_11_28_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_195_LC_11_28_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_195_LC_11_28_4.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_2_lut_3_lut_adj_195_LC_11_28_4 (
            .in0(N__37416),
            .in1(N__50068),
            .in2(_gnd_net_),
            .in3(N__49834),
            .lcout(n22_adj_724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_227_LC_11_29_6.C_ON=1'b0;
    defparam i6_4_lut_adj_227_LC_11_29_6.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_227_LC_11_29_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_227_LC_11_29_6 (
            .in0(N__39011),
            .in1(N__38807),
            .in2(N__38778),
            .in3(N__39026),
            .lcout(),
            .ltout(n16_adj_764_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_11_29_7.C_ON=1'b0;
    defparam i9_4_lut_LC_11_29_7.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_11_29_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_LC_11_29_7 (
            .in0(N__38870),
            .in1(N__37356),
            .in2(N__37350),
            .in3(N__38822),
            .lcout(n10978),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_32_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_32_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_32_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_32_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_224_LC_12_14_1.C_ON=1'b0;
    defparam i1_4_lut_adj_224_LC_12_14_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_224_LC_12_14_1.LUT_INIT=16'b0000011100000010;
    LogicCell40 i1_4_lut_adj_224_LC_12_14_1 (
            .in0(N__50044),
            .in1(N__49830),
            .in2(N__49588),
            .in3(N__37461),
            .lcout(n36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9315_3_lut_LC_12_14_3.C_ON=1'b0;
    defparam i9315_3_lut_LC_12_14_3.SEQ_MODE=4'b0000;
    defparam i9315_3_lut_LC_12_14_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i9315_3_lut_LC_12_14_3 (
            .in0(N__37544),
            .in1(N__38926),
            .in2(_gnd_net_),
            .in3(N__49033),
            .lcout(n13162),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9564_2_lut_3_lut_LC_12_15_2.C_ON=1'b0;
    defparam i9564_2_lut_3_lut_LC_12_15_2.SEQ_MODE=4'b0000;
    defparam i9564_2_lut_3_lut_LC_12_15_2.LUT_INIT=16'b0000000000010001;
    LogicCell40 i9564_2_lut_3_lut_LC_12_15_2 (
            .in0(N__47163),
            .in1(N__48133),
            .in2(_gnd_net_),
            .in3(N__47230),
            .lcout(state_7_N_167_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_188_LC_12_15_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_188_LC_12_15_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_188_LC_12_15_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_188_LC_12_15_3 (
            .in0(N__47231),
            .in1(N__47164),
            .in2(N__48147),
            .in3(N__49032),
            .lcout(n7166),
            .ltout(n7166_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2932_3_lut_4_lut_LC_12_15_4.C_ON=1'b0;
    defparam i2932_3_lut_4_lut_LC_12_15_4.SEQ_MODE=4'b0000;
    defparam i2932_3_lut_4_lut_LC_12_15_4.LUT_INIT=16'b1111111000000000;
    LogicCell40 i2932_3_lut_4_lut_LC_12_15_4 (
            .in0(N__40664),
            .in1(N__40442),
            .in2(N__37587),
            .in3(N__46944),
            .lcout(n6152),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_282_i8_2_lut_3_lut_LC_12_16_2.C_ON=1'b0;
    defparam equal_282_i8_2_lut_3_lut_LC_12_16_2.SEQ_MODE=4'b0000;
    defparam equal_282_i8_2_lut_3_lut_LC_12_16_2.LUT_INIT=16'b1111111110111011;
    LogicCell40 equal_282_i8_2_lut_3_lut_LC_12_16_2 (
            .in0(N__48699),
            .in1(N__50777),
            .in2(_gnd_net_),
            .in3(N__50573),
            .lcout(n8_adj_751),
            .ltout(n8_adj_751_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_171_LC_12_16_3.C_ON=1'b0;
    defparam i1_4_lut_adj_171_LC_12_16_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_171_LC_12_16_3.LUT_INIT=16'b0000100010101010;
    LogicCell40 i1_4_lut_adj_171_LC_12_16_3 (
            .in0(N__47476),
            .in1(N__43295),
            .in2(N__37566),
            .in3(N__39062),
            .lcout(),
            .ltout(n7294_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i11_LC_12_16_4.C_ON=1'b0;
    defparam pin_output_i0_i11_LC_12_16_4.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i11_LC_12_16_4.LUT_INIT=16'b0000110010101100;
    LogicCell40 pin_output_i0_i11_LC_12_16_4 (
            .in0(N__39063),
            .in1(N__37540),
            .in2(N__37563),
            .in3(N__46518),
            .lcout(pin_out_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48420),
            .ce(),
            .sr(_gnd_net_));
    defparam i2934_3_lut_4_lut_LC_12_16_6.C_ON=1'b0;
    defparam i2934_3_lut_4_lut_LC_12_16_6.SEQ_MODE=4'b0000;
    defparam i2934_3_lut_4_lut_LC_12_16_6.LUT_INIT=16'b1111111000000000;
    LogicCell40 i2934_3_lut_4_lut_LC_12_16_6 (
            .in0(N__40334),
            .in1(N__40657),
            .in2(N__40448),
            .in3(N__46915),
            .lcout(n6154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_284_i8_2_lut_3_lut_LC_12_17_0.C_ON=1'b0;
    defparam equal_284_i8_2_lut_3_lut_LC_12_17_0.SEQ_MODE=4'b0000;
    defparam equal_284_i8_2_lut_3_lut_LC_12_17_0.LUT_INIT=16'b1110111011111111;
    LogicCell40 equal_284_i8_2_lut_3_lut_LC_12_17_0 (
            .in0(N__48698),
            .in1(N__50772),
            .in2(_gnd_net_),
            .in3(N__50534),
            .lcout(n8_adj_744),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9272_2_lut_LC_12_17_4.C_ON=1'b0;
    defparam i9272_2_lut_LC_12_17_4.SEQ_MODE=4'b0000;
    defparam i9272_2_lut_LC_12_17_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i9272_2_lut_LC_12_17_4 (
            .in0(_gnd_net_),
            .in1(N__48482),
            .in2(_gnd_net_),
            .in3(N__48527),
            .lcout(),
            .ltout(n13048_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9443_4_lut_LC_12_17_5.C_ON=1'b0;
    defparam i9443_4_lut_LC_12_17_5.SEQ_MODE=4'b0000;
    defparam i9443_4_lut_LC_12_17_5.LUT_INIT=16'b0000000000000100;
    LogicCell40 i9443_4_lut_LC_12_17_5 (
            .in0(N__39053),
            .in1(N__47654),
            .in2(N__37464),
            .in3(N__48572),
            .lcout(n13264),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9434_3_lut_4_lut_LC_12_18_1.C_ON=1'b0;
    defparam i9434_3_lut_4_lut_LC_12_18_1.SEQ_MODE=4'b0000;
    defparam i9434_3_lut_4_lut_LC_12_18_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9434_3_lut_4_lut_LC_12_18_1 (
            .in0(N__48573),
            .in1(N__39054),
            .in2(N__48492),
            .in3(N__48534),
            .lcout(n13273),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_12_18_2.C_ON=1'b0;
    defparam i1_3_lut_LC_12_18_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_12_18_2.LUT_INIT=16'b0000000001100110;
    LogicCell40 i1_3_lut_LC_12_18_2 (
            .in0(N__50007),
            .in1(N__49771),
            .in2(_gnd_net_),
            .in3(N__49510),
            .lcout(n7231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1752_3_lut_LC_12_18_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1752_3_lut_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1752_3_lut_LC_12_18_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1752_3_lut_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__39729),
            .in2(N__38022),
            .in3(N__39525),
            .lcout(\nx.n2597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9524_3_lut_LC_12_18_7 .C_ON=1'b0;
    defparam \nx.i9524_3_lut_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.i9524_3_lut_LC_12_18_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.i9524_3_lut_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__38133),
            .in2(N__39324),
            .in3(N__39524),
            .lcout(\nx.n2601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1684_3_lut_LC_12_19_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1684_3_lut_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1684_3_lut_LC_12_19_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1684_3_lut_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__43233),
            .in2(N__41334),
            .in3(N__41660),
            .lcout(\nx.n2497 ),
            .ltout(\nx.n2497_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_3_lut_LC_12_19_2 .C_ON=1'b0;
    defparam \nx.i5_3_lut_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.i5_3_lut_LC_12_19_2 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i5_3_lut_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__37896),
            .in2(N__37641),
            .in3(N__37820),
            .lcout(),
            .ltout(\nx.n26_adj_611_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_24_LC_12_19_3 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_24_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_24_LC_12_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_24_LC_12_19_3  (
            .in0(N__37974),
            .in1(N__39376),
            .in2(N__37638),
            .in3(N__37635),
            .lcout(),
            .ltout(\nx.n38_adj_612_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_adj_48_LC_12_19_4 .C_ON=1'b0;
    defparam \nx.i20_4_lut_adj_48_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_adj_48_LC_12_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i20_4_lut_adj_48_LC_12_19_4  (
            .in0(N__37902),
            .in1(N__39606),
            .in2(N__37623),
            .in3(N__39330),
            .lcout(\nx.n2522 ),
            .ltout(\nx.n2522_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9522_3_lut_LC_12_19_5 .C_ON=1'b0;
    defparam \nx.i9522_3_lut_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9522_3_lut_LC_12_19_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \nx.i9522_3_lut_LC_12_19_5  (
            .in0(N__38121),
            .in1(N__38097),
            .in2(N__37620),
            .in3(_gnd_net_),
            .lcout(\nx.n2600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9532_3_lut_LC_12_19_6 .C_ON=1'b0;
    defparam \nx.i9532_3_lut_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9532_3_lut_LC_12_19_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.i9532_3_lut_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__37764),
            .in2(N__39273),
            .in3(N__39508),
            .lcout(\nx.n2605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_46_LC_12_19_7 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_46_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_46_LC_12_19_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_46_LC_12_19_7  (
            .in0(N__38120),
            .in1(N__38065),
            .in2(N__37755),
            .in3(N__39724),
            .lcout(\nx.n35_adj_639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_2_lut_LC_12_20_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_2_lut_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_2_lut_LC_12_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_2_lut_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__37891),
            .in2(_gnd_net_),
            .in3(N__37824),
            .lcout(\nx.n2577 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\nx.n10747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_3_lut_LC_12_20_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_3_lut_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_3_lut_LC_12_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_3_lut_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37819),
            .in3(N__37779),
            .lcout(\nx.n2576 ),
            .ltout(),
            .carryin(\nx.n10747 ),
            .carryout(\nx.n10748 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_4_lut_LC_12_20_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_4_lut_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_4_lut_LC_12_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_4_lut_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__45450),
            .in2(N__39296),
            .in3(N__37776),
            .lcout(\nx.n2575 ),
            .ltout(),
            .carryin(\nx.n10748 ),
            .carryout(\nx.n10749 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_5_lut_LC_12_20_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_5_lut_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_5_lut_LC_12_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_5_lut_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__45453),
            .in2(N__39638),
            .in3(N__37767),
            .lcout(\nx.n2574 ),
            .ltout(),
            .carryin(\nx.n10749 ),
            .carryout(\nx.n10750 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_6_lut_LC_12_20_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_6_lut_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_6_lut_LC_12_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_6_lut_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__45451),
            .in2(N__39272),
            .in3(N__37758),
            .lcout(\nx.n2573 ),
            .ltout(),
            .carryin(\nx.n10750 ),
            .carryout(\nx.n10751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_7_lut_LC_12_20_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_7_lut_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_7_lut_LC_12_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_7_lut_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__45454),
            .in2(N__37744),
            .in3(N__37713),
            .lcout(\nx.n2572 ),
            .ltout(),
            .carryin(\nx.n10751 ),
            .carryout(\nx.n10752 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_8_lut_LC_12_20_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_8_lut_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_8_lut_LC_12_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_8_lut_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__45452),
            .in2(N__39659),
            .in3(N__38145),
            .lcout(\nx.n2571 ),
            .ltout(),
            .carryin(\nx.n10752 ),
            .carryout(\nx.n10753 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_9_lut_LC_12_20_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_9_lut_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_9_lut_LC_12_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_9_lut_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(N__45455),
            .in2(N__39350),
            .in3(N__38136),
            .lcout(\nx.n2570 ),
            .ltout(),
            .carryin(\nx.n10753 ),
            .carryout(\nx.n10754 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_10_lut_LC_12_21_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_10_lut_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_10_lut_LC_12_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_10_lut_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__45440),
            .in2(N__39320),
            .in3(N__38124),
            .lcout(\nx.n2569 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\nx.n10755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_11_lut_LC_12_21_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_11_lut_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_11_lut_LC_12_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_11_lut_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(N__45025),
            .in2(N__38114),
            .in3(N__38088),
            .lcout(\nx.n2568 ),
            .ltout(),
            .carryin(\nx.n10755 ),
            .carryout(\nx.n10756 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_12_lut_LC_12_21_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_12_lut_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_12_lut_LC_12_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_12_lut_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(N__45441),
            .in2(N__39593),
            .in3(N__38073),
            .lcout(\nx.n2567 ),
            .ltout(),
            .carryin(\nx.n10756 ),
            .carryout(\nx.n10757 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_13_lut_LC_12_21_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_13_lut_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_13_lut_LC_12_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_13_lut_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(N__45026),
            .in2(N__38066),
            .in3(N__38025),
            .lcout(\nx.n2566 ),
            .ltout(),
            .carryin(\nx.n10757 ),
            .carryout(\nx.n10758 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_14_lut_LC_12_21_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_14_lut_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_14_lut_LC_12_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_14_lut_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(N__45442),
            .in2(N__39728),
            .in3(N__38010),
            .lcout(\nx.n2565 ),
            .ltout(),
            .carryin(\nx.n10758 ),
            .carryout(\nx.n10759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_15_lut_LC_12_21_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_15_lut_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_15_lut_LC_12_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_15_lut_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__45027),
            .in2(N__38007),
            .in3(N__37977),
            .lcout(\nx.n2564 ),
            .ltout(),
            .carryin(\nx.n10759 ),
            .carryout(\nx.n10760 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_16_lut_LC_12_21_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_16_lut_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_16_lut_LC_12_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_16_lut_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__45443),
            .in2(N__37973),
            .in3(N__37935),
            .lcout(\nx.n2563 ),
            .ltout(),
            .carryin(\nx.n10760 ),
            .carryout(\nx.n10761 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_17_lut_LC_12_21_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_17_lut_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_17_lut_LC_12_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_17_lut_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(N__45028),
            .in2(N__39380),
            .in3(N__38319),
            .lcout(\nx.n2562 ),
            .ltout(),
            .carryin(\nx.n10761 ),
            .carryout(\nx.n10762 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_18_lut_LC_12_22_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_18_lut_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_18_lut_LC_12_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_18_lut_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__38316),
            .in2(N__45438),
            .in3(N__38298),
            .lcout(\nx.n2561 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\nx.n10763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_19_lut_LC_12_22_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_19_lut_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_19_lut_LC_12_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_19_lut_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(N__38291),
            .in2(N__45437),
            .in3(N__38259),
            .lcout(\nx.n2560 ),
            .ltout(),
            .carryin(\nx.n10763 ),
            .carryout(\nx.n10764 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_20_lut_LC_12_22_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_20_lut_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_20_lut_LC_12_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_20_lut_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__38256),
            .in2(N__45439),
            .in3(N__38223),
            .lcout(\nx.n2559 ),
            .ltout(),
            .carryin(\nx.n10764 ),
            .carryout(\nx.n10765 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_21_lut_LC_12_22_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_21_lut_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_21_lut_LC_12_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_21_lut_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(N__45036),
            .in2(N__38220),
            .in3(N__38190),
            .lcout(\nx.n2558 ),
            .ltout(),
            .carryin(\nx.n10765 ),
            .carryout(\nx.n10766 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_22_lut_LC_12_22_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_22_lut_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_22_lut_LC_12_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_22_lut_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(N__45023),
            .in2(N__39693),
            .in3(N__38175),
            .lcout(\nx.n2557 ),
            .ltout(),
            .carryin(\nx.n10766 ),
            .carryout(\nx.n10767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_23_lut_LC_12_22_5 .C_ON=1'b0;
    defparam \nx.mod_5_add_1741_23_lut_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_23_lut_LC_12_22_5 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1741_23_lut_LC_12_22_5  (
            .in0(N__45024),
            .in1(N__41538),
            .in2(N__39549),
            .in3(N__38172),
            .lcout(\nx.n2588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_51_LC_12_22_6 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_51_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_51_LC_12_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_51_LC_12_22_6  (
            .in0(N__43852),
            .in1(N__43936),
            .in2(N__43451),
            .in3(N__43399),
            .lcout(\nx.n33_adj_644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_47_LC_12_22_7 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_47_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_47_LC_12_22_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_47_LC_12_22_7  (
            .in0(N__43899),
            .in1(N__44147),
            .in2(N__45810),
            .in3(N__38349),
            .lcout(\nx.n34_adj_641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1559_3_lut_LC_12_23_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1559_3_lut_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1559_3_lut_LC_12_23_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1559_3_lut_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(N__40057),
            .in2(N__40035),
            .in3(N__41932),
            .lcout(\nx.n2308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_LC_12_23_2 .C_ON=1'b0;
    defparam \nx.i16_4_lut_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_LC_12_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_LC_12_23_2  (
            .in0(N__39949),
            .in1(N__42208),
            .in2(N__38475),
            .in3(N__38466),
            .lcout(),
            .ltout(\nx.n34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_LC_12_23_3 .C_ON=1'b0;
    defparam \nx.i17_4_lut_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_LC_12_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_LC_12_23_3  (
            .in0(N__38403),
            .in1(N__38409),
            .in2(N__38343),
            .in3(N__38340),
            .lcout(\nx.n2225 ),
            .ltout(\nx.n2225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1556_3_lut_LC_12_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1556_3_lut_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1556_3_lut_LC_12_23_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1556_3_lut_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__39963),
            .in2(N__38331),
            .in3(N__39983),
            .lcout(\nx.n2305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1560_3_lut_LC_12_23_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1560_3_lut_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1560_3_lut_LC_12_23_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1560_3_lut_LC_12_23_5  (
            .in0(N__39804),
            .in1(N__39858),
            .in2(_gnd_net_),
            .in3(N__41928),
            .lcout(\nx.n2309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1558_3_lut_LC_12_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1558_3_lut_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1558_3_lut_LC_12_23_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1558_3_lut_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(N__39999),
            .in2(N__41957),
            .in3(N__40022),
            .lcout(\nx.n2307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1555_3_lut_LC_12_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1555_3_lut_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1555_3_lut_LC_12_23_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1555_3_lut_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(N__39950),
            .in2(N__39933),
            .in3(N__41933),
            .lcout(\nx.n2304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6426_2_lut_LC_12_24_0 .C_ON=1'b0;
    defparam \nx.i6426_2_lut_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.i6426_2_lut_LC_12_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \nx.i6426_2_lut_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__43567),
            .in2(_gnd_net_),
            .in3(N__43486),
            .lcout(\nx.n9650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_78_LC_12_24_1 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_78_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_78_LC_12_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_78_LC_12_24_1  (
            .in0(N__41506),
            .in1(N__40018),
            .in2(N__42124),
            .in3(N__42076),
            .lcout(\nx.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_77_LC_12_24_2 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_77_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_77_LC_12_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_77_LC_12_24_2  (
            .in0(N__40141),
            .in1(N__40090),
            .in2(N__42013),
            .in3(N__40376),
            .lcout(\nx.n28_adj_601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i12_LC_12_24_4.C_ON=1'b0;
    defparam neopxl_color_prev_i12_LC_12_24_4.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i12_LC_12_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 neopxl_color_prev_i12_LC_12_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38460),
            .lcout(neopxl_color_prev_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48439),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_LC_12_24_5 .C_ON=1'b0;
    defparam \nx.i12_4_lut_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_LC_12_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_LC_12_24_5  (
            .in0(N__40273),
            .in1(N__39910),
            .in2(N__42056),
            .in3(N__39982),
            .lcout(\nx.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_3_lut_adj_79_LC_12_24_7 .C_ON=1'b0;
    defparam \nx.i4_3_lut_adj_79_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.i4_3_lut_adj_79_LC_12_24_7 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \nx.i4_3_lut_adj_79_LC_12_24_7  (
            .in0(N__39857),
            .in1(_gnd_net_),
            .in2(N__40059),
            .in3(N__42169),
            .lcout(\nx.n22_adj_604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_223_LC_12_25_5.C_ON=1'b0;
    defparam i2_3_lut_adj_223_LC_12_25_5.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_223_LC_12_25_5.LUT_INIT=16'b0010001000000000;
    LogicCell40 i2_3_lut_adj_223_LC_12_25_5 (
            .in0(N__40806),
            .in1(N__47711),
            .in2(_gnd_net_),
            .in3(N__47678),
            .lcout(n7442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_counter_1104__i0_LC_12_26_0.C_ON=1'b1;
    defparam delay_counter_1104__i0_LC_12_26_0.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i0_LC_12_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i0_LC_12_26_0 (
            .in0(_gnd_net_),
            .in1(N__38396),
            .in2(_gnd_net_),
            .in3(N__38382),
            .lcout(delay_counter_0),
            .ltout(),
            .carryin(bfn_12_26_0_),
            .carryout(n10517),
            .clk(N__48445),
            .ce(N__40812),
            .sr(N__38976));
    defparam delay_counter_1104__i1_LC_12_26_1.C_ON=1'b1;
    defparam delay_counter_1104__i1_LC_12_26_1.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i1_LC_12_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i1_LC_12_26_1 (
            .in0(_gnd_net_),
            .in1(N__38379),
            .in2(_gnd_net_),
            .in3(N__38367),
            .lcout(delay_counter_1),
            .ltout(),
            .carryin(n10517),
            .carryout(n10518),
            .clk(N__48445),
            .ce(N__40812),
            .sr(N__38976));
    defparam delay_counter_1104__i2_LC_12_26_2.C_ON=1'b1;
    defparam delay_counter_1104__i2_LC_12_26_2.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i2_LC_12_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i2_LC_12_26_2 (
            .in0(_gnd_net_),
            .in1(N__38364),
            .in2(_gnd_net_),
            .in3(N__38352),
            .lcout(delay_counter_2),
            .ltout(),
            .carryin(n10518),
            .carryout(n10519),
            .clk(N__48445),
            .ce(N__40812),
            .sr(N__38976));
    defparam delay_counter_1104__i3_LC_12_26_3.C_ON=1'b1;
    defparam delay_counter_1104__i3_LC_12_26_3.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i3_LC_12_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i3_LC_12_26_3 (
            .in0(_gnd_net_),
            .in1(N__38613),
            .in2(_gnd_net_),
            .in3(N__38601),
            .lcout(delay_counter_3),
            .ltout(),
            .carryin(n10519),
            .carryout(n10520),
            .clk(N__48445),
            .ce(N__40812),
            .sr(N__38976));
    defparam delay_counter_1104__i4_LC_12_26_4.C_ON=1'b1;
    defparam delay_counter_1104__i4_LC_12_26_4.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i4_LC_12_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i4_LC_12_26_4 (
            .in0(_gnd_net_),
            .in1(N__38598),
            .in2(_gnd_net_),
            .in3(N__38586),
            .lcout(delay_counter_4),
            .ltout(),
            .carryin(n10520),
            .carryout(n10521),
            .clk(N__48445),
            .ce(N__40812),
            .sr(N__38976));
    defparam delay_counter_1104__i5_LC_12_26_5.C_ON=1'b1;
    defparam delay_counter_1104__i5_LC_12_26_5.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i5_LC_12_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i5_LC_12_26_5 (
            .in0(_gnd_net_),
            .in1(N__38583),
            .in2(_gnd_net_),
            .in3(N__38571),
            .lcout(delay_counter_5),
            .ltout(),
            .carryin(n10521),
            .carryout(n10522),
            .clk(N__48445),
            .ce(N__40812),
            .sr(N__38976));
    defparam delay_counter_1104__i6_LC_12_26_6.C_ON=1'b1;
    defparam delay_counter_1104__i6_LC_12_26_6.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i6_LC_12_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i6_LC_12_26_6 (
            .in0(_gnd_net_),
            .in1(N__38568),
            .in2(_gnd_net_),
            .in3(N__38556),
            .lcout(delay_counter_6),
            .ltout(),
            .carryin(n10522),
            .carryout(n10523),
            .clk(N__48445),
            .ce(N__40812),
            .sr(N__38976));
    defparam delay_counter_1104__i7_LC_12_26_7.C_ON=1'b1;
    defparam delay_counter_1104__i7_LC_12_26_7.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i7_LC_12_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i7_LC_12_26_7 (
            .in0(_gnd_net_),
            .in1(N__38553),
            .in2(_gnd_net_),
            .in3(N__38541),
            .lcout(delay_counter_7),
            .ltout(),
            .carryin(n10523),
            .carryout(n10524),
            .clk(N__48445),
            .ce(N__40812),
            .sr(N__38976));
    defparam delay_counter_1104__i8_LC_12_27_0.C_ON=1'b1;
    defparam delay_counter_1104__i8_LC_12_27_0.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i8_LC_12_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i8_LC_12_27_0 (
            .in0(_gnd_net_),
            .in1(N__38538),
            .in2(_gnd_net_),
            .in3(N__38526),
            .lcout(delay_counter_8),
            .ltout(),
            .carryin(bfn_12_27_0_),
            .carryout(n10525),
            .clk(N__48447),
            .ce(N__40820),
            .sr(N__38993));
    defparam delay_counter_1104__i9_LC_12_27_1.C_ON=1'b1;
    defparam delay_counter_1104__i9_LC_12_27_1.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i9_LC_12_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i9_LC_12_27_1 (
            .in0(_gnd_net_),
            .in1(N__38522),
            .in2(_gnd_net_),
            .in3(N__38508),
            .lcout(delay_counter_9),
            .ltout(),
            .carryin(n10525),
            .carryout(n10526),
            .clk(N__48447),
            .ce(N__40820),
            .sr(N__38993));
    defparam delay_counter_1104__i10_LC_12_27_2.C_ON=1'b1;
    defparam delay_counter_1104__i10_LC_12_27_2.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i10_LC_12_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i10_LC_12_27_2 (
            .in0(_gnd_net_),
            .in1(N__38505),
            .in2(_gnd_net_),
            .in3(N__38493),
            .lcout(delay_counter_10),
            .ltout(),
            .carryin(n10526),
            .carryout(n10527),
            .clk(N__48447),
            .ce(N__40820),
            .sr(N__38993));
    defparam delay_counter_1104__i11_LC_12_27_3.C_ON=1'b1;
    defparam delay_counter_1104__i11_LC_12_27_3.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i11_LC_12_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i11_LC_12_27_3 (
            .in0(_gnd_net_),
            .in1(N__38490),
            .in2(_gnd_net_),
            .in3(N__38478),
            .lcout(delay_counter_11),
            .ltout(),
            .carryin(n10527),
            .carryout(n10528),
            .clk(N__48447),
            .ce(N__40820),
            .sr(N__38993));
    defparam delay_counter_1104__i12_LC_12_27_4.C_ON=1'b1;
    defparam delay_counter_1104__i12_LC_12_27_4.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i12_LC_12_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i12_LC_12_27_4 (
            .in0(_gnd_net_),
            .in1(N__38760),
            .in2(_gnd_net_),
            .in3(N__38748),
            .lcout(delay_counter_12),
            .ltout(),
            .carryin(n10528),
            .carryout(n10529),
            .clk(N__48447),
            .ce(N__40820),
            .sr(N__38993));
    defparam delay_counter_1104__i13_LC_12_27_5.C_ON=1'b1;
    defparam delay_counter_1104__i13_LC_12_27_5.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i13_LC_12_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i13_LC_12_27_5 (
            .in0(_gnd_net_),
            .in1(N__38745),
            .in2(_gnd_net_),
            .in3(N__38733),
            .lcout(delay_counter_13),
            .ltout(),
            .carryin(n10529),
            .carryout(n10530),
            .clk(N__48447),
            .ce(N__40820),
            .sr(N__38993));
    defparam delay_counter_1104__i14_LC_12_27_6.C_ON=1'b1;
    defparam delay_counter_1104__i14_LC_12_27_6.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i14_LC_12_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i14_LC_12_27_6 (
            .in0(_gnd_net_),
            .in1(N__38730),
            .in2(_gnd_net_),
            .in3(N__38718),
            .lcout(delay_counter_14),
            .ltout(),
            .carryin(n10530),
            .carryout(n10531),
            .clk(N__48447),
            .ce(N__40820),
            .sr(N__38993));
    defparam delay_counter_1104__i15_LC_12_27_7.C_ON=1'b1;
    defparam delay_counter_1104__i15_LC_12_27_7.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i15_LC_12_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i15_LC_12_27_7 (
            .in0(_gnd_net_),
            .in1(N__38708),
            .in2(_gnd_net_),
            .in3(N__38694),
            .lcout(delay_counter_15),
            .ltout(),
            .carryin(n10531),
            .carryout(n10532),
            .clk(N__48447),
            .ce(N__40820),
            .sr(N__38993));
    defparam delay_counter_1104__i16_LC_12_28_0.C_ON=1'b1;
    defparam delay_counter_1104__i16_LC_12_28_0.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i16_LC_12_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i16_LC_12_28_0 (
            .in0(_gnd_net_),
            .in1(N__38690),
            .in2(_gnd_net_),
            .in3(N__38676),
            .lcout(delay_counter_16),
            .ltout(),
            .carryin(bfn_12_28_0_),
            .carryout(n10533),
            .clk(N__48448),
            .ce(N__40813),
            .sr(N__38989));
    defparam delay_counter_1104__i17_LC_12_28_1.C_ON=1'b1;
    defparam delay_counter_1104__i17_LC_12_28_1.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i17_LC_12_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i17_LC_12_28_1 (
            .in0(_gnd_net_),
            .in1(N__38669),
            .in2(_gnd_net_),
            .in3(N__38655),
            .lcout(delay_counter_17),
            .ltout(),
            .carryin(n10533),
            .carryout(n10534),
            .clk(N__48448),
            .ce(N__40813),
            .sr(N__38989));
    defparam delay_counter_1104__i18_LC_12_28_2.C_ON=1'b1;
    defparam delay_counter_1104__i18_LC_12_28_2.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i18_LC_12_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i18_LC_12_28_2 (
            .in0(_gnd_net_),
            .in1(N__38648),
            .in2(_gnd_net_),
            .in3(N__38634),
            .lcout(delay_counter_18),
            .ltout(),
            .carryin(n10534),
            .carryout(n10535),
            .clk(N__48448),
            .ce(N__40813),
            .sr(N__38989));
    defparam delay_counter_1104__i19_LC_12_28_3.C_ON=1'b1;
    defparam delay_counter_1104__i19_LC_12_28_3.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i19_LC_12_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i19_LC_12_28_3 (
            .in0(_gnd_net_),
            .in1(N__38630),
            .in2(_gnd_net_),
            .in3(N__38616),
            .lcout(delay_counter_19),
            .ltout(),
            .carryin(n10535),
            .carryout(n10536),
            .clk(N__48448),
            .ce(N__40813),
            .sr(N__38989));
    defparam delay_counter_1104__i20_LC_12_28_4.C_ON=1'b1;
    defparam delay_counter_1104__i20_LC_12_28_4.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i20_LC_12_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i20_LC_12_28_4 (
            .in0(_gnd_net_),
            .in1(N__38888),
            .in2(_gnd_net_),
            .in3(N__38874),
            .lcout(delay_counter_20),
            .ltout(),
            .carryin(n10536),
            .carryout(n10537),
            .clk(N__48448),
            .ce(N__40813),
            .sr(N__38989));
    defparam delay_counter_1104__i21_LC_12_28_5.C_ON=1'b1;
    defparam delay_counter_1104__i21_LC_12_28_5.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i21_LC_12_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i21_LC_12_28_5 (
            .in0(_gnd_net_),
            .in1(N__38871),
            .in2(_gnd_net_),
            .in3(N__38859),
            .lcout(delay_counter_21),
            .ltout(),
            .carryin(n10537),
            .carryout(n10538),
            .clk(N__48448),
            .ce(N__40813),
            .sr(N__38989));
    defparam delay_counter_1104__i22_LC_12_28_6.C_ON=1'b1;
    defparam delay_counter_1104__i22_LC_12_28_6.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i22_LC_12_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i22_LC_12_28_6 (
            .in0(_gnd_net_),
            .in1(N__38855),
            .in2(_gnd_net_),
            .in3(N__38841),
            .lcout(delay_counter_22),
            .ltout(),
            .carryin(n10538),
            .carryout(n10539),
            .clk(N__48448),
            .ce(N__40813),
            .sr(N__38989));
    defparam delay_counter_1104__i23_LC_12_28_7.C_ON=1'b1;
    defparam delay_counter_1104__i23_LC_12_28_7.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i23_LC_12_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i23_LC_12_28_7 (
            .in0(_gnd_net_),
            .in1(N__38838),
            .in2(_gnd_net_),
            .in3(N__38826),
            .lcout(delay_counter_23),
            .ltout(),
            .carryin(n10539),
            .carryout(n10540),
            .clk(N__48448),
            .ce(N__40813),
            .sr(N__38989));
    defparam delay_counter_1104__i24_LC_12_29_0.C_ON=1'b1;
    defparam delay_counter_1104__i24_LC_12_29_0.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i24_LC_12_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i24_LC_12_29_0 (
            .in0(_gnd_net_),
            .in1(N__38823),
            .in2(_gnd_net_),
            .in3(N__38811),
            .lcout(delay_counter_24),
            .ltout(),
            .carryin(bfn_12_29_0_),
            .carryout(n10541),
            .clk(N__48449),
            .ce(N__40824),
            .sr(N__38994));
    defparam delay_counter_1104__i25_LC_12_29_1.C_ON=1'b1;
    defparam delay_counter_1104__i25_LC_12_29_1.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i25_LC_12_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i25_LC_12_29_1 (
            .in0(_gnd_net_),
            .in1(N__38808),
            .in2(_gnd_net_),
            .in3(N__38796),
            .lcout(delay_counter_25),
            .ltout(),
            .carryin(n10541),
            .carryout(n10542),
            .clk(N__48449),
            .ce(N__40824),
            .sr(N__38994));
    defparam delay_counter_1104__i26_LC_12_29_2.C_ON=1'b1;
    defparam delay_counter_1104__i26_LC_12_29_2.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i26_LC_12_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i26_LC_12_29_2 (
            .in0(_gnd_net_),
            .in1(N__38793),
            .in2(_gnd_net_),
            .in3(N__38781),
            .lcout(delay_counter_26),
            .ltout(),
            .carryin(n10542),
            .carryout(n10543),
            .clk(N__48449),
            .ce(N__40824),
            .sr(N__38994));
    defparam delay_counter_1104__i27_LC_12_29_3.C_ON=1'b1;
    defparam delay_counter_1104__i27_LC_12_29_3.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i27_LC_12_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i27_LC_12_29_3 (
            .in0(_gnd_net_),
            .in1(N__38777),
            .in2(_gnd_net_),
            .in3(N__38763),
            .lcout(delay_counter_27),
            .ltout(),
            .carryin(n10543),
            .carryout(n10544),
            .clk(N__48449),
            .ce(N__40824),
            .sr(N__38994));
    defparam delay_counter_1104__i28_LC_12_29_4.C_ON=1'b1;
    defparam delay_counter_1104__i28_LC_12_29_4.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i28_LC_12_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i28_LC_12_29_4 (
            .in0(_gnd_net_),
            .in1(N__39042),
            .in2(_gnd_net_),
            .in3(N__39030),
            .lcout(delay_counter_28),
            .ltout(),
            .carryin(n10544),
            .carryout(n10545),
            .clk(N__48449),
            .ce(N__40824),
            .sr(N__38994));
    defparam delay_counter_1104__i29_LC_12_29_5.C_ON=1'b1;
    defparam delay_counter_1104__i29_LC_12_29_5.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i29_LC_12_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i29_LC_12_29_5 (
            .in0(_gnd_net_),
            .in1(N__39027),
            .in2(_gnd_net_),
            .in3(N__39015),
            .lcout(delay_counter_29),
            .ltout(),
            .carryin(n10545),
            .carryout(n10546),
            .clk(N__48449),
            .ce(N__40824),
            .sr(N__38994));
    defparam delay_counter_1104__i30_LC_12_29_6.C_ON=1'b1;
    defparam delay_counter_1104__i30_LC_12_29_6.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i30_LC_12_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i30_LC_12_29_6 (
            .in0(_gnd_net_),
            .in1(N__39012),
            .in2(_gnd_net_),
            .in3(N__39000),
            .lcout(delay_counter_30),
            .ltout(),
            .carryin(n10546),
            .carryout(n10547),
            .clk(N__48449),
            .ce(N__40824),
            .sr(N__38994));
    defparam delay_counter_1104__i31_LC_12_29_7.C_ON=1'b0;
    defparam delay_counter_1104__i31_LC_12_29_7.SEQ_MODE=4'b1000;
    defparam delay_counter_1104__i31_LC_12_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_1104__i31_LC_12_29_7 (
            .in0(_gnd_net_),
            .in1(N__47707),
            .in2(_gnd_net_),
            .in3(N__38997),
            .lcout(delay_counter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(N__40824),
            .sr(N__38994));
    defparam i1_3_lut_4_lut_adj_245_LC_13_14_0.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_245_LC_13_14_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_245_LC_13_14_0.LUT_INIT=16'b1100110011001000;
    LogicCell40 i1_3_lut_4_lut_adj_245_LC_13_14_0 (
            .in0(N__42262),
            .in1(N__46980),
            .in2(N__40665),
            .in3(N__46657),
            .lcout(n10_adj_779),
            .ltout(n10_adj_779_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_169_LC_13_14_1.C_ON=1'b0;
    defparam i1_4_lut_adj_169_LC_13_14_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_169_LC_13_14_1.LUT_INIT=16'b0000110001001100;
    LogicCell40 i1_4_lut_adj_169_LC_13_14_1 (
            .in0(N__42455),
            .in1(N__47505),
            .in2(N__38955),
            .in3(N__47994),
            .lcout(),
            .ltout(n7290_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i10_LC_13_14_2.C_ON=1'b0;
    defparam pin_output_i0_i10_LC_13_14_2.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i10_LC_13_14_2.LUT_INIT=16'b0000110010101100;
    LogicCell40 pin_output_i0_i10_LC_13_14_2 (
            .in0(N__38952),
            .in1(N__38927),
            .in2(N__38946),
            .in3(N__46535),
            .lcout(pin_out_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48428),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_230_LC_13_15_3.C_ON=1'b0;
    defparam i1_2_lut_adj_230_LC_13_15_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_230_LC_13_15_3.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_230_LC_13_15_3 (
            .in0(_gnd_net_),
            .in1(N__47168),
            .in2(_gnd_net_),
            .in3(N__47236),
            .lcout(n7135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_189_LC_13_15_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_189_LC_13_15_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_189_LC_13_15_4.LUT_INIT=16'b1111111011111111;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_189_LC_13_15_4 (
            .in0(N__47235),
            .in1(N__48137),
            .in2(N__47176),
            .in3(N__49017),
            .lcout(n7155),
            .ltout(n7155_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2954_3_lut_4_lut_LC_13_15_5.C_ON=1'b0;
    defparam i2954_3_lut_4_lut_LC_13_15_5.SEQ_MODE=4'b0000;
    defparam i2954_3_lut_4_lut_LC_13_15_5.LUT_INIT=16'b1111111000000000;
    LogicCell40 i2954_3_lut_4_lut_LC_13_15_5 (
            .in0(N__42252),
            .in1(N__42326),
            .in2(N__39087),
            .in3(N__46940),
            .lcout(n6174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2970_3_lut_4_lut_LC_13_16_0.C_ON=1'b0;
    defparam i2970_3_lut_4_lut_LC_13_16_0.SEQ_MODE=4'b0000;
    defparam i2970_3_lut_4_lut_LC_13_16_0.LUT_INIT=16'b1100110011001000;
    LogicCell40 i2970_3_lut_4_lut_LC_13_16_0 (
            .in0(N__42327),
            .in1(N__46970),
            .in2(N__40362),
            .in3(N__46776),
            .lcout(n6190),
            .ltout(n6190_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_197_LC_13_16_1.C_ON=1'b0;
    defparam i1_4_lut_adj_197_LC_13_16_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_197_LC_13_16_1.LUT_INIT=16'b0000101000101010;
    LogicCell40 i1_4_lut_adj_197_LC_13_16_1 (
            .in0(N__47458),
            .in1(N__42715),
            .in2(N__39075),
            .in3(N__47290),
            .lcout(n7334),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2950_3_lut_4_lut_LC_13_16_3.C_ON=1'b0;
    defparam i2950_3_lut_4_lut_LC_13_16_3.SEQ_MODE=4'b0000;
    defparam i2950_3_lut_4_lut_LC_13_16_3.LUT_INIT=16'b1111000011100000;
    LogicCell40 i2950_3_lut_4_lut_LC_13_16_3 (
            .in0(N__40351),
            .in1(N__42261),
            .in2(N__46979),
            .in3(N__40656),
            .lcout(n6170),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_217_LC_13_16_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_217_LC_13_16_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_217_LC_13_16_4.LUT_INIT=16'b0000000000000100;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_217_LC_13_16_4 (
            .in0(N__47238),
            .in1(N__49803),
            .in2(N__47181),
            .in3(N__48149),
            .lcout(n11481),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6193_2_lut_LC_13_17_0.C_ON=1'b0;
    defparam i6193_2_lut_LC_13_17_0.SEQ_MODE=4'b0000;
    defparam i6193_2_lut_LC_13_17_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i6193_2_lut_LC_13_17_0 (
            .in0(N__50771),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48697),
            .lcout(n9415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2966_3_lut_4_lut_LC_13_17_1.C_ON=1'b0;
    defparam i2966_3_lut_4_lut_LC_13_17_1.SEQ_MODE=4'b0000;
    defparam i2966_3_lut_4_lut_LC_13_17_1.LUT_INIT=16'b1111000011100000;
    LogicCell40 i2966_3_lut_4_lut_LC_13_17_1 (
            .in0(N__46774),
            .in1(N__40648),
            .in2(N__46978),
            .in3(N__40354),
            .lcout(n6186),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i404_4_lut_LC_13_17_2.C_ON=1'b0;
    defparam i404_4_lut_LC_13_17_2.SEQ_MODE=4'b0000;
    defparam i404_4_lut_LC_13_17_2.LUT_INIT=16'b1100110011001000;
    LogicCell40 i404_4_lut_LC_13_17_2 (
            .in0(N__40609),
            .in1(N__39248),
            .in2(N__50358),
            .in3(N__48920),
            .lcout(n2337),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2962_3_lut_4_lut_LC_13_17_4.C_ON=1'b0;
    defparam i2962_3_lut_4_lut_LC_13_17_4.SEQ_MODE=4'b0000;
    defparam i2962_3_lut_4_lut_LC_13_17_4.LUT_INIT=16'b1111111000000000;
    LogicCell40 i2962_3_lut_4_lut_LC_13_17_4 (
            .in0(N__40353),
            .in1(N__46775),
            .in2(N__46745),
            .in3(N__46969),
            .lcout(n6182),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_270_i8_2_lut_3_lut_LC_13_17_5.C_ON=1'b0;
    defparam equal_270_i8_2_lut_3_lut_LC_13_17_5.SEQ_MODE=4'b0000;
    defparam equal_270_i8_2_lut_3_lut_LC_13_17_5.LUT_INIT=16'b1101110111111111;
    LogicCell40 equal_270_i8_2_lut_3_lut_LC_13_17_5 (
            .in0(N__48696),
            .in1(N__50770),
            .in2(_gnd_net_),
            .in3(N__50533),
            .lcout(n8_adj_723),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_0__bdd_4_lut_LC_13_17_6.C_ON=1'b0;
    defparam current_pin_0__bdd_4_lut_LC_13_17_6.SEQ_MODE=4'b0000;
    defparam current_pin_0__bdd_4_lut_LC_13_17_6.LUT_INIT=16'b1011101111000000;
    LogicCell40 current_pin_0__bdd_4_lut_LC_13_17_6 (
            .in0(N__40703),
            .in1(N__50262),
            .in2(N__39194),
            .in3(N__48919),
            .lcout(),
            .ltout(n13480_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13480_bdd_4_lut_LC_13_17_7.C_ON=1'b0;
    defparam n13480_bdd_4_lut_LC_13_17_7.SEQ_MODE=4'b0000;
    defparam n13480_bdd_4_lut_LC_13_17_7.LUT_INIT=16'b1111001011000010;
    LogicCell40 n13480_bdd_4_lut_LC_13_17_7 (
            .in0(N__39249),
            .in1(N__50348),
            .in2(N__39231),
            .in3(N__40583),
            .lcout(n13483),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_13_18_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_13_18_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_13_18_1.LUT_INIT=16'b0001000100000000;
    LogicCell40 i1_2_lut_3_lut_LC_13_18_1 (
            .in0(N__50005),
            .in1(N__49758),
            .in2(_gnd_net_),
            .in3(N__49508),
            .lcout(),
            .ltout(current_pin_7__N_157_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16_4_lut_LC_13_18_2.C_ON=1'b0;
    defparam i16_4_lut_LC_13_18_2.SEQ_MODE=4'b0000;
    defparam i16_4_lut_LC_13_18_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i16_4_lut_LC_13_18_2 (
            .in0(N__47617),
            .in1(N__39093),
            .in2(N__39228),
            .in3(N__50006),
            .lcout(n45_adj_772),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i356_3_lut_4_lut_LC_13_18_4.C_ON=1'b0;
    defparam i356_3_lut_4_lut_LC_13_18_4.SEQ_MODE=4'b0000;
    defparam i356_3_lut_4_lut_LC_13_18_4.LUT_INIT=16'b1100110011001000;
    LogicCell40 i356_3_lut_4_lut_LC_13_18_4 (
            .in0(N__47797),
            .in1(N__39225),
            .in2(N__42626),
            .in3(N__42831),
            .lcout(),
            .ltout(n2289_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_13_18_5.C_ON=1'b0;
    defparam i10_4_lut_LC_13_18_5.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_13_18_5.LUT_INIT=16'b1111110011111000;
    LogicCell40 i10_4_lut_LC_13_18_5 (
            .in0(N__47992),
            .in1(N__39195),
            .in2(N__39153),
            .in3(N__40610),
            .lcout(n39),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i392_4_lut_LC_13_18_7.C_ON=1'b0;
    defparam i392_4_lut_LC_13_18_7.SEQ_MODE=4'b0000;
    defparam i392_4_lut_LC_13_18_7.LUT_INIT=16'b1111000011100000;
    LogicCell40 i392_4_lut_LC_13_18_7 (
            .in0(N__47991),
            .in1(N__50616),
            .in2(N__39150),
            .in3(N__47796),
            .lcout(n2325),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9515_3_lut_LC_13_19_0.C_ON=1'b0;
    defparam i9515_3_lut_LC_13_19_0.SEQ_MODE=4'b0000;
    defparam i9515_3_lut_LC_13_19_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 i9515_3_lut_LC_13_19_0 (
            .in0(N__50756),
            .in1(N__39108),
            .in2(_gnd_net_),
            .in3(N__39561),
            .lcout(),
            .ltout(n13364_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i37_4_lut_LC_13_19_1.C_ON=1'b0;
    defparam i37_4_lut_LC_13_19_1.SEQ_MODE=4'b0000;
    defparam i37_4_lut_LC_13_19_1.LUT_INIT=16'b0110011000111100;
    LogicCell40 i37_4_lut_LC_13_19_1 (
            .in0(N__47808),
            .in1(N__46451),
            .in2(N__39096),
            .in3(N__48682),
            .lcout(n150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6204_2_lut_LC_13_19_3.C_ON=1'b0;
    defparam i6204_2_lut_LC_13_19_3.SEQ_MODE=4'b0000;
    defparam i6204_2_lut_LC_13_19_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 i6204_2_lut_LC_13_19_3 (
            .in0(N__50337),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49016),
            .lcout(n9426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9511_3_lut_LC_13_19_4.C_ON=1'b0;
    defparam i9511_3_lut_LC_13_19_4.SEQ_MODE=4'b0000;
    defparam i9511_3_lut_LC_13_19_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 i9511_3_lut_LC_13_19_4 (
            .in0(N__50569),
            .in1(N__40959),
            .in2(_gnd_net_),
            .in3(N__39570),
            .lcout(n13360),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1762_3_lut_LC_13_19_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1762_3_lut_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1762_3_lut_LC_13_19_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1762_3_lut_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__39555),
            .in2(N__39297),
            .in3(N__39507),
            .lcout(\nx.n2607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1682_3_lut_LC_13_20_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1682_3_lut_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1682_3_lut_LC_13_20_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1682_3_lut_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__41881),
            .in2(N__41301),
            .in3(N__41653),
            .lcout(\nx.n2495 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9538_3_lut_LC_13_20_1 .C_ON=1'b0;
    defparam \nx.i9538_3_lut_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9538_3_lut_LC_13_20_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.i9538_3_lut_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__40998),
            .in2(N__41663),
            .in3(N__41012),
            .lcout(\nx.n2503 ),
            .ltout(\nx.n2503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_44_LC_13_20_2 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_44_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_44_LC_13_20_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_44_LC_13_20_2  (
            .in0(N__39268),
            .in1(N__39316),
            .in2(N__39333),
            .in3(N__39292),
            .lcout(\nx.n36_adj_636 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9540_3_lut_LC_13_20_3 .C_ON=1'b0;
    defparam \nx.i9540_3_lut_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9540_3_lut_LC_13_20_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.i9540_3_lut_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__43663),
            .in2(N__41664),
            .in3(N__41451),
            .lcout(\nx.n2502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1695_rep_30_3_lut_LC_13_20_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1695_rep_30_3_lut_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1695_rep_30_3_lut_LC_13_20_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1695_rep_30_3_lut_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__41163),
            .in2(N__41203),
            .in3(N__41640),
            .lcout(\nx.n2508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9534_3_lut_LC_13_20_5 .C_ON=1'b0;
    defparam \nx.i9534_3_lut_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9534_3_lut_LC_13_20_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.i9534_3_lut_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__41085),
            .in2(N__41662),
            .in3(N__41109),
            .lcout(\nx.n2506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_205_LC_13_20_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_205_LC_13_20_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_205_LC_13_20_6.LUT_INIT=16'b1100110010001000;
    LogicCell40 i1_2_lut_3_lut_adj_205_LC_13_20_6 (
            .in0(N__49753),
            .in1(N__39778),
            .in2(_gnd_net_),
            .in3(N__50001),
            .lcout(n22_adj_730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1685_3_lut_LC_13_20_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1685_3_lut_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1685_3_lut_LC_13_20_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1685_3_lut_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__41366),
            .in2(N__41665),
            .in3(N__41346),
            .lcout(\nx.n2498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1622_3_lut_LC_13_21_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1622_3_lut_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1622_3_lut_LC_13_21_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1622_3_lut_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__43941),
            .in2(N__43917),
            .in3(N__44081),
            .lcout(\nx.n2403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1623_3_lut_LC_13_21_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1623_3_lut_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1623_3_lut_LC_13_21_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1623_3_lut_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__43956),
            .in2(N__43986),
            .in3(N__44082),
            .lcout(\nx.n2404 ),
            .ltout(\nx.n2404_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_61_LC_13_21_3 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_61_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_61_LC_13_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_61_LC_13_21_3  (
            .in0(N__43232),
            .in1(N__41104),
            .in2(N__39705),
            .in3(N__41362),
            .lcout(\nx.n34_adj_657 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_57_LC_13_21_4 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_57_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_57_LC_13_21_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i1_2_lut_adj_57_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41537),
            .in3(N__39686),
            .lcout(),
            .ltout(\nx.n22_adj_637_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_45_LC_13_21_5 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_45_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_45_LC_13_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_45_LC_13_21_5  (
            .in0(N__39663),
            .in1(N__39586),
            .in2(N__39642),
            .in3(N__39639),
            .lcout(\nx.n37_adj_638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9544_3_lut_LC_13_21_6 .C_ON=1'b0;
    defparam \nx.i9544_3_lut_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9544_3_lut_LC_13_21_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.i9544_3_lut_LC_13_21_6  (
            .in0(N__41669),
            .in1(N__41394),
            .in2(N__41423),
            .in3(_gnd_net_),
            .lcout(\nx.n2500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1618_3_lut_LC_13_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1618_3_lut_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1618_3_lut_LC_13_21_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1618_3_lut_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__43752),
            .in2(N__44116),
            .in3(N__43766),
            .lcout(\nx.n2399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1626_3_lut_LC_13_22_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1626_3_lut_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1626_3_lut_LC_13_22_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1626_3_lut_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__43425),
            .in2(N__44117),
            .in3(N__43447),
            .lcout(\nx.n2407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1627_3_lut_LC_13_22_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1627_3_lut_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1627_3_lut_LC_13_22_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1627_3_lut_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__43490),
            .in2(N__43470),
            .in3(N__44086),
            .lcout(\nx.n2408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1553_3_lut_LC_13_22_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1553_3_lut_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1553_3_lut_LC_13_22_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1553_3_lut_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__39891),
            .in2(N__39918),
            .in3(N__41953),
            .lcout(\nx.n2302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1551_3_lut_LC_13_22_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1551_3_lut_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1551_3_lut_LC_13_22_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1551_3_lut_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__40278),
            .in2(N__41976),
            .in3(N__40251),
            .lcout(\nx.n2300 ),
            .ltout(\nx.n2300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_50_LC_13_22_4 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_50_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_50_LC_13_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_50_LC_13_22_4  (
            .in0(N__43810),
            .in1(N__43975),
            .in2(N__39879),
            .in3(N__43369),
            .lcout(),
            .ltout(\nx.n32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_53_LC_13_22_5 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_53_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_53_LC_13_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_53_LC_13_22_5  (
            .in0(N__39876),
            .in1(N__39870),
            .in2(N__39864),
            .in3(N__42144),
            .lcout(\nx.n2324 ),
            .ltout(\nx.n2324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9497_3_lut_LC_13_22_6 .C_ON=1'b0;
    defparam \nx.i9497_3_lut_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9497_3_lut_LC_13_22_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.i9497_3_lut_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(N__43353),
            .in2(N__39861),
            .in3(N__43370),
            .lcout(\nx.n2405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9489_3_lut_LC_13_22_7 .C_ON=1'b0;
    defparam \nx.i9489_3_lut_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.i9489_3_lut_LC_13_22_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.i9489_3_lut_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(N__43853),
            .in2(N__43833),
            .in3(N__44090),
            .lcout(\nx.n2401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_2_lut_LC_13_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_2_lut_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_2_lut_LC_13_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_2_lut_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__39856),
            .in2(_gnd_net_),
            .in3(N__39798),
            .lcout(\nx.n2277 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\nx.n10690 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_3_lut_LC_13_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_3_lut_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_3_lut_LC_13_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_3_lut_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__40058),
            .in2(_gnd_net_),
            .in3(N__40026),
            .lcout(\nx.n2276 ),
            .ltout(),
            .carryin(\nx.n10690 ),
            .carryout(\nx.n10691 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_4_lut_LC_13_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_4_lut_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_4_lut_LC_13_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_4_lut_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__45571),
            .in2(N__40023),
            .in3(N__39993),
            .lcout(\nx.n2275 ),
            .ltout(),
            .carryin(\nx.n10691 ),
            .carryout(\nx.n10692 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_5_lut_LC_13_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_5_lut_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_5_lut_LC_13_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_5_lut_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(N__44644),
            .in2(N__41513),
            .in3(N__39990),
            .lcout(\nx.n2274 ),
            .ltout(),
            .carryin(\nx.n10692 ),
            .carryout(\nx.n10693 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_6_lut_LC_13_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_6_lut_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_6_lut_LC_13_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_6_lut_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__45572),
            .in2(N__39987),
            .in3(N__39957),
            .lcout(\nx.n2273 ),
            .ltout(),
            .carryin(\nx.n10693 ),
            .carryout(\nx.n10694 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_7_lut_LC_13_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_7_lut_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_7_lut_LC_13_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_7_lut_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__44645),
            .in2(N__39954),
            .in3(N__39924),
            .lcout(\nx.n2272 ),
            .ltout(),
            .carryin(\nx.n10694 ),
            .carryout(\nx.n10695 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_8_lut_LC_13_23_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_8_lut_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_8_lut_LC_13_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_8_lut_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__42209),
            .in2(N__45019),
            .in3(N__39921),
            .lcout(\nx.n2271 ),
            .ltout(),
            .carryin(\nx.n10695 ),
            .carryout(\nx.n10696 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_9_lut_LC_13_23_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_9_lut_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_9_lut_LC_13_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_9_lut_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__39911),
            .in2(N__45731),
            .in3(N__39885),
            .lcout(\nx.n2270 ),
            .ltout(),
            .carryin(\nx.n10696 ),
            .carryout(\nx.n10697 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_10_lut_LC_13_24_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_10_lut_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_10_lut_LC_13_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_10_lut_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__45218),
            .in2(N__42129),
            .in3(N__39882),
            .lcout(\nx.n2269 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\nx.n10698 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_11_lut_LC_13_24_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_11_lut_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_11_lut_LC_13_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_11_lut_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__45227),
            .in2(N__40277),
            .in3(N__40242),
            .lcout(\nx.n2268 ),
            .ltout(),
            .carryin(\nx.n10698 ),
            .carryout(\nx.n10699 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_12_lut_LC_13_24_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_12_lut_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_12_lut_LC_13_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_12_lut_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__45219),
            .in2(N__42089),
            .in3(N__40239),
            .lcout(\nx.n2267 ),
            .ltout(),
            .carryin(\nx.n10699 ),
            .carryout(\nx.n10700 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_13_lut_LC_13_24_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_13_lut_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_13_lut_LC_13_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_13_lut_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__42052),
            .in2(N__45568),
            .in3(N__40236),
            .lcout(\nx.n2266 ),
            .ltout(),
            .carryin(\nx.n10700 ),
            .carryout(\nx.n10701 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_14_lut_LC_13_24_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_14_lut_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_14_lut_LC_13_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_14_lut_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__45223),
            .in2(N__42182),
            .in3(N__40233),
            .lcout(\nx.n2265 ),
            .ltout(),
            .carryin(\nx.n10701 ),
            .carryout(\nx.n10702 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_15_lut_LC_13_24_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_15_lut_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_15_lut_LC_13_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_15_lut_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__40229),
            .in2(N__45569),
            .in3(N__40194),
            .lcout(\nx.n2264 ),
            .ltout(),
            .carryin(\nx.n10702 ),
            .carryout(\nx.n10703 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_16_lut_LC_13_24_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_16_lut_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_16_lut_LC_13_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_16_lut_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__40191),
            .in2(N__45570),
            .in3(N__40155),
            .lcout(\nx.n2263 ),
            .ltout(),
            .carryin(\nx.n10703 ),
            .carryout(\nx.n10704 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_17_lut_LC_13_24_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_17_lut_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_17_lut_LC_13_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_17_lut_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__45231),
            .in2(N__40152),
            .in3(N__40110),
            .lcout(\nx.n2262 ),
            .ltout(),
            .carryin(\nx.n10704 ),
            .carryout(\nx.n10705 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_18_lut_LC_13_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_18_lut_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_18_lut_LC_13_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_18_lut_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__44859),
            .in2(N__40107),
            .in3(N__40065),
            .lcout(\nx.n2261 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\nx.n10706 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_19_lut_LC_13_25_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_19_lut_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_19_lut_LC_13_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_19_lut_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__44860),
            .in2(N__42020),
            .in3(N__40062),
            .lcout(\nx.n2260 ),
            .ltout(),
            .carryin(\nx.n10706 ),
            .carryout(\nx.n10707 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_20_lut_LC_13_25_2 .C_ON=1'b0;
    defparam \nx.mod_5_add_1540_20_lut_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_20_lut_LC_13_25_2 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_1540_20_lut_LC_13_25_2  (
            .in0(N__44861),
            .in1(N__41975),
            .in2(N__40383),
            .in3(N__40365),
            .lcout(\nx.n2291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1628_3_lut_LC_13_25_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1628_3_lut_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1628_3_lut_LC_13_25_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1628_3_lut_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(N__43509),
            .in2(N__44123),
            .in3(N__43571),
            .lcout(\nx.n2409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2958_3_lut_4_lut_LC_14_15_0.C_ON=1'b0;
    defparam i2958_3_lut_4_lut_LC_14_15_0.SEQ_MODE=4'b0000;
    defparam i2958_3_lut_4_lut_LC_14_15_0.LUT_INIT=16'b1100110011000100;
    LogicCell40 i2958_3_lut_4_lut_LC_14_15_0 (
            .in0(N__50128),
            .in1(N__46941),
            .in2(N__42264),
            .in3(N__40346),
            .lcout(n6178),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i9_LC_14_15_1.C_ON=1'b0;
    defparam pin_output_i0_i9_LC_14_15_1.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i9_LC_14_15_1.LUT_INIT=16'b0101000011011000;
    LogicCell40 pin_output_i0_i9_LC_14_15_1 (
            .in0(N__40287),
            .in1(N__40296),
            .in2(N__42494),
            .in3(N__46517),
            .lcout(pin_out_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48429),
            .ce(),
            .sr(_gnd_net_));
    defparam i2946_3_lut_4_lut_LC_14_15_2.C_ON=1'b0;
    defparam i2946_3_lut_4_lut_LC_14_15_2.SEQ_MODE=4'b0000;
    defparam i2946_3_lut_4_lut_LC_14_15_2.LUT_INIT=16'b1100110011001000;
    LogicCell40 i2946_3_lut_4_lut_LC_14_15_2 (
            .in0(N__42260),
            .in1(N__46942),
            .in2(N__46746),
            .in3(N__40347),
            .lcout(n6166),
            .ltout(n6166_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_167_LC_14_15_3.C_ON=1'b0;
    defparam i1_4_lut_adj_167_LC_14_15_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_167_LC_14_15_3.LUT_INIT=16'b0000110001001100;
    LogicCell40 i1_4_lut_adj_167_LC_14_15_3 (
            .in0(N__42456),
            .in1(N__47526),
            .in2(N__40290),
            .in3(N__42726),
            .lcout(n7286),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_282_i7_2_lut_LC_14_15_4.C_ON=1'b0;
    defparam equal_282_i7_2_lut_LC_14_15_4.SEQ_MODE=4'b0000;
    defparam equal_282_i7_2_lut_LC_14_15_4.LUT_INIT=16'b1100110011111111;
    LogicCell40 equal_282_i7_2_lut_LC_14_15_4 (
            .in0(_gnd_net_),
            .in1(N__48691),
            .in2(_gnd_net_),
            .in3(N__50758),
            .lcout(n7_adj_753),
            .ltout(n7_adj_753_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2944_3_lut_4_lut_LC_14_15_5.C_ON=1'b0;
    defparam i2944_3_lut_4_lut_LC_14_15_5.SEQ_MODE=4'b0000;
    defparam i2944_3_lut_4_lut_LC_14_15_5.LUT_INIT=16'b1010101010101000;
    LogicCell40 i2944_3_lut_4_lut_LC_14_15_5 (
            .in0(N__46943),
            .in1(N__46743),
            .in2(N__40281),
            .in3(N__46677),
            .lcout(n6164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i13_LC_14_15_7.C_ON=1'b0;
    defparam pin_output_i0_i13_LC_14_15_7.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i13_LC_14_15_7.LUT_INIT=16'b0101000011011000;
    LogicCell40 pin_output_i0_i13_LC_14_15_7 (
            .in0(N__42270),
            .in1(N__42284),
            .in2(N__48073),
            .in3(N__46516),
            .lcout(pin_out_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48429),
            .ce(),
            .sr(_gnd_net_));
    defparam i2968_3_lut_4_lut_LC_14_16_0.C_ON=1'b0;
    defparam i2968_3_lut_4_lut_LC_14_16_0.SEQ_MODE=4'b0000;
    defparam i2968_3_lut_4_lut_LC_14_16_0.LUT_INIT=16'b1100110011001000;
    LogicCell40 i2968_3_lut_4_lut_LC_14_16_0 (
            .in0(N__42324),
            .in1(N__46916),
            .in2(N__46688),
            .in3(N__46788),
            .lcout(n6188),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_1098_i21_2_lut_LC_14_16_2.C_ON=1'b0;
    defparam equal_1098_i21_2_lut_LC_14_16_2.SEQ_MODE=4'b0000;
    defparam equal_1098_i21_2_lut_LC_14_16_2.LUT_INIT=16'b1111111101010101;
    LogicCell40 equal_1098_i21_2_lut_LC_14_16_2 (
            .in0(N__50354),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50557),
            .lcout(n21_adj_714),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_238_LC_14_16_3.C_ON=1'b0;
    defparam i12_4_lut_adj_238_LC_14_16_3.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_238_LC_14_16_3.LUT_INIT=16'b1110111011101100;
    LogicCell40 i12_4_lut_adj_238_LC_14_16_3 (
            .in0(N__40479),
            .in1(N__40671),
            .in2(N__49349),
            .in3(N__47795),
            .lcout(n41),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_1100_i21_2_lut_LC_14_16_6.C_ON=1'b0;
    defparam equal_1100_i21_2_lut_LC_14_16_6.SEQ_MODE=4'b0000;
    defparam equal_1100_i21_2_lut_LC_14_16_6.LUT_INIT=16'b1010101011111111;
    LogicCell40 equal_1100_i21_2_lut_LC_14_16_6 (
            .in0(N__50355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50558),
            .lcout(n21_adj_741),
            .ltout(n21_adj_741_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_LC_14_16_7.C_ON=1'b0;
    defparam i2_3_lut_LC_14_16_7.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_14_16_7.LUT_INIT=16'b1111111111111100;
    LogicCell40 i2_3_lut_LC_14_16_7 (
            .in0(_gnd_net_),
            .in1(N__40449),
            .in2(N__40404),
            .in3(N__48148),
            .lcout(n7128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_879_i9_2_lut_LC_14_17_0.C_ON=1'b0;
    defparam equal_879_i9_2_lut_LC_14_17_0.SEQ_MODE=4'b0000;
    defparam equal_879_i9_2_lut_LC_14_17_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 equal_879_i9_2_lut_LC_14_17_0 (
            .in0(_gnd_net_),
            .in1(N__50263),
            .in2(_gnd_net_),
            .in3(N__48921),
            .lcout(n9_adj_733),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_903_i11_2_lut_4_lut_LC_14_17_1.C_ON=1'b0;
    defparam equal_903_i11_2_lut_4_lut_LC_14_17_1.SEQ_MODE=4'b0000;
    defparam equal_903_i11_2_lut_4_lut_LC_14_17_1.LUT_INIT=16'b1111111111011111;
    LogicCell40 equal_903_i11_2_lut_4_lut_LC_14_17_1 (
            .in0(N__50264),
            .in1(N__50722),
            .in2(N__48994),
            .in3(N__50544),
            .lcout(n11_adj_743),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_231_LC_14_17_2.C_ON=1'b0;
    defparam i1_2_lut_adj_231_LC_14_17_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_231_LC_14_17_2.LUT_INIT=16'b1111111101010101;
    LogicCell40 i1_2_lut_adj_231_LC_14_17_2 (
            .in0(N__48666),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47263),
            .lcout(n14_adj_752),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_274_i8_2_lut_3_lut_LC_14_17_3.C_ON=1'b0;
    defparam equal_274_i8_2_lut_3_lut_LC_14_17_3.SEQ_MODE=4'b0000;
    defparam equal_274_i8_2_lut_3_lut_LC_14_17_3.LUT_INIT=16'b1110111011111111;
    LogicCell40 equal_274_i8_2_lut_3_lut_LC_14_17_3 (
            .in0(N__50532),
            .in1(N__50726),
            .in2(_gnd_net_),
            .in3(N__48671),
            .lcout(n8_adj_746),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_215_LC_14_17_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_215_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_215_LC_14_17_4.LUT_INIT=16'b1111111111111101;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_215_LC_14_17_4 (
            .in0(N__50721),
            .in1(N__50531),
            .in2(N__48695),
            .in3(N__47264),
            .lcout(n7150),
            .ltout(n7150_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i422_4_lut_LC_14_17_5.C_ON=1'b0;
    defparam i422_4_lut_LC_14_17_5.SEQ_MODE=4'b0000;
    defparam i422_4_lut_LC_14_17_5.LUT_INIT=16'b1111011100000000;
    LogicCell40 i422_4_lut_LC_14_17_5 (
            .in0(N__50265),
            .in1(N__49004),
            .in2(N__40710),
            .in3(N__40707),
            .lcout(n2355),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_273_i7_2_lut_LC_14_17_6.C_ON=1'b0;
    defparam equal_273_i7_2_lut_LC_14_17_6.SEQ_MODE=4'b0000;
    defparam equal_273_i7_2_lut_LC_14_17_6.LUT_INIT=16'b1111010111110101;
    LogicCell40 equal_273_i7_2_lut_LC_14_17_6 (
            .in0(N__48670),
            .in1(_gnd_net_),
            .in2(N__50757),
            .in3(_gnd_net_),
            .lcout(n7_adj_719),
            .ltout(n7_adj_719_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2964_3_lut_4_lut_LC_14_17_7.C_ON=1'b0;
    defparam i2964_3_lut_4_lut_LC_14_17_7.SEQ_MODE=4'b0000;
    defparam i2964_3_lut_4_lut_LC_14_17_7.LUT_INIT=16'b1100110011001000;
    LogicCell40 i2964_3_lut_4_lut_LC_14_17_7 (
            .in0(N__40655),
            .in1(N__46977),
            .in2(N__40614),
            .in3(N__46687),
            .lcout(n6184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i410_4_lut_LC_14_18_0.C_ON=1'b0;
    defparam i410_4_lut_LC_14_18_0.SEQ_MODE=4'b0000;
    defparam i410_4_lut_LC_14_18_0.LUT_INIT=16'b1110000011110000;
    LogicCell40 i410_4_lut_LC_14_18_0 (
            .in0(N__40611),
            .in1(N__50353),
            .in2(N__40593),
            .in3(N__48985),
            .lcout(),
            .ltout(n2343_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_LC_14_18_1.C_ON=1'b0;
    defparam i24_4_lut_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_14_18_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i24_4_lut_LC_14_18_1 (
            .in0(N__40563),
            .in1(N__42918),
            .in2(N__40557),
            .in3(N__47034),
            .lcout(n53_adj_769),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_LC_14_18_4.C_ON=1'b0;
    defparam i14_4_lut_LC_14_18_4.SEQ_MODE=4'b0000;
    defparam i14_4_lut_LC_14_18_4.LUT_INIT=16'b1110111011101010;
    LogicCell40 i14_4_lut_LC_14_18_4 (
            .in0(N__40554),
            .in1(N__40548),
            .in2(N__48197),
            .in3(N__47798),
            .lcout(n43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_235_LC_14_18_6.C_ON=1'b0;
    defparam i1_4_lut_adj_235_LC_14_18_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_235_LC_14_18_6.LUT_INIT=16'b1111000011100000;
    LogicCell40 i1_4_lut_adj_235_LC_14_18_6 (
            .in0(N__42765),
            .in1(N__50352),
            .in2(N__40986),
            .in3(N__48984),
            .lcout(n2361),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_237_LC_14_19_0.C_ON=1'b0;
    defparam i4_4_lut_adj_237_LC_14_19_0.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_237_LC_14_19_0.LUT_INIT=16'b1111111111100000;
    LogicCell40 i4_4_lut_adj_237_LC_14_19_0 (
            .in0(N__42927),
            .in1(N__47799),
            .in2(N__40518),
            .in3(N__40485),
            .lcout(n33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_0__bdd_4_lut_9624_LC_14_19_1.C_ON=1'b0;
    defparam current_pin_0__bdd_4_lut_9624_LC_14_19_1.SEQ_MODE=4'b0000;
    defparam current_pin_0__bdd_4_lut_9624_LC_14_19_1.LUT_INIT=16'b1011110010110000;
    LogicCell40 current_pin_0__bdd_4_lut_9624_LC_14_19_1 (
            .in0(N__40928),
            .in1(N__50333),
            .in2(N__49040),
            .in3(N__42807),
            .lcout(),
            .ltout(n13474_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13474_bdd_4_lut_LC_14_19_2.C_ON=1'b0;
    defparam n13474_bdd_4_lut_LC_14_19_2.SEQ_MODE=4'b0000;
    defparam n13474_bdd_4_lut_LC_14_19_2.LUT_INIT=16'b1110010111100000;
    LogicCell40 n13474_bdd_4_lut_LC_14_19_2 (
            .in0(N__50334),
            .in1(N__40953),
            .in2(N__40989),
            .in3(N__40985),
            .lcout(n13477),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_236_LC_14_19_4.C_ON=1'b0;
    defparam i1_4_lut_adj_236_LC_14_19_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_236_LC_14_19_4.LUT_INIT=16'b1100100011001100;
    LogicCell40 i1_4_lut_adj_236_LC_14_19_4 (
            .in0(N__50335),
            .in1(N__40952),
            .in2(N__42768),
            .in3(N__49014),
            .lcout(n2367),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i446_4_lut_LC_14_19_5.C_ON=1'b0;
    defparam i446_4_lut_LC_14_19_5.SEQ_MODE=4'b0000;
    defparam i446_4_lut_LC_14_19_5.LUT_INIT=16'b1011000011110000;
    LogicCell40 i446_4_lut_LC_14_19_5 (
            .in0(N__42766),
            .in1(N__50336),
            .in2(N__40932),
            .in3(N__49015),
            .lcout(),
            .ltout(n2379_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i23_4_lut_LC_14_19_6.C_ON=1'b0;
    defparam i23_4_lut_LC_14_19_6.SEQ_MODE=4'b0000;
    defparam i23_4_lut_LC_14_19_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i23_4_lut_LC_14_19_6 (
            .in0(N__40911),
            .in1(N__40905),
            .in2(N__40899),
            .in3(N__40896),
            .lcout(n52_adj_770),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_209_LC_14_20_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_209_LC_14_20_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_209_LC_14_20_0.LUT_INIT=16'b1110111000000000;
    LogicCell40 i1_2_lut_3_lut_adj_209_LC_14_20_0 (
            .in0(N__49985),
            .in1(N__49775),
            .in2(_gnd_net_),
            .in3(N__40887),
            .lcout(n22_adj_732),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_219_LC_14_20_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_219_LC_14_20_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_219_LC_14_20_1.LUT_INIT=16'b0000000010001000;
    LogicCell40 i1_2_lut_3_lut_adj_219_LC_14_20_1 (
            .in0(N__49774),
            .in1(N__49984),
            .in2(_gnd_net_),
            .in3(N__49553),
            .lcout(n7232),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i26_4_lut_LC_14_20_4.C_ON=1'b0;
    defparam i26_4_lut_LC_14_20_4.SEQ_MODE=4'b0000;
    defparam i26_4_lut_LC_14_20_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i26_4_lut_LC_14_20_4 (
            .in0(N__47727),
            .in1(N__40773),
            .in2(N__43332),
            .in3(N__40764),
            .lcout(n55_adj_767),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_201_LC_14_20_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_201_LC_14_20_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_201_LC_14_20_5.LUT_INIT=16'b1010100010101000;
    LogicCell40 i1_2_lut_3_lut_adj_201_LC_14_20_5 (
            .in0(N__40755),
            .in1(N__49986),
            .in2(N__49811),
            .in3(_gnd_net_),
            .lcout(n22_adj_728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_212_LC_14_20_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_212_LC_14_20_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_212_LC_14_20_6.LUT_INIT=16'b1111101111111111;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_212_LC_14_20_6 (
            .in0(N__47265),
            .in1(N__50755),
            .in2(N__48702),
            .in3(N__50556),
            .lcout(n7145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_2_lut_LC_14_21_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_2_lut_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_2_lut_LC_14_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_2_lut_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__41283),
            .in2(_gnd_net_),
            .in3(N__41211),
            .lcout(\nx.n2477 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\nx.n10727 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_3_lut_LC_14_21_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_3_lut_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_3_lut_LC_14_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_3_lut_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41204),
            .in3(N__41157),
            .lcout(\nx.n2476 ),
            .ltout(),
            .carryin(\nx.n10727 ),
            .carryout(\nx.n10728 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_4_lut_LC_14_21_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_4_lut_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_4_lut_LC_14_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_4_lut_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__45444),
            .in2(N__41146),
            .in3(N__41112),
            .lcout(\nx.n2475 ),
            .ltout(),
            .carryin(\nx.n10728 ),
            .carryout(\nx.n10729 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_5_lut_LC_14_21_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_5_lut_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_5_lut_LC_14_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_5_lut_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__45447),
            .in2(N__41108),
            .in3(N__41079),
            .lcout(\nx.n2474 ),
            .ltout(),
            .carryin(\nx.n10729 ),
            .carryout(\nx.n10730 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_6_lut_LC_14_21_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_6_lut_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_6_lut_LC_14_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_6_lut_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__45445),
            .in2(N__43595),
            .in3(N__41064),
            .lcout(\nx.n2473 ),
            .ltout(),
            .carryin(\nx.n10730 ),
            .carryout(\nx.n10731 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_7_lut_LC_14_21_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_7_lut_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_7_lut_LC_14_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_7_lut_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__45448),
            .in2(N__41059),
            .in3(N__41016),
            .lcout(\nx.n2472 ),
            .ltout(),
            .carryin(\nx.n10731 ),
            .carryout(\nx.n10732 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_8_lut_LC_14_21_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_8_lut_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_8_lut_LC_14_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_8_lut_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__45446),
            .in2(N__41013),
            .in3(N__40992),
            .lcout(\nx.n2471 ),
            .ltout(),
            .carryin(\nx.n10732 ),
            .carryout(\nx.n10733 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_9_lut_LC_14_21_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_9_lut_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_9_lut_LC_14_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_9_lut_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__45449),
            .in2(N__43667),
            .in3(N__41445),
            .lcout(\nx.n2470 ),
            .ltout(),
            .carryin(\nx.n10733 ),
            .carryout(\nx.n10734 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_10_lut_LC_14_22_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_10_lut_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_10_lut_LC_14_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_10_lut_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(N__43616),
            .in2(N__45732),
            .in3(N__41430),
            .lcout(\nx.n2469 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\nx.n10735 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_11_lut_LC_14_22_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_11_lut_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_11_lut_LC_14_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_11_lut_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(N__45584),
            .in2(N__41422),
            .in3(N__41388),
            .lcout(\nx.n2468 ),
            .ltout(),
            .carryin(\nx.n10735 ),
            .carryout(\nx.n10736 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_12_lut_LC_14_22_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_12_lut_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_12_lut_LC_14_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_12_lut_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(N__45588),
            .in2(N__43688),
            .in3(N__41370),
            .lcout(\nx.n2467 ),
            .ltout(),
            .carryin(\nx.n10736 ),
            .carryout(\nx.n10737 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_13_lut_LC_14_22_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_13_lut_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_13_lut_LC_14_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_13_lut_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(N__45585),
            .in2(N__41367),
            .in3(N__41337),
            .lcout(\nx.n2466 ),
            .ltout(),
            .carryin(\nx.n10737 ),
            .carryout(\nx.n10738 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_14_lut_LC_14_22_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_14_lut_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_14_lut_LC_14_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_14_lut_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__45589),
            .in2(N__43228),
            .in3(N__41319),
            .lcout(\nx.n2465 ),
            .ltout(),
            .carryin(\nx.n10738 ),
            .carryout(\nx.n10739 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_15_lut_LC_14_22_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_15_lut_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_15_lut_LC_14_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_15_lut_LC_14_22_5  (
            .in0(_gnd_net_),
            .in1(N__45586),
            .in2(N__43198),
            .in3(N__41304),
            .lcout(\nx.n2464 ),
            .ltout(),
            .carryin(\nx.n10739 ),
            .carryout(\nx.n10740 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_16_lut_LC_14_22_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_16_lut_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_16_lut_LC_14_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_16_lut_LC_14_22_6  (
            .in0(_gnd_net_),
            .in1(N__45590),
            .in2(N__41882),
            .in3(N__41286),
            .lcout(\nx.n2463 ),
            .ltout(),
            .carryin(\nx.n10740 ),
            .carryout(\nx.n10741 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_17_lut_LC_14_22_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_17_lut_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_17_lut_LC_14_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_17_lut_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(N__45587),
            .in2(N__41847),
            .in3(N__41814),
            .lcout(\nx.n2462 ),
            .ltout(),
            .carryin(\nx.n10741 ),
            .carryout(\nx.n10742 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_18_lut_LC_14_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_18_lut_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_18_lut_LC_14_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_18_lut_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__45576),
            .in2(N__41811),
            .in3(N__41775),
            .lcout(\nx.n2461 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\nx.n10743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_19_lut_LC_14_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_19_lut_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_19_lut_LC_14_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_19_lut_LC_14_23_1  (
            .in0(_gnd_net_),
            .in1(N__45578),
            .in2(N__41772),
            .in3(N__41733),
            .lcout(\nx.n2460 ),
            .ltout(),
            .carryin(\nx.n10743 ),
            .carryout(\nx.n10744 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_20_lut_LC_14_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_20_lut_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_20_lut_LC_14_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_20_lut_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(N__45577),
            .in2(N__41730),
            .in3(N__41688),
            .lcout(\nx.n2459 ),
            .ltout(),
            .carryin(\nx.n10744 ),
            .carryout(\nx.n10745 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_21_lut_LC_14_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_21_lut_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_21_lut_LC_14_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_21_lut_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(N__45579),
            .in2(N__41473),
            .in3(N__41673),
            .lcout(\nx.n2458 ),
            .ltout(),
            .carryin(\nx.n10745 ),
            .carryout(\nx.n10746 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_22_lut_LC_14_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_add_1674_22_lut_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_22_lut_LC_14_23_4 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1674_22_lut_LC_14_23_4  (
            .in0(N__45580),
            .in1(N__44006),
            .in2(N__41670),
            .in3(N__41541),
            .lcout(\nx.n2489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1557_3_lut_LC_14_23_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1557_3_lut_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1557_3_lut_LC_14_23_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1557_3_lut_LC_14_23_5  (
            .in0(_gnd_net_),
            .in1(N__41514),
            .in2(N__41487),
            .in3(N__41973),
            .lcout(\nx.n2306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1610_3_lut_LC_14_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1610_3_lut_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1610_3_lut_LC_14_23_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1610_3_lut_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(N__45777),
            .in2(N__45806),
            .in3(N__44098),
            .lcout(\nx.n2391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1554_3_lut_LC_14_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1554_3_lut_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1554_3_lut_LC_14_23_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1554_3_lut_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__42222),
            .in2(N__42213),
            .in3(N__41972),
            .lcout(\nx.n2303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1548_3_lut_LC_14_24_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1548_3_lut_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1548_3_lut_LC_14_24_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1548_3_lut_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(N__42189),
            .in2(N__41991),
            .in3(N__42183),
            .lcout(\nx.n2297 ),
            .ltout(\nx.n2297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_52_LC_14_24_2 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_52_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_52_LC_14_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_52_LC_14_24_2  (
            .in0(N__46039),
            .in1(N__43726),
            .in2(N__42156),
            .in3(N__42153),
            .lcout(\nx.n31_adj_645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1552_3_lut_LC_14_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1552_3_lut_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1552_3_lut_LC_14_24_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1552_3_lut_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(N__42135),
            .in2(N__41990),
            .in3(N__42128),
            .lcout(\nx.n2301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1550_3_lut_LC_14_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1550_3_lut_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1550_3_lut_LC_14_24_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1550_3_lut_LC_14_24_4  (
            .in0(_gnd_net_),
            .in1(N__42099),
            .in2(N__42093),
            .in3(N__41981),
            .lcout(\nx.n2299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1549_3_lut_LC_14_24_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1549_3_lut_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1549_3_lut_LC_14_24_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1549_3_lut_LC_14_24_5  (
            .in0(N__42063),
            .in1(_gnd_net_),
            .in2(N__41989),
            .in3(N__42057),
            .lcout(\nx.n2298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1543_3_lut_LC_14_24_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1543_3_lut_LC_14_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1543_3_lut_LC_14_24_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1543_3_lut_LC_14_24_6  (
            .in0(_gnd_net_),
            .in1(N__42030),
            .in2(N__42024),
            .in3(N__41977),
            .lcout(\nx.n2292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1615_3_lut_LC_14_24_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1615_3_lut_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1615_3_lut_LC_14_24_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1615_3_lut_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(N__45990),
            .in2(N__46008),
            .in3(N__44099),
            .lcout(\nx.n2396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9330_4_lut_LC_14_28_3.C_ON=1'b0;
    defparam i9330_4_lut_LC_14_28_3.SEQ_MODE=4'b0000;
    defparam i9330_4_lut_LC_14_28_3.LUT_INIT=16'b1111100011101100;
    LogicCell40 i9330_4_lut_LC_14_28_3 (
            .in0(N__46218),
            .in1(N__46238),
            .in2(N__46278),
            .in3(N__46257),
            .lcout(),
            .ltout(n13177_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9331_3_lut_LC_14_28_4.C_ON=1'b0;
    defparam i9331_3_lut_LC_14_28_4.SEQ_MODE=4'b0000;
    defparam i9331_3_lut_LC_14_28_4.LUT_INIT=16'b0000111101010101;
    LogicCell40 i9331_3_lut_LC_14_28_4 (
            .in0(N__42333),
            .in1(_gnd_net_),
            .in2(N__42354),
            .in3(N__46353),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9329_4_lut_LC_14_28_6.C_ON=1'b0;
    defparam i9329_4_lut_LC_14_28_6.SEQ_MODE=4'b0000;
    defparam i9329_4_lut_LC_14_28_6.LUT_INIT=16'b1011101100100000;
    LogicCell40 i9329_4_lut_LC_14_28_6 (
            .in0(N__46256),
            .in1(N__46217),
            .in2(N__46239),
            .in3(N__46274),
            .lcout(n13176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_173_LC_15_15_1.C_ON=1'b0;
    defparam i1_4_lut_adj_173_LC_15_15_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_173_LC_15_15_1.LUT_INIT=16'b0010001000101010;
    LogicCell40 i1_4_lut_adj_173_LC_15_15_1 (
            .in0(N__47524),
            .in1(N__42303),
            .in2(N__42641),
            .in3(N__43319),
            .lcout(n7298),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2952_3_lut_4_lut_LC_15_15_2.C_ON=1'b0;
    defparam i2952_3_lut_4_lut_LC_15_15_2.SEQ_MODE=4'b0000;
    defparam i2952_3_lut_4_lut_LC_15_15_2.LUT_INIT=16'b1111111000000000;
    LogicCell40 i2952_3_lut_4_lut_LC_15_15_2 (
            .in0(N__46669),
            .in1(N__42325),
            .in2(N__42263),
            .in3(N__46871),
            .lcout(n6172),
            .ltout(n6172_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i12_LC_15_15_3.C_ON=1'b0;
    defparam pin_output_i0_i12_LC_15_15_3.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i12_LC_15_15_3.LUT_INIT=16'b0100010011100100;
    LogicCell40 pin_output_i0_i12_LC_15_15_3 (
            .in0(N__42297),
            .in1(N__48028),
            .in2(N__42291),
            .in3(N__46487),
            .lcout(pin_out_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48434),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_175_LC_15_15_4.C_ON=1'b0;
    defparam i1_4_lut_adj_175_LC_15_15_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_175_LC_15_15_4.LUT_INIT=16'b0010101000001010;
    LogicCell40 i1_4_lut_adj_175_LC_15_15_4 (
            .in0(N__47525),
            .in1(N__50342),
            .in2(N__42288),
            .in3(N__48096),
            .lcout(n7302),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2956_3_lut_4_lut_LC_15_15_5.C_ON=1'b0;
    defparam i2956_3_lut_4_lut_LC_15_15_5.SEQ_MODE=4'b0000;
    defparam i2956_3_lut_4_lut_LC_15_15_5.LUT_INIT=16'b1111000011010000;
    LogicCell40 i2956_3_lut_4_lut_LC_15_15_5 (
            .in0(N__50129),
            .in1(N__42256),
            .in2(N__46927),
            .in3(N__46670),
            .lcout(n6176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_181_LC_15_16_0.C_ON=1'b0;
    defparam i1_4_lut_adj_181_LC_15_16_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_181_LC_15_16_0.LUT_INIT=16'b0010001000101010;
    LogicCell40 i1_4_lut_adj_181_LC_15_16_0 (
            .in0(N__47519),
            .in1(N__46592),
            .in2(N__42633),
            .in3(N__42974),
            .lcout(n7314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_177_LC_15_16_1.C_ON=1'b0;
    defparam i1_4_lut_adj_177_LC_15_16_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_177_LC_15_16_1.LUT_INIT=16'b0000010011001100;
    LogicCell40 i1_4_lut_adj_177_LC_15_16_1 (
            .in0(N__43318),
            .in1(N__47523),
            .in2(N__47997),
            .in3(N__42518),
            .lcout(),
            .ltout(n7306_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i14_LC_15_16_2.C_ON=1'b0;
    defparam pin_output_i0_i14_LC_15_16_2.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i14_LC_15_16_2.LUT_INIT=16'b0000110010101100;
    LogicCell40 pin_output_i0_i14_LC_15_16_2 (
            .in0(N__42519),
            .in1(N__47839),
            .in2(N__42510),
            .in3(N__46482),
            .lcout(pin_out_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48430),
            .ce(),
            .sr(_gnd_net_));
    defparam i9314_3_lut_LC_15_16_3.C_ON=1'b0;
    defparam i9314_3_lut_LC_15_16_3.SEQ_MODE=4'b0000;
    defparam i9314_3_lut_LC_15_16_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i9314_3_lut_LC_15_16_3 (
            .in0(N__42487),
            .in1(N__42400),
            .in2(_gnd_net_),
            .in3(N__48995),
            .lcout(),
            .ltout(n13161_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13468_bdd_4_lut_LC_15_16_4.C_ON=1'b0;
    defparam n13468_bdd_4_lut_LC_15_16_4.SEQ_MODE=4'b0000;
    defparam n13468_bdd_4_lut_LC_15_16_4.LUT_INIT=16'b1110111001010000;
    LogicCell40 n13468_bdd_4_lut_LC_15_16_4 (
            .in0(N__50565),
            .in1(N__42471),
            .in2(N__42459),
            .in3(N__48006),
            .lcout(n13471),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_165_LC_15_16_6.C_ON=1'b0;
    defparam i1_4_lut_adj_165_LC_15_16_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_165_LC_15_16_6.LUT_INIT=16'b0011000001110000;
    LogicCell40 i1_4_lut_adj_165_LC_15_16_6 (
            .in0(N__42454),
            .in1(N__42425),
            .in2(N__47534),
            .in3(N__42625),
            .lcout(),
            .ltout(n7282_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i8_LC_15_16_7.C_ON=1'b0;
    defparam pin_output_i0_i8_LC_15_16_7.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i8_LC_15_16_7.LUT_INIT=16'b0100111101000000;
    LogicCell40 pin_output_i0_i8_LC_15_16_7 (
            .in0(N__46481),
            .in1(N__42426),
            .in2(N__42414),
            .in3(N__42401),
            .lcout(pin_out_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48430),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_186_LC_15_17_2.C_ON=1'b0;
    defparam i1_4_lut_adj_186_LC_15_17_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_186_LC_15_17_2.LUT_INIT=16'b0000101000101010;
    LogicCell40 i1_4_lut_adj_186_LC_15_17_2 (
            .in0(N__47506),
            .in1(N__47996),
            .in2(N__42387),
            .in3(N__42972),
            .lcout(),
            .ltout(n7322_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i18_LC_15_17_3.C_ON=1'b0;
    defparam pin_output_i0_i18_LC_15_17_3.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i18_LC_15_17_3.LUT_INIT=16'b0000110010101100;
    LogicCell40 pin_output_i0_i18_LC_15_17_3 (
            .in0(N__42386),
            .in1(N__42538),
            .in2(N__42372),
            .in3(N__46483),
            .lcout(pin_out_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48424),
            .ce(),
            .sr(_gnd_net_));
    defparam i9513_3_lut_LC_15_17_4.C_ON=1'b0;
    defparam i9513_3_lut_LC_15_17_4.SEQ_MODE=4'b0000;
    defparam i9513_3_lut_LC_15_17_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 i9513_3_lut_LC_15_17_4 (
            .in0(N__42369),
            .in1(N__50713),
            .in2(_gnd_net_),
            .in3(N__42363),
            .lcout(n13362),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_276_i8_2_lut_3_lut_LC_15_17_6.C_ON=1'b0;
    defparam equal_276_i8_2_lut_3_lut_LC_15_17_6.SEQ_MODE=4'b0000;
    defparam equal_276_i8_2_lut_3_lut_LC_15_17_6.LUT_INIT=16'b1011101111111111;
    LogicCell40 equal_276_i8_2_lut_3_lut_LC_15_17_6 (
            .in0(N__48680),
            .in1(N__50714),
            .in2(_gnd_net_),
            .in3(N__50535),
            .lcout(n8_adj_747),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_15_17_7.C_ON=1'b0;
    defparam i2_4_lut_LC_15_17_7.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_15_17_7.LUT_INIT=16'b1100110011000100;
    LogicCell40 i2_4_lut_LC_15_17_7 (
            .in0(N__50130),
            .in1(N__47271),
            .in2(N__46692),
            .in3(N__46777),
            .lcout(n12135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i20_LC_15_18_0.C_ON=1'b0;
    defparam pin_output_i0_i20_LC_15_18_0.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i20_LC_15_18_0.LUT_INIT=16'b0101000011011000;
    LogicCell40 pin_output_i0_i20_LC_15_18_0 (
            .in0(N__42561),
            .in1(N__42575),
            .in2(N__42863),
            .in3(N__46450),
            .lcout(pin_out_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48431),
            .ce(),
            .sr(_gnd_net_));
    defparam i452_3_lut_4_lut_LC_15_18_1.C_ON=1'b0;
    defparam i452_3_lut_4_lut_LC_15_18_1.SEQ_MODE=4'b0000;
    defparam i452_3_lut_4_lut_LC_15_18_1.LUT_INIT=16'b1111000011100000;
    LogicCell40 i452_3_lut_4_lut_LC_15_18_1 (
            .in0(N__42830),
            .in1(N__42609),
            .in2(N__49233),
            .in3(N__49123),
            .lcout(n2385),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i440_3_lut_LC_15_18_2.C_ON=1'b0;
    defparam i440_3_lut_LC_15_18_2.SEQ_MODE=4'b0000;
    defparam i440_3_lut_LC_15_18_2.LUT_INIT=16'b1100110010001000;
    LogicCell40 i440_3_lut_LC_15_18_2 (
            .in0(N__47993),
            .in1(N__42800),
            .in2(_gnd_net_),
            .in3(N__42767),
            .lcout(n2373),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i16_LC_15_18_4.C_ON=1'b0;
    defparam pin_output_i0_i16_LC_15_18_4.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i16_LC_15_18_4.LUT_INIT=16'b0100010011100100;
    LogicCell40 pin_output_i0_i16_LC_15_18_4 (
            .in0(N__42735),
            .in1(N__43085),
            .in2(N__46602),
            .in3(N__46448),
            .lcout(pin_out_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48431),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_184_LC_15_18_5.C_ON=1'b0;
    defparam i1_4_lut_adj_184_LC_15_18_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_184_LC_15_18_5.LUT_INIT=16'b0100010001001100;
    LogicCell40 i1_4_lut_adj_184_LC_15_18_5 (
            .in0(N__42665),
            .in1(N__47494),
            .in2(N__42725),
            .in3(N__42973),
            .lcout(),
            .ltout(n7318_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i17_LC_15_18_6.C_ON=1'b0;
    defparam pin_output_i0_i17_LC_15_18_6.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i17_LC_15_18_6.LUT_INIT=16'b0000101011001010;
    LogicCell40 pin_output_i0_i17_LC_15_18_6 (
            .in0(N__43048),
            .in1(N__42666),
            .in2(N__42648),
            .in3(N__46449),
            .lcout(pin_out_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48431),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_193_LC_15_18_7.C_ON=1'b0;
    defparam i1_4_lut_adj_193_LC_15_18_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_193_LC_15_18_7.LUT_INIT=16'b0001111100000000;
    LogicCell40 i1_4_lut_adj_193_LC_15_18_7 (
            .in0(N__47298),
            .in1(N__42610),
            .in2(N__42576),
            .in3(N__47493),
            .lcout(n7330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_0__bdd_4_lut_9596_LC_15_19_1.C_ON=1'b0;
    defparam current_pin_0__bdd_4_lut_9596_LC_15_19_1.SEQ_MODE=4'b0000;
    defparam current_pin_0__bdd_4_lut_9596_LC_15_19_1.LUT_INIT=16'b1110001011001100;
    LogicCell40 current_pin_0__bdd_4_lut_9596_LC_15_19_1 (
            .in0(N__42542),
            .in1(N__49000),
            .in2(N__42998),
            .in3(N__50346),
            .lcout(),
            .ltout(n13438_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13438_bdd_4_lut_LC_15_19_2.C_ON=1'b0;
    defparam n13438_bdd_4_lut_LC_15_19_2.SEQ_MODE=4'b0000;
    defparam n13438_bdd_4_lut_LC_15_19_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n13438_bdd_4_lut_LC_15_19_2 (
            .in0(N__50347),
            .in1(N__43084),
            .in2(N__43068),
            .in3(N__43052),
            .lcout(),
            .ltout(n13441_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9295_3_lut_LC_15_19_3.C_ON=1'b0;
    defparam i9295_3_lut_LC_15_19_3.SEQ_MODE=4'b0000;
    defparam i9295_3_lut_LC_15_19_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 i9295_3_lut_LC_15_19_3 (
            .in0(_gnd_net_),
            .in1(N__43338),
            .in2(N__43029),
            .in3(N__50536),
            .lcout(),
            .ltout(n13142_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9514_4_lut_LC_15_19_4.C_ON=1'b0;
    defparam i9514_4_lut_LC_15_19_4.SEQ_MODE=4'b0000;
    defparam i9514_4_lut_LC_15_19_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 i9514_4_lut_LC_15_19_4 (
            .in0(N__48681),
            .in1(N__50759),
            .in2(N__43026),
            .in3(N__43023),
            .lcout(n149),
            .ltout(n149_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i19_LC_15_19_5.C_ON=1'b0;
    defparam pin_output_i0_i19_LC_15_19_5.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i19_LC_15_19_5.LUT_INIT=16'b0000110010101010;
    LogicCell40 pin_output_i0_i19_LC_15_19_5 (
            .in0(N__42994),
            .in1(N__42948),
            .in2(N__43014),
            .in3(N__42933),
            .lcout(pin_out_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48435),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_190_LC_15_19_7.C_ON=1'b0;
    defparam i1_4_lut_adj_190_LC_15_19_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_190_LC_15_19_7.LUT_INIT=16'b0100000011110000;
    LogicCell40 i1_4_lut_adj_190_LC_15_19_7 (
            .in0(N__42978),
            .in1(N__43289),
            .in2(N__47527),
            .in3(N__42947),
            .lcout(n7326),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_887_i11_2_lut_4_lut_LC_15_20_0.C_ON=1'b0;
    defparam equal_887_i11_2_lut_4_lut_LC_15_20_0.SEQ_MODE=4'b0000;
    defparam equal_887_i11_2_lut_4_lut_LC_15_20_0.LUT_INIT=16'b1111111111111011;
    LogicCell40 equal_887_i11_2_lut_4_lut_LC_15_20_0 (
            .in0(N__50345),
            .in1(N__48999),
            .in2(N__50567),
            .in3(N__50761),
            .lcout(n11_adj_734),
            .ltout(n11_adj_734_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_241_LC_15_20_1.C_ON=1'b0;
    defparam i7_4_lut_adj_241_LC_15_20_1.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_241_LC_15_20_1.LUT_INIT=16'b1111111110101000;
    LogicCell40 i7_4_lut_adj_241_LC_15_20_1 (
            .in0(N__49191),
            .in1(N__49141),
            .in2(N__42921),
            .in3(N__46992),
            .lcout(n36_adj_773),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Mux_35_i19_3_lut_LC_15_20_4.C_ON=1'b0;
    defparam Mux_35_i19_3_lut_LC_15_20_4.SEQ_MODE=4'b0000;
    defparam Mux_35_i19_3_lut_LC_15_20_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 Mux_35_i19_3_lut_LC_15_20_4 (
            .in0(N__42898),
            .in1(N__42856),
            .in2(_gnd_net_),
            .in3(N__48996),
            .lcout(),
            .ltout(n19_adj_735_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9294_4_lut_LC_15_20_5.C_ON=1'b0;
    defparam i9294_4_lut_LC_15_20_5.SEQ_MODE=4'b0000;
    defparam i9294_4_lut_LC_15_20_5.LUT_INIT=16'b0100010011110000;
    LogicCell40 i9294_4_lut_LC_15_20_5 (
            .in0(N__48997),
            .in1(N__47323),
            .in2(N__43341),
            .in3(N__50343),
            .lcout(n13141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_783_i11_2_lut_4_lut_LC_15_20_6.C_ON=1'b0;
    defparam equal_783_i11_2_lut_4_lut_LC_15_20_6.SEQ_MODE=4'b0000;
    defparam equal_783_i11_2_lut_4_lut_LC_15_20_6.LUT_INIT=16'b1111111111101111;
    LogicCell40 equal_783_i11_2_lut_4_lut_LC_15_20_6 (
            .in0(N__50344),
            .in1(N__48998),
            .in2(N__50566),
            .in3(N__50760),
            .lcout(n11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_183_LC_15_20_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_183_LC_15_20_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_183_LC_15_20_7.LUT_INIT=16'b1110111000000000;
    LogicCell40 i1_2_lut_3_lut_adj_183_LC_15_20_7 (
            .in0(N__49923),
            .in1(N__49722),
            .in2(_gnd_net_),
            .in3(N__49516),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_179_LC_15_21_4.C_ON=1'b0;
    defparam i1_4_lut_adj_179_LC_15_21_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_179_LC_15_21_4.LUT_INIT=16'b0010000010101010;
    LogicCell40 i1_4_lut_adj_179_LC_15_21_4 (
            .in0(N__47518),
            .in1(N__43323),
            .in2(N__43299),
            .in3(N__43250),
            .lcout(),
            .ltout(n7310_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i15_LC_15_21_5.C_ON=1'b0;
    defparam pin_output_i0_i15_LC_15_21_5.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i15_LC_15_21_5.LUT_INIT=16'b0000110010101100;
    LogicCell40 pin_output_i0_i15_LC_15_21_5 (
            .in0(N__43251),
            .in1(N__47869),
            .in2(N__43236),
            .in3(N__46488),
            .lcout(pin_out_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48440),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i14_LC_15_21_7.C_ON=1'b0;
    defparam neopxl_color_i14_LC_15_21_7.SEQ_MODE=4'b1000;
    defparam neopxl_color_i14_LC_15_21_7.LUT_INIT=16'b1011111100000010;
    LogicCell40 neopxl_color_i14_LC_15_21_7 (
            .in0(N__49554),
            .in1(N__49956),
            .in2(N__49757),
            .in3(N__43149),
            .lcout(neopxl_color_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48440),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1617_3_lut_LC_15_22_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1617_3_lut_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1617_3_lut_LC_15_22_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i1617_3_lut_LC_15_22_1  (
            .in0(N__44113),
            .in1(_gnd_net_),
            .in2(N__43737),
            .in3(N__43710),
            .lcout(\nx.n2398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1616_3_lut_LC_15_22_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1616_3_lut_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1616_3_lut_LC_15_22_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1616_3_lut_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__46047),
            .in2(N__46023),
            .in3(N__44109),
            .lcout(\nx.n2397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i14_LC_15_22_3.C_ON=1'b0;
    defparam neopxl_color_prev_i14_LC_15_22_3.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i14_LC_15_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 neopxl_color_prev_i14_LC_15_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43159),
            .lcout(neopxl_color_prev_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48444),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1619_3_lut_LC_15_22_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1619_3_lut_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1619_3_lut_LC_15_22_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1619_3_lut_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__43785),
            .in2(N__43815),
            .in3(N__44115),
            .lcout(\nx.n2400 ),
            .ltout(\nx.n2400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_62_LC_15_22_5 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_62_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_62_LC_15_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_62_LC_15_22_5  (
            .in0(N__43591),
            .in1(N__43615),
            .in2(N__43671),
            .in3(N__43668),
            .lcout(\nx.n35_adj_658 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1621_3_lut_LC_15_22_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1621_3_lut_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1621_3_lut_LC_15_22_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \nx.mod_5_i1621_3_lut_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__44114),
            .in2(N__43872),
            .in3(N__43894),
            .lcout(\nx.n2402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1625_rep_47_3_lut_LC_15_22_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1625_rep_47_3_lut_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1625_rep_47_3_lut_LC_15_22_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1625_rep_47_3_lut_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(N__43380),
            .in2(N__44128),
            .in3(N__43410),
            .lcout(\nx.n2406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_2_lut_LC_15_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_2_lut_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_2_lut_LC_15_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_2_lut_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__43572),
            .in2(_gnd_net_),
            .in3(N__43497),
            .lcout(\nx.n2377 ),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\nx.n10708 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_3_lut_LC_15_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_3_lut_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_3_lut_LC_15_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_3_lut_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43494),
            .in3(N__43455),
            .lcout(\nx.n2376 ),
            .ltout(),
            .carryin(\nx.n10708 ),
            .carryout(\nx.n10709 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_4_lut_LC_15_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_4_lut_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_4_lut_LC_15_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_4_lut_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__45677),
            .in2(N__43452),
            .in3(N__43413),
            .lcout(\nx.n2375 ),
            .ltout(),
            .carryin(\nx.n10709 ),
            .carryout(\nx.n10710 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_5_lut_LC_15_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_5_lut_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_5_lut_LC_15_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_5_lut_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__45679),
            .in2(N__43409),
            .in3(N__43374),
            .lcout(\nx.n2374 ),
            .ltout(),
            .carryin(\nx.n10710 ),
            .carryout(\nx.n10711 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_6_lut_LC_15_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_6_lut_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_6_lut_LC_15_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_6_lut_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(N__45678),
            .in2(N__43371),
            .in3(N__43989),
            .lcout(\nx.n2373 ),
            .ltout(),
            .carryin(\nx.n10711 ),
            .carryout(\nx.n10712 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_7_lut_LC_15_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_7_lut_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_7_lut_LC_15_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_7_lut_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__45680),
            .in2(N__43985),
            .in3(N__43944),
            .lcout(\nx.n2372 ),
            .ltout(),
            .carryin(\nx.n10712 ),
            .carryout(\nx.n10713 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_8_lut_LC_15_23_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_8_lut_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_8_lut_LC_15_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_8_lut_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__43940),
            .in2(N__45756),
            .in3(N__43902),
            .lcout(\nx.n2371 ),
            .ltout(),
            .carryin(\nx.n10713 ),
            .carryout(\nx.n10714 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_9_lut_LC_15_23_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_9_lut_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_9_lut_LC_15_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_9_lut_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__45684),
            .in2(N__43898),
            .in3(N__43863),
            .lcout(\nx.n2370 ),
            .ltout(),
            .carryin(\nx.n10714 ),
            .carryout(\nx.n10715 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_10_lut_LC_15_24_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_10_lut_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_10_lut_LC_15_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_10_lut_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__45414),
            .in2(N__43860),
            .in3(N__43818),
            .lcout(\nx.n2369 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\nx.n10716 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_11_lut_LC_15_24_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_11_lut_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_11_lut_LC_15_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_11_lut_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__45433),
            .in2(N__43811),
            .in3(N__43776),
            .lcout(\nx.n2368 ),
            .ltout(),
            .carryin(\nx.n10716 ),
            .carryout(\nx.n10717 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_12_lut_LC_15_24_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_12_lut_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_12_lut_LC_15_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_12_lut_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__45415),
            .in2(N__43773),
            .in3(N__43740),
            .lcout(\nx.n2367 ),
            .ltout(),
            .carryin(\nx.n10717 ),
            .carryout(\nx.n10718 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_13_lut_LC_15_24_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_13_lut_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_13_lut_LC_15_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_13_lut_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__45434),
            .in2(N__43733),
            .in3(N__43701),
            .lcout(\nx.n2366 ),
            .ltout(),
            .carryin(\nx.n10718 ),
            .carryout(\nx.n10719 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_14_lut_LC_15_24_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_14_lut_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_14_lut_LC_15_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_14_lut_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__45416),
            .in2(N__46046),
            .in3(N__46011),
            .lcout(\nx.n2365 ),
            .ltout(),
            .carryin(\nx.n10719 ),
            .carryout(\nx.n10720 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_15_lut_LC_15_24_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_15_lut_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_15_lut_LC_15_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_15_lut_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__45435),
            .in2(N__46007),
            .in3(N__45984),
            .lcout(\nx.n2364 ),
            .ltout(),
            .carryin(\nx.n10720 ),
            .carryout(\nx.n10721 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_16_lut_LC_15_24_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_16_lut_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_16_lut_LC_15_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_16_lut_LC_15_24_6  (
            .in0(_gnd_net_),
            .in1(N__45417),
            .in2(N__45981),
            .in3(N__45948),
            .lcout(\nx.n2363 ),
            .ltout(),
            .carryin(\nx.n10721 ),
            .carryout(\nx.n10722 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_17_lut_LC_15_24_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_17_lut_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_17_lut_LC_15_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_17_lut_LC_15_24_7  (
            .in0(_gnd_net_),
            .in1(N__45436),
            .in2(N__45945),
            .in3(N__45900),
            .lcout(\nx.n2362 ),
            .ltout(),
            .carryin(\nx.n10722 ),
            .carryout(\nx.n10723 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_18_lut_LC_15_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_18_lut_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_18_lut_LC_15_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_18_lut_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(N__45411),
            .in2(N__45897),
            .in3(N__45855),
            .lcout(\nx.n2361 ),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(\nx.n10724 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_19_lut_LC_15_25_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_19_lut_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_19_lut_LC_15_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_19_lut_LC_15_25_1  (
            .in0(_gnd_net_),
            .in1(N__45432),
            .in2(N__45852),
            .in3(N__45813),
            .lcout(\nx.n2360 ),
            .ltout(),
            .carryin(\nx.n10724 ),
            .carryout(\nx.n10725 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_20_lut_LC_15_25_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_20_lut_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_20_lut_LC_15_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_20_lut_LC_15_25_2  (
            .in0(_gnd_net_),
            .in1(N__45412),
            .in2(N__45805),
            .in3(N__45768),
            .lcout(\nx.n2359 ),
            .ltout(),
            .carryin(\nx.n10725 ),
            .carryout(\nx.n10726 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_21_lut_LC_15_25_3 .C_ON=1'b0;
    defparam \nx.mod_5_add_1607_21_lut_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_21_lut_LC_15_25_3 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1607_21_lut_LC_15_25_3  (
            .in0(N__45413),
            .in1(N__44148),
            .in2(N__44130),
            .in3(N__44013),
            .lcout(\nx.n2390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i0_LC_15_26_0.C_ON=1'b1;
    defparam blink_counter_1105__i0_LC_15_26_0.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i0_LC_15_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i0_LC_15_26_0 (
            .in0(_gnd_net_),
            .in1(N__46119),
            .in2(_gnd_net_),
            .in3(N__46113),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(n10548),
            .clk(N__48450),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i1_LC_15_26_1.C_ON=1'b1;
    defparam blink_counter_1105__i1_LC_15_26_1.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i1_LC_15_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i1_LC_15_26_1 (
            .in0(_gnd_net_),
            .in1(N__46110),
            .in2(_gnd_net_),
            .in3(N__46104),
            .lcout(n25),
            .ltout(),
            .carryin(n10548),
            .carryout(n10549),
            .clk(N__48450),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i2_LC_15_26_2.C_ON=1'b1;
    defparam blink_counter_1105__i2_LC_15_26_2.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i2_LC_15_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i2_LC_15_26_2 (
            .in0(_gnd_net_),
            .in1(N__46101),
            .in2(_gnd_net_),
            .in3(N__46095),
            .lcout(n24),
            .ltout(),
            .carryin(n10549),
            .carryout(n10550),
            .clk(N__48450),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i3_LC_15_26_3.C_ON=1'b1;
    defparam blink_counter_1105__i3_LC_15_26_3.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i3_LC_15_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i3_LC_15_26_3 (
            .in0(_gnd_net_),
            .in1(N__46092),
            .in2(_gnd_net_),
            .in3(N__46086),
            .lcout(n23),
            .ltout(),
            .carryin(n10550),
            .carryout(n10551),
            .clk(N__48450),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i4_LC_15_26_4.C_ON=1'b1;
    defparam blink_counter_1105__i4_LC_15_26_4.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i4_LC_15_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i4_LC_15_26_4 (
            .in0(_gnd_net_),
            .in1(N__46083),
            .in2(_gnd_net_),
            .in3(N__46077),
            .lcout(n22),
            .ltout(),
            .carryin(n10551),
            .carryout(n10552),
            .clk(N__48450),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i5_LC_15_26_5.C_ON=1'b1;
    defparam blink_counter_1105__i5_LC_15_26_5.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i5_LC_15_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i5_LC_15_26_5 (
            .in0(_gnd_net_),
            .in1(N__46074),
            .in2(_gnd_net_),
            .in3(N__46068),
            .lcout(n21_adj_737),
            .ltout(),
            .carryin(n10552),
            .carryout(n10553),
            .clk(N__48450),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i6_LC_15_26_6.C_ON=1'b1;
    defparam blink_counter_1105__i6_LC_15_26_6.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i6_LC_15_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i6_LC_15_26_6 (
            .in0(_gnd_net_),
            .in1(N__46065),
            .in2(_gnd_net_),
            .in3(N__46059),
            .lcout(n20),
            .ltout(),
            .carryin(n10553),
            .carryout(n10554),
            .clk(N__48450),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i7_LC_15_26_7.C_ON=1'b1;
    defparam blink_counter_1105__i7_LC_15_26_7.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i7_LC_15_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i7_LC_15_26_7 (
            .in0(_gnd_net_),
            .in1(N__46056),
            .in2(_gnd_net_),
            .in3(N__46050),
            .lcout(n19_adj_718),
            .ltout(),
            .carryin(n10554),
            .carryout(n10555),
            .clk(N__48450),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i8_LC_15_27_0.C_ON=1'b1;
    defparam blink_counter_1105__i8_LC_15_27_0.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i8_LC_15_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i8_LC_15_27_0 (
            .in0(_gnd_net_),
            .in1(N__46200),
            .in2(_gnd_net_),
            .in3(N__46194),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_15_27_0_),
            .carryout(n10556),
            .clk(N__48451),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i9_LC_15_27_1.C_ON=1'b1;
    defparam blink_counter_1105__i9_LC_15_27_1.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i9_LC_15_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i9_LC_15_27_1 (
            .in0(_gnd_net_),
            .in1(N__46191),
            .in2(_gnd_net_),
            .in3(N__46185),
            .lcout(n17),
            .ltout(),
            .carryin(n10556),
            .carryout(n10557),
            .clk(N__48451),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i10_LC_15_27_2.C_ON=1'b1;
    defparam blink_counter_1105__i10_LC_15_27_2.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i10_LC_15_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i10_LC_15_27_2 (
            .in0(_gnd_net_),
            .in1(N__46182),
            .in2(_gnd_net_),
            .in3(N__46176),
            .lcout(n16),
            .ltout(),
            .carryin(n10557),
            .carryout(n10558),
            .clk(N__48451),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i11_LC_15_27_3.C_ON=1'b1;
    defparam blink_counter_1105__i11_LC_15_27_3.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i11_LC_15_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i11_LC_15_27_3 (
            .in0(_gnd_net_),
            .in1(N__46173),
            .in2(_gnd_net_),
            .in3(N__46167),
            .lcout(n15_adj_759),
            .ltout(),
            .carryin(n10558),
            .carryout(n10559),
            .clk(N__48451),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i12_LC_15_27_4.C_ON=1'b1;
    defparam blink_counter_1105__i12_LC_15_27_4.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i12_LC_15_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i12_LC_15_27_4 (
            .in0(_gnd_net_),
            .in1(N__46164),
            .in2(_gnd_net_),
            .in3(N__46158),
            .lcout(n14_adj_745),
            .ltout(),
            .carryin(n10559),
            .carryout(n10560),
            .clk(N__48451),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i13_LC_15_27_5.C_ON=1'b1;
    defparam blink_counter_1105__i13_LC_15_27_5.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i13_LC_15_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i13_LC_15_27_5 (
            .in0(_gnd_net_),
            .in1(N__46155),
            .in2(_gnd_net_),
            .in3(N__46149),
            .lcout(n13),
            .ltout(),
            .carryin(n10560),
            .carryout(n10561),
            .clk(N__48451),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i14_LC_15_27_6.C_ON=1'b1;
    defparam blink_counter_1105__i14_LC_15_27_6.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i14_LC_15_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i14_LC_15_27_6 (
            .in0(_gnd_net_),
            .in1(N__46146),
            .in2(_gnd_net_),
            .in3(N__46140),
            .lcout(n12),
            .ltout(),
            .carryin(n10561),
            .carryout(n10562),
            .clk(N__48451),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i15_LC_15_27_7.C_ON=1'b1;
    defparam blink_counter_1105__i15_LC_15_27_7.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i15_LC_15_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i15_LC_15_27_7 (
            .in0(_gnd_net_),
            .in1(N__46137),
            .in2(_gnd_net_),
            .in3(N__46131),
            .lcout(n11_adj_758),
            .ltout(),
            .carryin(n10562),
            .carryout(n10563),
            .clk(N__48451),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i16_LC_15_28_0.C_ON=1'b1;
    defparam blink_counter_1105__i16_LC_15_28_0.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i16_LC_15_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i16_LC_15_28_0 (
            .in0(_gnd_net_),
            .in1(N__46128),
            .in2(_gnd_net_),
            .in3(N__46122),
            .lcout(n10_adj_757),
            .ltout(),
            .carryin(bfn_15_28_0_),
            .carryout(n10564),
            .clk(N__48452),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i17_LC_15_28_1.C_ON=1'b1;
    defparam blink_counter_1105__i17_LC_15_28_1.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i17_LC_15_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i17_LC_15_28_1 (
            .in0(_gnd_net_),
            .in1(N__46314),
            .in2(_gnd_net_),
            .in3(N__46308),
            .lcout(n9),
            .ltout(),
            .carryin(n10564),
            .carryout(n10565),
            .clk(N__48452),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i18_LC_15_28_2.C_ON=1'b1;
    defparam blink_counter_1105__i18_LC_15_28_2.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i18_LC_15_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i18_LC_15_28_2 (
            .in0(_gnd_net_),
            .in1(N__46305),
            .in2(_gnd_net_),
            .in3(N__46299),
            .lcout(n8_adj_755),
            .ltout(),
            .carryin(n10565),
            .carryout(n10566),
            .clk(N__48452),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i19_LC_15_28_3.C_ON=1'b1;
    defparam blink_counter_1105__i19_LC_15_28_3.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i19_LC_15_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i19_LC_15_28_3 (
            .in0(_gnd_net_),
            .in1(N__46296),
            .in2(_gnd_net_),
            .in3(N__46290),
            .lcout(n7),
            .ltout(),
            .carryin(n10566),
            .carryout(n10567),
            .clk(N__48452),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i20_LC_15_28_4.C_ON=1'b1;
    defparam blink_counter_1105__i20_LC_15_28_4.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i20_LC_15_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i20_LC_15_28_4 (
            .in0(_gnd_net_),
            .in1(N__46287),
            .in2(_gnd_net_),
            .in3(N__46281),
            .lcout(n6_adj_756),
            .ltout(),
            .carryin(n10567),
            .carryout(n10568),
            .clk(N__48452),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i21_LC_15_28_5.C_ON=1'b1;
    defparam blink_counter_1105__i21_LC_15_28_5.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i21_LC_15_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i21_LC_15_28_5 (
            .in0(_gnd_net_),
            .in1(N__46273),
            .in2(_gnd_net_),
            .in3(N__46260),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n10568),
            .carryout(n10569),
            .clk(N__48452),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i22_LC_15_28_6.C_ON=1'b1;
    defparam blink_counter_1105__i22_LC_15_28_6.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i22_LC_15_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i22_LC_15_28_6 (
            .in0(_gnd_net_),
            .in1(N__46255),
            .in2(_gnd_net_),
            .in3(N__46242),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n10569),
            .carryout(n10570),
            .clk(N__48452),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i23_LC_15_28_7.C_ON=1'b1;
    defparam blink_counter_1105__i23_LC_15_28_7.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i23_LC_15_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i23_LC_15_28_7 (
            .in0(_gnd_net_),
            .in1(N__46234),
            .in2(_gnd_net_),
            .in3(N__46221),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n10570),
            .carryout(n10571),
            .clk(N__48452),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i24_LC_15_29_0.C_ON=1'b1;
    defparam blink_counter_1105__i24_LC_15_29_0.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i24_LC_15_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i24_LC_15_29_0 (
            .in0(_gnd_net_),
            .in1(N__46216),
            .in2(_gnd_net_),
            .in3(N__46203),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_15_29_0_),
            .carryout(n10572),
            .clk(N__48453),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1105__i25_LC_15_29_1.C_ON=1'b0;
    defparam blink_counter_1105__i25_LC_15_29_1.SEQ_MODE=4'b1000;
    defparam blink_counter_1105__i25_LC_15_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_1105__i25_LC_15_29_1 (
            .in0(_gnd_net_),
            .in1(N__46352),
            .in2(_gnd_net_),
            .in3(N__46356),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48453),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_1103__i0_LC_16_14_0.C_ON=1'b0;
    defparam counter_1103__i0_LC_16_14_0.SEQ_MODE=4'b1000;
    defparam counter_1103__i0_LC_16_14_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 counter_1103__i0_LC_16_14_0 (
            .in0(N__46578),
            .in1(N__49412),
            .in2(_gnd_net_),
            .in3(N__46341),
            .lcout(counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48441),
            .ce(N__47530),
            .sr(_gnd_net_));
    defparam counter_1103_add_4_2_lut_LC_16_15_0.C_ON=1'b1;
    defparam counter_1103_add_4_2_lut_LC_16_15_0.SEQ_MODE=4'b0000;
    defparam counter_1103_add_4_2_lut_LC_16_15_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_1103_add_4_2_lut_LC_16_15_0 (
            .in0(_gnd_net_),
            .in1(N__47570),
            .in2(N__47630),
            .in3(N__46335),
            .lcout(n45),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(n10510),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_1103__i1_LC_16_15_1.C_ON=1'b1;
    defparam counter_1103__i1_LC_16_15_1.SEQ_MODE=4'b1000;
    defparam counter_1103__i1_LC_16_15_1.LUT_INIT=16'b1100101000111010;
    LogicCell40 counter_1103__i1_LC_16_15_1 (
            .in0(N__46567),
            .in1(N__48177),
            .in2(N__46928),
            .in3(N__46332),
            .lcout(counter_1),
            .ltout(),
            .carryin(n10510),
            .carryout(n10511),
            .clk(N__48438),
            .ce(N__47538),
            .sr(_gnd_net_));
    defparam counter_1103__i2_LC_16_15_2.C_ON=1'b1;
    defparam counter_1103__i2_LC_16_15_2.SEQ_MODE=4'b1000;
    defparam counter_1103__i2_LC_16_15_2.LUT_INIT=16'b1110001000101110;
    LogicCell40 counter_1103__i2_LC_16_15_2 (
            .in0(N__46579),
            .in1(N__46878),
            .in2(N__47556),
            .in3(N__46329),
            .lcout(counter_2),
            .ltout(),
            .carryin(n10511),
            .carryout(n10512),
            .clk(N__48438),
            .ce(N__47538),
            .sr(_gnd_net_));
    defparam counter_1103__i3_LC_16_15_3.C_ON=1'b1;
    defparam counter_1103__i3_LC_16_15_3.SEQ_MODE=4'b1000;
    defparam counter_1103__i3_LC_16_15_3.LUT_INIT=16'b1100101000111010;
    LogicCell40 counter_1103__i3_LC_16_15_3 (
            .in0(N__46568),
            .in1(N__47598),
            .in2(N__46929),
            .in3(N__46326),
            .lcout(counter_3),
            .ltout(),
            .carryin(n10512),
            .carryout(n10513),
            .clk(N__48438),
            .ce(N__47538),
            .sr(_gnd_net_));
    defparam counter_1103__i4_LC_16_15_4.C_ON=1'b1;
    defparam counter_1103__i4_LC_16_15_4.SEQ_MODE=4'b1000;
    defparam counter_1103__i4_LC_16_15_4.LUT_INIT=16'b1110001000101110;
    LogicCell40 counter_1103__i4_LC_16_15_4 (
            .in0(N__46580),
            .in1(N__46882),
            .in2(N__47586),
            .in3(N__46323),
            .lcout(counter_4),
            .ltout(),
            .carryin(n10513),
            .carryout(n10514),
            .clk(N__48438),
            .ce(N__47538),
            .sr(_gnd_net_));
    defparam counter_1103__i5_LC_16_15_5.C_ON=1'b1;
    defparam counter_1103__i5_LC_16_15_5.SEQ_MODE=4'b1000;
    defparam counter_1103__i5_LC_16_15_5.LUT_INIT=16'b1100101000111010;
    LogicCell40 counter_1103__i5_LC_16_15_5 (
            .in0(N__46569),
            .in1(N__48162),
            .in2(N__46930),
            .in3(N__46320),
            .lcout(counter_5),
            .ltout(),
            .carryin(n10514),
            .carryout(n10515),
            .clk(N__48438),
            .ce(N__47538),
            .sr(_gnd_net_));
    defparam counter_1103__i6_LC_16_15_6.C_ON=1'b1;
    defparam counter_1103__i6_LC_16_15_6.SEQ_MODE=4'b1000;
    defparam counter_1103__i6_LC_16_15_6.LUT_INIT=16'b1110001000101110;
    LogicCell40 counter_1103__i6_LC_16_15_6 (
            .in0(N__46581),
            .in1(N__46886),
            .in2(N__47172),
            .in3(N__46317),
            .lcout(counter_6),
            .ltout(),
            .carryin(n10515),
            .carryout(n10516),
            .clk(N__48438),
            .ce(N__47538),
            .sr(_gnd_net_));
    defparam counter_1103__i7_LC_16_15_7.C_ON=1'b0;
    defparam counter_1103__i7_LC_16_15_7.SEQ_MODE=4'b1000;
    defparam counter_1103__i7_LC_16_15_7.LUT_INIT=16'b1100101000111010;
    LogicCell40 counter_1103__i7_LC_16_15_7 (
            .in0(N__46570),
            .in1(N__47229),
            .in2(N__46931),
            .in3(N__46986),
            .lcout(counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48438),
            .ce(N__47538),
            .sr(_gnd_net_));
    defparam i3_3_lut_LC_16_16_1.C_ON=1'b0;
    defparam i3_3_lut_LC_16_16_1.SEQ_MODE=4'b0000;
    defparam i3_3_lut_LC_16_16_1.LUT_INIT=16'b1111111111101110;
    LogicCell40 i3_3_lut_LC_16_16_1 (
            .in0(N__47156),
            .in1(N__49999),
            .in2(_gnd_net_),
            .in3(N__48132),
            .lcout(),
            .ltout(n8_adj_763_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9579_4_lut_LC_16_16_2.C_ON=1'b0;
    defparam i9579_4_lut_LC_16_16_2.SEQ_MODE=4'b0000;
    defparam i9579_4_lut_LC_16_16_2.LUT_INIT=16'b1010101010101011;
    LogicCell40 i9579_4_lut_LC_16_16_2 (
            .in0(N__47105),
            .in1(N__47225),
            .in2(N__46983),
            .in3(N__49526),
            .lcout(n7223),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_199_LC_16_16_4.C_ON=1'b0;
    defparam i2_3_lut_adj_199_LC_16_16_4.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_199_LC_16_16_4.LUT_INIT=16'b0000000001000100;
    LogicCell40 i2_3_lut_adj_199_LC_16_16_4 (
            .in0(N__46787),
            .in1(N__50125),
            .in2(_gnd_net_),
            .in3(N__46679),
            .lcout(n12208),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam state_7__I_0_205_i16_1_lut_LC_16_16_5.C_ON=1'b0;
    defparam state_7__I_0_205_i16_1_lut_LC_16_16_5.SEQ_MODE=4'b0000;
    defparam state_7__I_0_205_i16_1_lut_LC_16_16_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 state_7__I_0_205_i16_1_lut_LC_16_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49406),
            .lcout(current_pin_7__N_155),
            .ltout(current_pin_7__N_155_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2960_3_lut_4_lut_LC_16_16_6.C_ON=1'b0;
    defparam i2960_3_lut_4_lut_LC_16_16_6.SEQ_MODE=4'b0000;
    defparam i2960_3_lut_4_lut_LC_16_16_6.LUT_INIT=16'b1111000011100000;
    LogicCell40 i2960_3_lut_4_lut_LC_16_16_6 (
            .in0(N__46786),
            .in1(N__46744),
            .in2(N__46695),
            .in3(N__46678),
            .lcout(n6180),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_220_LC_16_16_7.C_ON=1'b0;
    defparam i2_3_lut_adj_220_LC_16_16_7.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_220_LC_16_16_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i2_3_lut_adj_220_LC_16_16_7 (
            .in0(N__49527),
            .in1(N__50000),
            .in2(_gnd_net_),
            .in3(N__49807),
            .lcout(n6971),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4169_2_lut_LC_16_17_0.C_ON=1'b0;
    defparam i4169_2_lut_LC_16_17_0.SEQ_MODE=4'b0000;
    defparam i4169_2_lut_LC_16_17_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 i4169_2_lut_LC_16_17_0 (
            .in0(_gnd_net_),
            .in1(N__49410),
            .in2(_gnd_net_),
            .in3(N__48233),
            .lcout(n7401),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4263_4_lut_LC_16_17_3.C_ON=1'b0;
    defparam i4263_4_lut_LC_16_17_3.SEQ_MODE=4'b0000;
    defparam i4263_4_lut_LC_16_17_3.LUT_INIT=16'b1011000011110100;
    LogicCell40 i4263_4_lut_LC_16_17_3 (
            .in0(N__46542),
            .in1(N__47528),
            .in2(N__47324),
            .in3(N__46475),
            .lcout(),
            .ltout(n7500_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i22_LC_16_17_4.C_ON=1'b0;
    defparam pin_output_i0_i22_LC_16_17_4.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i22_LC_16_17_4.LUT_INIT=16'b0101000001110000;
    LogicCell40 pin_output_i0_i22_LC_16_17_4 (
            .in0(N__47529),
            .in1(N__47346),
            .in2(N__47340),
            .in3(N__49411),
            .lcout(pin_out_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48427),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_233_LC_16_17_5.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_233_LC_16_17_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_233_LC_16_17_5.LUT_INIT=16'b0000111100001011;
    LogicCell40 i1_3_lut_4_lut_adj_233_LC_16_17_5 (
            .in0(N__47294),
            .in1(N__50315),
            .in2(N__49413),
            .in3(N__48955),
            .lcout(n4_adj_778),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_216_LC_16_17_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_216_LC_16_17_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_216_LC_16_17_6.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1_2_lut_3_lut_adj_216_LC_16_17_6 (
            .in0(N__48474),
            .in1(N__48519),
            .in2(_gnd_net_),
            .in3(N__48553),
            .lcout(n7142),
            .ltout(n7142_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_234_LC_16_17_7.C_ON=1'b0;
    defparam i1_2_lut_adj_234_LC_16_17_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_234_LC_16_17_7.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_234_LC_16_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47241),
            .in3(N__48645),
            .lcout(n14_adj_717),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam state__i2_LC_16_18_0.C_ON=1'b0;
    defparam state__i2_LC_16_18_0.SEQ_MODE=4'b1000;
    defparam state__i2_LC_16_18_0.LUT_INIT=16'b0011001100110010;
    LogicCell40 state__i2_LC_16_18_0 (
            .in0(N__47237),
            .in1(N__50016),
            .in2(N__47180),
            .in3(N__48150),
            .lcout(state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48436),
            .ce(N__50820),
            .sr(N__48213));
    defparam i9575_2_lut_3_lut_LC_16_18_5.C_ON=1'b0;
    defparam i9575_2_lut_3_lut_LC_16_18_5.SEQ_MODE=4'b0000;
    defparam i9575_2_lut_3_lut_LC_16_18_5.LUT_INIT=16'b0000000000010001;
    LogicCell40 i9575_2_lut_3_lut_LC_16_18_5 (
            .in0(N__50015),
            .in1(N__49751),
            .in2(_gnd_net_),
            .in3(N__49489),
            .lcout(n73),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_239_LC_16_19_0.C_ON=1'b0;
    defparam i2_4_lut_adj_239_LC_16_19_0.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_239_LC_16_19_0.LUT_INIT=16'b1111111111011111;
    LogicCell40 i2_4_lut_adj_239_LC_16_19_0 (
            .in0(N__49003),
            .in1(N__47780),
            .in2(N__50338),
            .in3(N__50611),
            .lcout(),
            .ltout(n12123_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_LC_16_19_1.C_ON=1'b0;
    defparam i19_4_lut_LC_16_19_1.SEQ_MODE=4'b0000;
    defparam i19_4_lut_LC_16_19_1.LUT_INIT=16'b1111111111101100;
    LogicCell40 i19_4_lut_LC_16_19_1 (
            .in0(N__47088),
            .in1(N__47043),
            .in2(N__47037),
            .in3(N__49056),
            .lcout(n48_adj_771),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i380_3_lut_LC_16_19_2.C_ON=1'b0;
    defparam i380_3_lut_LC_16_19_2.SEQ_MODE=4'b0000;
    defparam i380_3_lut_LC_16_19_2.LUT_INIT=16'b1010101010001000;
    LogicCell40 i380_3_lut_LC_16_19_2 (
            .in0(N__47022),
            .in1(N__47742),
            .in2(_gnd_net_),
            .in3(N__47779),
            .lcout(n2313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9297_4_lut_LC_16_19_5.C_ON=1'b0;
    defparam i9297_4_lut_LC_16_19_5.SEQ_MODE=4'b0000;
    defparam i9297_4_lut_LC_16_19_5.LUT_INIT=16'b0010001011100010;
    LogicCell40 i9297_4_lut_LC_16_19_5 (
            .in0(N__48717),
            .in1(N__50287),
            .in2(N__47927),
            .in3(N__49001),
            .lcout(),
            .ltout(n13144_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9442_4_lut_LC_16_19_6.C_ON=1'b0;
    defparam i9442_4_lut_LC_16_19_6.SEQ_MODE=4'b0000;
    defparam i9442_4_lut_LC_16_19_6.LUT_INIT=16'b0101000001000100;
    LogicCell40 i9442_4_lut_LC_16_19_6 (
            .in0(N__50752),
            .in1(N__49152),
            .in2(N__47811),
            .in3(N__50537),
            .lcout(n13279),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_791_i15_4_lut_LC_16_19_7.C_ON=1'b0;
    defparam equal_791_i15_4_lut_LC_16_19_7.SEQ_MODE=4'b0000;
    defparam equal_791_i15_4_lut_LC_16_19_7.LUT_INIT=16'b1111111011111111;
    LogicCell40 equal_791_i15_4_lut_LC_16_19_7 (
            .in0(N__47778),
            .in1(N__50288),
            .in2(N__50615),
            .in3(N__49002),
            .lcout(n15_adj_750),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_243_LC_16_20_0.C_ON=1'b0;
    defparam i1_4_lut_adj_243_LC_16_20_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_243_LC_16_20_0.LUT_INIT=16'b1100111110001111;
    LogicCell40 i1_4_lut_adj_243_LC_16_20_0 (
            .in0(N__47741),
            .in1(N__48747),
            .in2(N__49772),
            .in3(N__49143),
            .lcout(n30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_242_LC_16_20_1.C_ON=1'b0;
    defparam i2_3_lut_adj_242_LC_16_20_1.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_242_LC_16_20_1.LUT_INIT=16'b0010001000110011;
    LogicCell40 i2_3_lut_adj_242_LC_16_20_1 (
            .in0(N__47718),
            .in1(N__49517),
            .in2(_gnd_net_),
            .in3(N__47685),
            .lcout(n6_adj_766),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam state__i1_LC_16_20_3.C_ON=1'b0;
    defparam state__i1_LC_16_20_3.SEQ_MODE=4'b1000;
    defparam state__i1_LC_16_20_3.LUT_INIT=16'b0111010001000100;
    LogicCell40 state__i1_LC_16_20_3 (
            .in0(N__49749),
            .in1(N__49955),
            .in2(N__47664),
            .in3(N__47643),
            .lcout(state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48442),
            .ce(N__50816),
            .sr(N__50787));
    defparam state__i0_LC_16_20_4.C_ON=1'b0;
    defparam state__i0_LC_16_20_4.SEQ_MODE=4'b1000;
    defparam state__i0_LC_16_20_4.LUT_INIT=16'b0101010100010001;
    LogicCell40 state__i0_LC_16_20_4 (
            .in0(N__49954),
            .in1(N__49750),
            .in2(_gnd_net_),
            .in3(N__47631),
            .lcout(state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48442),
            .ce(N__50816),
            .sr(N__50787));
    defparam i4_4_lut_adj_246_LC_17_15_0.C_ON=1'b0;
    defparam i4_4_lut_adj_246_LC_17_15_0.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_246_LC_17_15_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i4_4_lut_adj_246_LC_17_15_0 (
            .in0(N__47597),
            .in1(N__47582),
            .in2(N__47571),
            .in3(N__47549),
            .lcout(),
            .ltout(n10_adj_762_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_3_lut_adj_247_LC_17_15_1.C_ON=1'b0;
    defparam i5_3_lut_adj_247_LC_17_15_1.SEQ_MODE=4'b0000;
    defparam i5_3_lut_adj_247_LC_17_15_1.LUT_INIT=16'b1111111111111100;
    LogicCell40 i5_3_lut_adj_247_LC_17_15_1 (
            .in0(_gnd_net_),
            .in1(N__48176),
            .in2(N__48165),
            .in3(N__48161),
            .lcout(n18_adj_742),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_895_i11_2_lut_4_lut_LC_17_15_6.C_ON=1'b0;
    defparam equal_895_i11_2_lut_4_lut_LC_17_15_6.SEQ_MODE=4'b0000;
    defparam equal_895_i11_2_lut_4_lut_LC_17_15_6.LUT_INIT=16'b1111111111101111;
    LogicCell40 equal_895_i11_2_lut_4_lut_LC_17_15_6 (
            .in0(N__50499),
            .in1(N__48913),
            .in2(N__50332),
            .in3(N__50753),
            .lcout(n11_adj_739),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_LC_17_16_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_17_16_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_17_16_0.LUT_INIT=16'b0000000010000000;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_17_16_0 (
            .in0(N__50492),
            .in1(N__48845),
            .in2(N__50754),
            .in3(N__48646),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9317_3_lut_LC_17_16_1.C_ON=1'b0;
    defparam i9317_3_lut_LC_17_16_1.SEQ_MODE=4'b0000;
    defparam i9317_3_lut_LC_17_16_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i9317_3_lut_LC_17_16_1 (
            .in0(N__48843),
            .in1(N__48077),
            .in2(_gnd_net_),
            .in3(N__48038),
            .lcout(),
            .ltout(n13164_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_1__bdd_4_lut_LC_17_16_2.C_ON=1'b0;
    defparam current_pin_1__bdd_4_lut_LC_17_16_2.SEQ_MODE=4'b0000;
    defparam current_pin_1__bdd_4_lut_LC_17_16_2.LUT_INIT=16'b1110110001100100;
    LogicCell40 current_pin_1__bdd_4_lut_LC_17_16_2 (
            .in0(N__50491),
            .in1(N__50204),
            .in2(N__48009),
            .in3(N__47820),
            .lcout(n13468),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_280_i6_2_lut_LC_17_16_4.C_ON=1'b0;
    defparam equal_280_i6_2_lut_LC_17_16_4.SEQ_MODE=4'b0000;
    defparam equal_280_i6_2_lut_LC_17_16_4.LUT_INIT=16'b1111111100110011;
    LogicCell40 equal_280_i6_2_lut_LC_17_16_4 (
            .in0(_gnd_net_),
            .in1(N__50205),
            .in2(_gnd_net_),
            .in3(N__48844),
            .lcout(n6_adj_748),
            .ltout(n6_adj_748_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i488_4_lut_LC_17_16_5.C_ON=1'b0;
    defparam i488_4_lut_LC_17_16_5.SEQ_MODE=4'b0000;
    defparam i488_4_lut_LC_17_16_5.LUT_INIT=16'b1010101010101000;
    LogicCell40 i488_4_lut_LC_17_16_5 (
            .in0(N__47928),
            .in1(N__50595),
            .in2(N__47886),
            .in3(N__49146),
            .lcout(n2421),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9318_3_lut_LC_17_16_7.C_ON=1'b0;
    defparam i9318_3_lut_LC_17_16_7.SEQ_MODE=4'b0000;
    defparam i9318_3_lut_LC_17_16_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 i9318_3_lut_LC_17_16_7 (
            .in0(N__48842),
            .in1(N__47883),
            .in2(_gnd_net_),
            .in3(N__47843),
            .lcout(n13165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_i0_i0_LC_17_17_0.C_ON=1'b1;
    defparam current_pin_i0_i0_LC_17_17_0.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i0_LC_17_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i0_LC_17_17_0 (
            .in0(_gnd_net_),
            .in1(N__48894),
            .in2(_gnd_net_),
            .in3(N__47814),
            .lcout(current_pin_0),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(n10384),
            .clk(N__48433),
            .ce(N__48234),
            .sr(N__48222));
    defparam current_pin_i0_i1_LC_17_17_1.C_ON=1'b1;
    defparam current_pin_i0_i1_LC_17_17_1.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i1_LC_17_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i1_LC_17_17_1 (
            .in0(_gnd_net_),
            .in1(N__50316),
            .in2(_gnd_net_),
            .in3(N__48711),
            .lcout(current_pin_1),
            .ltout(),
            .carryin(n10384),
            .carryout(n10385),
            .clk(N__48433),
            .ce(N__48234),
            .sr(N__48222));
    defparam current_pin_i0_i2_LC_17_17_2.C_ON=1'b1;
    defparam current_pin_i0_i2_LC_17_17_2.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i2_LC_17_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i2_LC_17_17_2 (
            .in0(_gnd_net_),
            .in1(N__50490),
            .in2(_gnd_net_),
            .in3(N__48708),
            .lcout(current_pin_2),
            .ltout(),
            .carryin(n10385),
            .carryout(n10386),
            .clk(N__48433),
            .ce(N__48234),
            .sr(N__48222));
    defparam current_pin_i0_i3_LC_17_17_3.C_ON=1'b1;
    defparam current_pin_i0_i3_LC_17_17_3.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i3_LC_17_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i3_LC_17_17_3 (
            .in0(_gnd_net_),
            .in1(N__50712),
            .in2(_gnd_net_),
            .in3(N__48705),
            .lcout(current_pin_3),
            .ltout(),
            .carryin(n10386),
            .carryout(n10387),
            .clk(N__48433),
            .ce(N__48234),
            .sr(N__48222));
    defparam current_pin_i0_i4_LC_17_17_4.C_ON=1'b1;
    defparam current_pin_i0_i4_LC_17_17_4.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i4_LC_17_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i4_LC_17_17_4 (
            .in0(_gnd_net_),
            .in1(N__48647),
            .in2(_gnd_net_),
            .in3(N__48576),
            .lcout(current_pin_4),
            .ltout(),
            .carryin(n10387),
            .carryout(n10388),
            .clk(N__48433),
            .ce(N__48234),
            .sr(N__48222));
    defparam current_pin_i0_i5_LC_17_17_5.C_ON=1'b1;
    defparam current_pin_i0_i5_LC_17_17_5.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i5_LC_17_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i5_LC_17_17_5 (
            .in0(_gnd_net_),
            .in1(N__48559),
            .in2(_gnd_net_),
            .in3(N__48537),
            .lcout(current_pin_5),
            .ltout(),
            .carryin(n10388),
            .carryout(n10389),
            .clk(N__48433),
            .ce(N__48234),
            .sr(N__48222));
    defparam current_pin_i0_i6_LC_17_17_6.C_ON=1'b1;
    defparam current_pin_i0_i6_LC_17_17_6.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i6_LC_17_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i6_LC_17_17_6 (
            .in0(_gnd_net_),
            .in1(N__48526),
            .in2(_gnd_net_),
            .in3(N__48498),
            .lcout(current_pin_6),
            .ltout(),
            .carryin(n10389),
            .carryout(n10390),
            .clk(N__48433),
            .ce(N__48234),
            .sr(N__48222));
    defparam current_pin_i0_i7_LC_17_17_7.C_ON=1'b0;
    defparam current_pin_i0_i7_LC_17_17_7.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i7_LC_17_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i7_LC_17_17_7 (
            .in0(_gnd_net_),
            .in1(N__48481),
            .in2(_gnd_net_),
            .in3(N__48495),
            .lcout(current_pin_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48433),
            .ce(N__48234),
            .sr(N__48222));
    defparam i4172_2_lut_LC_17_18_1.C_ON=1'b0;
    defparam i4172_2_lut_LC_17_18_1.SEQ_MODE=4'b0000;
    defparam i4172_2_lut_LC_17_18_1.LUT_INIT=16'b0101010100000000;
    LogicCell40 i4172_2_lut_LC_17_18_1 (
            .in0(N__49752),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50815),
            .lcout(n7409),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_LC_17_18_2.C_ON=1'b0;
    defparam i13_4_lut_LC_17_18_2.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_17_18_2.LUT_INIT=16'b1111111111001000;
    LogicCell40 i13_4_lut_LC_17_18_2 (
            .in0(N__49145),
            .in1(N__49290),
            .in2(N__48201),
            .in3(N__49368),
            .lcout(n42),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_LC_17_18_3.C_ON=1'b0;
    defparam i11_4_lut_LC_17_18_3.SEQ_MODE=4'b0000;
    defparam i11_4_lut_LC_17_18_3.LUT_INIT=16'b1110111011101100;
    LogicCell40 i11_4_lut_LC_17_18_3 (
            .in0(N__49263),
            .in1(N__49359),
            .in2(N__49350),
            .in3(N__49144),
            .lcout(),
            .ltout(n40_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i25_4_lut_LC_17_18_4.C_ON=1'b0;
    defparam i25_4_lut_LC_17_18_4.SEQ_MODE=4'b0000;
    defparam i25_4_lut_LC_17_18_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i25_4_lut_LC_17_18_4 (
            .in0(N__49323),
            .in1(N__49311),
            .in2(N__49305),
            .in3(N__49302),
            .lcout(n54_adj_768),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_0__bdd_4_lut_9619_LC_17_19_0.C_ON=1'b0;
    defparam current_pin_0__bdd_4_lut_9619_LC_17_19_0.SEQ_MODE=4'b0000;
    defparam current_pin_0__bdd_4_lut_9619_LC_17_19_0.LUT_INIT=16'b1011101111000000;
    LogicCell40 current_pin_0__bdd_4_lut_9619_LC_17_19_0 (
            .in0(N__49283),
            .in1(N__50284),
            .in2(N__49259),
            .in3(N__48968),
            .lcout(),
            .ltout(n13444_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13444_bdd_4_lut_LC_17_19_1.C_ON=1'b0;
    defparam n13444_bdd_4_lut_LC_17_19_1.SEQ_MODE=4'b0000;
    defparam n13444_bdd_4_lut_LC_17_19_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n13444_bdd_4_lut_LC_17_19_1 (
            .in0(N__50285),
            .in1(N__49226),
            .in2(N__49194),
            .in3(N__49187),
            .lcout(n13447),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_919_i15_4_lut_LC_17_19_4.C_ON=1'b0;
    defparam equal_919_i15_4_lut_LC_17_19_4.SEQ_MODE=4'b0000;
    defparam equal_919_i15_4_lut_LC_17_19_4.LUT_INIT=16'b1111111011111111;
    LogicCell40 equal_919_i15_4_lut_LC_17_19_4 (
            .in0(N__49142),
            .in1(N__50286),
            .in2(N__50607),
            .in3(N__48969),
            .lcout(),
            .ltout(n15_adj_749_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_adj_240_LC_17_19_5.C_ON=1'b0;
    defparam i8_4_lut_adj_240_LC_17_19_5.SEQ_MODE=4'b0000;
    defparam i8_4_lut_adj_240_LC_17_19_5.LUT_INIT=16'b1110110010100000;
    LogicCell40 i8_4_lut_adj_240_LC_17_19_5 (
            .in0(N__48774),
            .in1(N__49095),
            .in2(N__49065),
            .in3(N__49062),
            .lcout(n37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Mux_34_i19_3_lut_LC_17_19_7.C_ON=1'b0;
    defparam Mux_34_i19_3_lut_LC_17_19_7.SEQ_MODE=4'b0000;
    defparam Mux_34_i19_3_lut_LC_17_19_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 Mux_34_i19_3_lut_LC_17_19_7 (
            .in0(N__48967),
            .in1(N__48773),
            .in2(_gnd_net_),
            .in3(N__48746),
            .lcout(n19_adj_715),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9261_4_lut_4_lut_LC_17_20_5.C_ON=1'b0;
    defparam i9261_4_lut_4_lut_LC_17_20_5.SEQ_MODE=4'b0000;
    defparam i9261_4_lut_4_lut_LC_17_20_5.LUT_INIT=16'b1110100010101000;
    LogicCell40 i9261_4_lut_4_lut_LC_17_20_5 (
            .in0(N__49524),
            .in1(N__49941),
            .in2(N__49796),
            .in3(N__50859),
            .lcout(),
            .ltout(n13037_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_244_LC_17_20_6.C_ON=1'b0;
    defparam i2_4_lut_adj_244_LC_17_20_6.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_244_LC_17_20_6.LUT_INIT=16'b0000111100001110;
    LogicCell40 i2_4_lut_adj_244_LC_17_20_6 (
            .in0(N__50853),
            .in1(N__50844),
            .in2(N__50832),
            .in3(N__50829),
            .lcout(n7249),
            .ltout(n7249_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4158_2_lut_4_lut_LC_17_20_7.C_ON=1'b0;
    defparam i4158_2_lut_4_lut_LC_17_20_7.SEQ_MODE=4'b0000;
    defparam i4158_2_lut_4_lut_LC_17_20_7.LUT_INIT=16'b0000000000100000;
    LogicCell40 i4158_2_lut_4_lut_LC_17_20_7 (
            .in0(N__49525),
            .in1(N__49942),
            .in2(N__50790),
            .in3(N__49697),
            .lcout(n7395),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_927_i10_2_lut_LC_18_16_2.C_ON=1'b0;
    defparam equal_927_i10_2_lut_LC_18_16_2.SEQ_MODE=4'b0000;
    defparam equal_927_i10_2_lut_LC_18_16_2.LUT_INIT=16'b1100110011111111;
    LogicCell40 equal_927_i10_2_lut_LC_18_16_2 (
            .in0(_gnd_net_),
            .in1(N__50687),
            .in2(_gnd_net_),
            .in3(N__50444),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6234_2_lut_LC_18_16_5.C_ON=1'b0;
    defparam i6234_2_lut_LC_18_16_5.SEQ_MODE=4'b0000;
    defparam i6234_2_lut_LC_18_16_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 i6234_2_lut_LC_18_16_5 (
            .in0(N__50445),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50256),
            .lcout(n9456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_218_LC_18_18_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_218_LC_18_18_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_218_LC_18_18_5.LUT_INIT=16'b1111111110111011;
    LogicCell40 i1_2_lut_3_lut_adj_218_LC_18_18_5 (
            .in0(N__50014),
            .in1(N__49773),
            .in2(_gnd_net_),
            .in3(N__49509),
            .lcout(n15_adj_721),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
