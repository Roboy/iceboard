// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Thu Feb  6 13:05:38 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, INLC_c_0, INHC_c_0, 
        INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, n36530, GHB, 
        GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire h1, h2, h3, n15, n14;
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(116[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(117[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(126[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(223[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(225[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(226[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(227[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(228[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(229[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(231[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(232[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(233[22:35])
    
    wire n41281, n41280, n36240;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(263[22:33])
    
    wire n41694;
    wire [7:0]data;   // verilog/TinyFPGA_B.v(326[14:18])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(350[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(358[15:20])
    
    wire pwm_setpoint_23__N_215;
    wire [23:0]pwm_setpoint_23__N_191;
    
    wire n46663, n40892, n33, n32, n31, n30, n29, n28, n27, 
        n26, n25, n24, n23, n22, n21, n20, n19, n18, n4;
    wire [7:0]commutation_state_7__N_216;
    
    wire commutation_state_7__N_224;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(222[11:28])
    
    wire n861, n10, GHA_N_367, GLA_N_384, GHB_N_389, GLB_N_398, 
        GHC_N_403, GLC_N_412, dti_N_416, RX_N_10, n1617;
    wire [31:0]motor_state_23__N_123;
    wire [32:0]encoder0_position_scaled_23__N_51;
    
    wire encoder1_position_scaled_23__N_279;
    wire [31:0]encoder1_position_scaled_23__N_75;
    wire [23:0]displacement_23__N_99;
    
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
        n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
        n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
        n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
        n50106, n1195, n4_adj_5096, n516, n41279, n1658;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(224[11:28])
    
    wire n41278;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n41277, n40891, n4_adj_5097, n41693, n17, n16, n15_adj_5098, 
        n14_adj_5099, n834, n833, n832, n831, n830, n829, n828, 
        n40890;
    wire [3:0]state_3__N_528;
    
    wire n40889, n40888, n41276, n27954, n50220, n41081, n6935, 
        n41080, n41079, n29671, n41275, n40456, n13, n41274, n41931, 
        n41078, n41077, n6662, n41076, n41273, n41930, n10_adj_5100, 
        n731, n41929, n29670, n29669, n3684, n41928, n36608, n4_adj_5101, 
        n41927, n8, n41926, n41925, n41692, n29668, n29667, n29666, 
        n29665, n41691, n40404, n41690, n29664, n29663, n29662, 
        n45289, n41272, n41689, n41075, n41271, n29661, n29660, 
        n29659, n29658, n29657, n41924, n41688, n29656, n29655, 
        n41687, n41686, n41270, n41269, n41685, n41268, n29654, 
        n29653, n41923, n41074, n41922, n41684, n41267, n53039, 
        n41683, n41073, n29652, n41921;
    wire [2:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n29651, n41920, n29650, n41682, n29649, n41072, n41071, 
        n41681, n41919, n41266, n41680, n3, n4_adj_5102, n5, n6, 
        n7, n8_adj_5103, n9, n10_adj_5104, n11, n12, n13_adj_5105, 
        n14_adj_5106, n15_adj_5107, n16_adj_5108, n17_adj_5109, n18_adj_5110, 
        n19_adj_5111, n20_adj_5112, n21_adj_5113, n22_adj_5114, n23_adj_5115, 
        n24_adj_5116, n25_adj_5117, n41070, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n40455, n41265, n36384, n41679, n41069, n40454;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n41264, n41068, n41067, n41263, n41918, n41678, n122, 
        n123, n41677, n41676, n41675, n41674, n41917, n41916, 
        n41673, n41262, n41261, n41066, n41915, n41672, n41260, 
        n29648, n46756, n29647, n41671, n41670, n41065, n41669, 
        n41914, n771, n41913, n41259, n41258, n41064, n41912, 
        n41063, n41062, n41061, n41060, n40453, n41257, n41911, 
        n41256, n40403, n41059, n41668, n51552, n41058, n41910, 
        n41667, n41057, n41255, n21721, n41909, n41254, n41253, 
        n41056, n41908, n41252, n41251, n41055, n40452, n41666, 
        n41665, n41054, n41250, n41249, n41053, n41664, n41907, 
        n41248, n40451, n47281, n41052, n41247, n41663, n41051, 
        n41906, n41662, n41246, n41245, n41905, n41050, n46745, 
        n41244, n41049, n41904, n41903, n41902, n41048, n41901, 
        n41243, n40450, n40695, n40694, n40388, n40449, n41661, 
        n40402, n40448, n46666, n41047, n41660, n40693, n46671, 
        n41659, n35272, n41658, n40692, n41242, n40691, n41241, 
        n41240, n41046, n41239, n41045, n41657, n41656, n41655, 
        n40447, n41238, n41044, n40690, n41043, n36536, n41654, 
        n41653, n41042, n40689, n36532, n40688, n40687, n41652, 
        n41651, n40686, n40446, n36510, n41650, n40401, n40445, 
        n41237, n41649, n40444, n40443, n40685, n41648, n40442, 
        n36244, n41236, n41647, n41235, n41234, n41041, n41233, 
        n41428, n41040, n41039, n41038, n41646, n41427, n41426, 
        n41645, n40684, n41232, n41037, n41644, n41231, n41425, 
        n41424, n41230, n40683, n41643, n41036, n41035, n40682, 
        n41642, n41034, n40400, n36490, n40441, n36488, n41423, 
        n40681, n41229, n41422, n41033, n40440, n40680, n40439, 
        n40438, n41641, n40437, n41032, n41228, n40387, n36484, 
        n41640, n41227, n36520, n41639, n41638, n41637, n40436, 
        n41636, n41421, n41226, n40679, n41420, n41225, n41419, 
        n40678, n40677, n41635, n41634, n41418, n36522, n40676, 
        n41224, n40675, n41417, n41416, n40674, n41223, n41222, 
        n41221, n41633, n41220, n41415, n41414, n41413, n41632, 
        n41412, n41219, n40552, n41411, n41410, n41218, n41217, 
        n40673, n41409, n41631, n41630, n41408, n41216, n41629, 
        n41628, n41407, n41627, n35426, n41215, n40551, n40550, 
        n41626, n41406, n41214, n41213, n46395, n113, n41212, 
        n41405, n52505, n114, n41625, n40435, n41624, n41404, 
        n41211, n41210, n41403, n41623, n2, n29646, n29645, n29644, 
        n29643, n7287, n7286, n7285, n7283, n7282, n41209, n41622, 
        n41621, n41620, n41619, n3303, n14_adj_5118;
    wire [31:0]\FRAME_MATCHER.state_31__N_2788 ;
    
    wire n41618, n10_adj_5119, n41617, n41208, n41616, n53005, n41615, 
        n41614, n41207, n41613, n40549, n41206, n41612, n41205, 
        n41611, n41610, n40434, n41609, n41608, n40433, n41204, 
        n41607, n40399, n41203, n41202, n40386, n41606, n41201, 
        n41200, n41605, n41604, n41603, n41602, n41199, n40548, 
        n41198, n41601, n41600, n41599, n41598, n4_adj_5120, n41197, 
        n29642, n29639, n4452, n40432, n40431, n40430, n41196, 
        n52089, n41195, n41194, n41193, n41192, n41191, n41190, 
        n41189, n41188, n41187, n4_adj_5121, n10_adj_5122, n52972, 
        n5_adj_5123, n29638, n29637, n40429, n29636, n29635, n29634, 
        n29633, \FRAME_MATCHER.i_31__N_2626 , n46749, n36189, n46425, 
        n27761, n46765, n45528, n44751, n36412, n41176, n652, 
        n29632, n625, n623, n622, n621, n41175, n36430, n53345, 
        n46713, n46728, n15_adj_5124, n25_adj_5125, n24_adj_5126, 
        n23_adj_5127, n22_adj_5128, n21_adj_5129, n20_adj_5130, n19_adj_5131, 
        n18_adj_5132, n17_adj_5133, n16_adj_5134, n29631, n29630, 
        n29629, n29628, n29627, n29626, n29625, n29624, n29623, 
        n29622, n29621, n29620, n29619, n29618, n29617, n29616, 
        n15_adj_5135, n14_adj_5136, n13_adj_5137, n12_adj_5138, n11_adj_5139, 
        n10_adj_5140, n9_adj_5141, n41174, n41173, n40428, n14_adj_5142, 
        n41172, n8_adj_5143, n7_adj_5144, n6_adj_5145, n5_adj_5146, 
        n4_adj_5147, n3_adj_5148, n5741, n40427, n10_adj_5149, n30125, 
        n30122, n30121, n46786, n30120, n30119, n41171, n30118, 
        n30117, n29615, n30116, n25316, n30115, n30114, n29614, 
        n30113, n30112, n30111, n30110, n30109, n30108, n30107, 
        n30106, n30105, n41170, n15_adj_5150, n30104, n30103, n30102, 
        n53344, n30101, n30100, n30099, n30098, n30097, n30096, 
        n30095, n30094, n30093, n30092;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev, n30091, n36402, n30090, n30089, n30088, n30087, 
        n30086, n12_adj_5151, n30085, n30084, n30083, n30082, n30081, 
        n30080, n30079, n30078, direction_N_3907, n30077, n30076, 
        n30075, n30074, n30073, n30072, n30071, n30070, n30069, 
        n30068, n63, n30067, n30066, n30065, n30064, n30063, n30062, 
        n30061, n30060, n30059, n30058, n30057, n30056, n30055, 
        n30054, n30053, n30052, n41169, n30051, n30050, n30049, 
        n41168, n41167, n50212, n30048, n30047;
    wire [1:0]a_new_adj_5272;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev_adj_5153, n30046, n1910, n30045, n30044, n35513, 
        n11_adj_5154, n10_adj_5155, n30043, n30042, n30041, n30040, 
        n30039, n30038, n30037, n30036, n4_adj_5156, direction_N_3907_adj_5157, 
        n30035, n30034, n30033, n30032, n30031, n30030, n30029, 
        n30028, n30027, n30026, n30025, n30024, n30023, n30022, 
        n30021, n30020, n30019, n30018, n30017, n30016, n30015, 
        n30014, n30013, n30012, n41166, n30011, n30010, n30009, 
        n30008, n30007, n30006, n30005, n30004, n30003, n30002, 
        n30001, n30000, n29999, n29998, n9_adj_5158, rw;
    wire [7:0]state_adj_5296;   // verilog/eeprom.v(23[11:16])
    
    wire n8_adj_5161, n7_adj_5162, n6_adj_5163, n5_adj_5164, n4_adj_5165, 
        n3_adj_5166, n2_adj_5167, n29997, n29996, n29995, n29994, 
        n29993, n29991, n29990, n29989, n29988, n29987, n29986, 
        n29985, n29984, n29983, n29982, n52940, n29981, n29980, 
        n29979, n29978, n29977, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n29976, n29975, n29974, n29973, n29972, n29971, n29970, 
        n29969, n41165, n35507, n41164, n29968, n29967, n46392, 
        n29966, n29965;
    wire [2:0]r_SM_Main_2__N_3542;
    
    wire n29964, n29963, n29962, n29613, n29961, n29960, n29959, 
        n29958, n29957, n29956, n29955, n29954, n29953, n29952, 
        n29951, n29950, n29949;
    wire [2:0]r_SM_Main_adj_5305;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5307;   // verilog/uart_tx.v(33[16:27])
    
    wire n40426, n40398;
    wire [2:0]r_SM_Main_2__N_3613;
    
    wire n29948, n40385, n48426, n46691, n29947, n36376, n29946, 
        n29945, n29944, n29943, n29942, n29941, n29940, n29939, 
        n29938, n29937, n29936, n29935, n29934, n29933, n29932, 
        n29931, n29930, n29929, n29928, n29927, n29926, n29925, 
        n29612;
    wire [7:0]state_adj_5316;   // verilog/i2c_controller.v(33[12:17])
    
    wire n29924, n29923;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n29922, n29921, n29920, n29919, enable_slow_N_4190, n40457, 
        n29918, n29917, n29916, n29915;
    wire [7:0]state_7__N_4087;
    
    wire n29914, n29913, n29611, n6387, n29912, n29911, n29910, 
        n29909, n29908, n29907, n29906, n29905, n29904;
    wire [7:0]state_7__N_4103;
    
    wire n29903, n29902, n29901, n29900, n29899, n29898, n29897, 
        n41163, n41162, n41161, n36372, n46818, n29896, n29895, 
        n36378, n46682, n29894, n29893, n29892, n29610, n29609, 
        n29608, n29607, n29606, n29891, n45591, n6970, n29890, 
        n29889, n29888, n29887, n29886, n29885, n29884, n29883, 
        n29882, n29881, n29880, n29879, n29878, n29877, n29876, 
        n29875, n29874, n29252, n29873, n29872, n29871, n29870, 
        n29869, n29868, n29867, n29866, n29865, n29864, n29863, 
        n29862, n29861, n29860, n29859, n29858, n29857, n29856, 
        n29855, n41160, n41159, n29854, n29853, n896, n897, n898, 
        n899, n900, n901, n29852, n927, n928, n929, n930, n931, 
        n932, n933, n934, n935, n936, n937, n938, n939, n940, 
        n941, n942, n943, n944, n945, n946, n947, n948, n949, 
        n950, n951, n952, n953, n954, n955, n956, n957, n960, 
        n995, n996, n997, n998, n999, n1000, n1001, n1026, n1027, 
        n1028, n1029, n1030, n1031, n1032, n1033, n1059, n1093_adj_5173, 
        n1094_adj_5174, n1095_adj_5175, n1096_adj_5176, n1097_adj_5177, 
        n1098_adj_5178, n1099_adj_5179, n1100_adj_5180, n1101_adj_5181, 
        n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
        n1133, n1158, n20247, n1193, n1194, n1195_adj_5182, n1196, 
        n1197, n1198, n1199, n1200, n1201, n1224, n1225, n1226, 
        n1227, n1228, n1229, n1230, n1231, n1232, n1233, n52524, 
        n1257, n1292, n1293, n1294, n1295, n1296, n1297, n1298, 
        n1299, n1300, n1301, n1323, n1324, n1325, n1326, n1327, 
        n1328, n1329, n1330, n1331, n1332, n1333, n1356, n1391, 
        n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
        n1400, n1401, n1422, n1423, n1424, n1425, n1426, n1427, 
        n1428, n1429, n1430, n1431, n1432, n1433, n1455, n1490, 
        n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
        n1499, n1500, n1501, n1521, n1522, n1523, n1524, n1525, 
        n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
        n1554, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
        n1596, n1597, n1598, n1599, n1600, n1601, n1620, n1621, 
        n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
        n1630, n1631, n1632, n1633, n1653_adj_5183, n27762, n1688, 
        n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
        n1697, n1698, n1699, n1700, n1701, n1719, n1720, n1721, 
        n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
        n1730, n1731, n1732, n1733, n1752, n1787, n1788, n1789, 
        n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, 
        n1798, n1799, n1800, n1801, n1818, n1819, n1820, n1821, 
        n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
        n1830, n1831, n1832, n1833, n36398, n1851, n1886, n1887, 
        n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, 
        n1896, n1897, n1898, n1899, n1900, n1901, n29851, n29186, 
        n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, 
        n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
        n1933, n1950, n29175, n1985, n1986, n1987, n1988, n1989, 
        n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
        n1998, n1999, n2000, n2001, n2016, n2017, n2018, n2019, 
        n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
        n2028, n2029, n2030, n2031, n2032, n2033, n2049, n2084, 
        n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
        n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, 
        n2101, n29165, n2115, n2116, n2117, n2118, n2119, n2120, 
        n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, 
        n2129, n2130, n2131, n2132, n2133, n29850, n2148, n29849, 
        n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, 
        n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, 
        n2199, n2200, n2201, n45179, n2214, n2215, n2216, n2217, 
        n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, 
        n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, 
        n2247, n29848, n29137, n2282, n2283, n2284, n2285, n2286, 
        n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
        n2295, n2296, n2297, n2298, n2299, n2300, n2301, n40425, 
        n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
        n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, 
        n2329, n2330, n2331, n2332, n2333, n2346, n8_adj_5184, 
        n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
        n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
        n2397, n2398, n2399, n2400, n2401, n40397, n2412, n2413, 
        n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, 
        n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, 
        n2430, n2431, n2432, n2433, n2445, n2480, n2481, n2482, 
        n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
        n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
        n2499, n2500, n2501, n2511, n2512, n2513, n2514, n2515, 
        n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, 
        n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, 
        n2532, n2533, n2544, n29106, n29394, n2579, n2580, n2581, 
        n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, 
        n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, 
        n2598, n2599, n2600, n2601, n2610, n2611, n2612, n2613, 
        n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, 
        n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
        n2630, n2631, n2632, n2633, n44527, n2643, n45588, n2678, 
        n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
        n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, 
        n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2709, 
        n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
        n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, 
        n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
        n2742, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
        n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, 
        n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
        n2800, n2801, n2808, n2809, n2810, n2811, n2812, n2813, 
        n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, 
        n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
        n2830, n2831, n2832, n2833, n2841, n29375, n2876, n2877, 
        n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
        n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
        n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
        n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, 
        n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, 
        n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, 
        n2931, n2932, n2933, n2940, n2975, n2976, n2977, n2978, 
        n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
        n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, 
        n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3006, 
        n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, 
        n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
        n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, 
        n3031, n3032, n3033, n3039, n29048, n3074, n3075, n3076, 
        n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, 
        n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
        n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, 
        n3101, n3105, n3106, n3107, n3108, n3109, n3110, n3111, 
        n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, 
        n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, 
        n3128, n3129, n3130, n3131, n3132, n3133, n53043, n3138, 
        n29044, n3173, n3174, n3175, n3176, n3177, n3178, n3179, 
        n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, 
        n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, 
        n3196, n3197, n3198, n3199, n3200, n3201, n3204, n3205, 
        n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, 
        n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, 
        n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, 
        n3230, n3231, n3232, n3233, n53077, n3237, n3272, n3273, 
        n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
        n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
        n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3298, 
        n3299, n3300, n3301, n24_adj_5185, n47661, n62, n27787, 
        n27790, n49269, n41158, n52615, n5_adj_5186, n49261, n49255, 
        n52908, n7_adj_5187, n63_adj_5188, n49249, n29600, n49243, 
        n27911, n29598, n29597, n29596, n49237, n29595, n29594, 
        n49235, n49231, n41157, n52491, n27946, n27898, n49225, 
        n7284, n6_adj_5189, n12_adj_5190, n41156, n53403, n48, n49, 
        n50, n51, n52, n53, n54, n55, n41155, n41154, n51822, 
        n52590, n41550, n41549, n49213, n41548, n41547, n7_adj_5191, 
        n8_adj_5192, n51830, n4_adj_5193, n49207, n49201, n49195, 
        n49189, n49187, n49185, n29591, n29587, n29583, n29582, 
        n29579, n29578, n29575, n29570, n29569, n29567, n29566, 
        n29565, n29564, n29563, n29561, n49163, n41153, n41152, 
        n41151, n40788, n40787, n49157, n49151, n29560, n29559, 
        n29558, n29557, n29556, n29555, n41546, n29544, n49145, 
        n49143, n52874, n49135, n2_adj_5194, n3_adj_5195, n4_adj_5196, 
        n5_adj_5197, n6_adj_5198, n7_adj_5199, n8_adj_5200, n9_adj_5201, 
        n10_adj_5202, n11_adj_5203, n12_adj_5204, n13_adj_5205, n14_adj_5206, 
        n15_adj_5207, n16_adj_5208, n17_adj_5209, n18_adj_5210, n19_adj_5211, 
        n20_adj_5212, n21_adj_5213, n22_adj_5214, n23_adj_5215, n24_adj_5216, 
        n25_adj_5217, n26_adj_5218, n27_adj_5219, n28_adj_5220, n29_adj_5221, 
        n30_adj_5222, n31_adj_5223, n32_adj_5224, n33_adj_5225, n49127, 
        n48551, n40786, n40785, n49121, n40784, n41545, n41150, 
        n49115, n49113, n40424, n41544, n41149, n41543, n49107, 
        n36382, n49105, n40783, n40782, n49103, n41148, n40781, 
        n40780, n41147, n41146, n49089, n41542, n41541, n41145, 
        n41540, n41539, n40423, n40422, n41538, n40421, n41537, 
        n41536, n41144, n49083, n41143, n41142, n41141, n41140, 
        n41535, n41139, n41138, n41534, n41533, n41532, n51973, 
        n41137, n41136, n41135, n41531, n41530, n41529, n41528, 
        n41527, n40769, n41134, n40768, n40767, n41133, n52571, 
        n40766, n40765, n41526, n41525, n36322, n40764, n40763, 
        n40762, n41132, n49071, n40761, n41131, n41524, n41130, 
        n40760, n40759, n41129, n41128, n41127, n40758, n41126, 
        n41125, n41124, n40757, n41123, n40756, n41122, n40755, 
        n40754, n41121, n40753, n48537, n40752, n49065, n40751, 
        n41120, n46814, n40396, n13_adj_5226, n40750, n40749, n21_adj_5227, 
        n23_adj_5228, n25_adj_5229, n27_adj_5230, n29_adj_5231, n31_adj_5232, 
        n41119, n41, n36300, n41321, n59, n61, n49061, n49055, 
        n49053, n51971, n49043, n10_adj_5233, n52553, n49037, n52846, 
        n5_adj_5234, n7_adj_5235, n4_adj_5236, n49031, n41320, n50269, 
        n50265, n40420, n41319, n49025, n49021, n41318, n48513, 
        n49005, n48999, n48993, n48989, n48985, n41118, n45417, 
        n46774, n41317, n46452, n48975, n50243, n46434, n41316, 
        n46432, n48969, n48965, n51345, n48955, n52807, n48949, 
        n46413, n27765, n50239, n48489, n48943, n50236, n41315, 
        n41314, n44955, n41117, n25059, n46401, n41116, n46394, 
        n48931, n41313, n48925, n41312, n48915, n48911, n41311, 
        n41310, n40419, n41309, n50228, n48901, n47488, n48891, 
        n52784, n48889, n48883, n50223, n52752, n48879, n36316, 
        n41308, n41307, n41306, n41115, n40384, n51326, n48871, 
        n51325, n40395, n41114, n40418, n48865, n41113, n40417, 
        n51324, n47921, n29542, n29541, n48861, n51323, n40416, 
        n29540, n48855, n48853, n29539, n41305, n51322, n51321, 
        n48841, n41112, n51320, n48835, n48829, n48827, n41111, 
        n29538, n41304, n51311, n48821, n52719, n48817, n48815, 
        n41110, n41724, n41303, n41723, n40415, n41722, n41109, 
        n41302, n41108, n40414, n41721, n48803, n41720, n41107, 
        n40383, n40394, n41106, n48797, n41719, n48795, n41301, 
        n48789, n40413, n41718, n40412, n48787, n41300, n41105, 
        n41299, n41298, n48777, n41297, n48771, n41104, n40393, 
        n40411, n40392, n41103, n40391, n41708, n27903, n27784, 
        n48765, n36442, n41296, n41295, n41102, n36256, n41707, 
        n41294, n41101, n52520, n48755, n48751, n40390, n41706, 
        n41705, n40410, n48745, n41704, n40409, n41100, n48737, 
        n40408, n36250, n48731, n48725, n40407, n41703, n41293, 
        n40406, n40382, n41099, n41292, n41098, n40389, n48719, 
        n25095, n48713, n48711, n40381, n48707, n52689, n41702, 
        n41291, n41701, n48699, n48691, n41097, n41096, n41290, 
        n41700, n41095, n41094, n48685, n48679, n48677, n48070, 
        n40897, n48673, n36246, n41699, n41698, n48661, n41697, 
        n41696, n41289, n48651, n48649, n48647, n48645, n40405, 
        n48643, n48641, n41288, n48639, n48637, n45526, n48635, 
        n48631, n48629, n41093, n48627, n40896, n41092, n41695, 
        n48623, n41287, n41286, n48621, n52665, n51281, n48617, 
        n48615, n40895, n40894, n41285, n48611, n48607, n48601, 
        n41284, n40893, n41283, n48595, n48589, n8_adj_5237, n45520, 
        n48583, n48581, n7_adj_5238, n41282, n52641;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i16107_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n44527), .I3(GND_net), .O(n29629));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16108_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n44527), .I3(GND_net), .O(n29630));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16109_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n44527), .I3(GND_net), .O(n29631));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16326_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n48489), .I3(GND_net), 
            .O(n29848));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16327_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n48489), .I3(GND_net), 
            .O(n29849));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16110_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n44527), .I3(GND_net), .O(n29632));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16110_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE dti_177 (.Q(dti), .C(CLK_c), .E(n29044), .D(dti_N_416));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i16111_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n44527), .I3(GND_net), .O(n29633));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16112_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n44527), .I3(GND_net), .O(n29634));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16113_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n44527), .I3(GND_net), .O(n29635));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16114_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n44527), .I3(GND_net), .O(n29636));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16115_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n44527), .I3(GND_net), .O(n29637));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16116_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n44527), .I3(GND_net), .O(n29638));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n40896), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(CLK_c), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(CLK_c), .D(displacement_23__N_99[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i16328_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n48489), .I3(GND_net), 
            .O(n29850));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16328_3_lut.LUT_INIT = 16'hacac;
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4103[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i16117_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n44527), .I3(GND_net), .O(n29639));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16117_3_lut.LUT_INIT = 16'hacac;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i16329_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n48489), .I3(GND_net), 
            .O(n29851));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16330_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n48489), .I3(GND_net), 
            .O(n29852));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16331_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n48489), .I3(GND_net), 
            .O(n29853));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n41121), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n48489));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i16332_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n48489), .I3(GND_net), 
            .O(n29854));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16332_3_lut.LUT_INIT = 16'hacac;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.\state[0] (state[0]), .\state[1] (state[1]), 
            .n44527(n44527), .GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .timer({timer}), .n29252(n29252), .neopxl_color({neopxl_color}), 
            .n29639(n29639), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n29638(n29638), .n29637(n29637), .n29636(n29636), .n29635(n29635), 
            .n29634(n29634), .n29633(n29633), .n29632(n29632), .n29631(n29631), 
            .n29630(n29630), .n29629(n29629), .n29628(n29628), .n29627(n29627), 
            .n29626(n29626), .n29625(n29625), .n29624(n29624), .n29623(n29623), 
            .n29622(n29622), .n29621(n29621), .n29620(n29620), .n29619(n29619), 
            .n29618(n29618), .n29617(n29617), .n29616(n29616), .n29615(n29615), 
            .n29614(n29614), .n29613(n29613), .n29612(n29612), .n29611(n29611), 
            .n29610(n29610), .n29609(n29609), .\state_3__N_528[1] (state_3__N_528[1]), 
            .LED_c(LED_c), .n29544(n29544), .n29539(n29539), .NEOPXL_c(NEOPXL_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[24] 49[2])
    SB_LUT4 i16333_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n29106), .I3(GND_net), .O(n29855));   // verilog/coms.v(127[12] 300[6])
    defparam i16333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16334_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n29106), .I3(GND_net), .O(n29856));   // verilog/coms.v(127[12] 300[6])
    defparam i16334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16335_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n29106), .I3(GND_net), .O(n29857));   // verilog/coms.v(127[12] 300[6])
    defparam i16335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(n771), .I1(n63_adj_5188), .I2(n114), .I3(n45588), 
            .O(n5_adj_5234));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut.LUT_INIT = 16'hcc04;
    SB_LUT4 i3_4_lut (.I0(n7_adj_5191), .I1(\FRAME_MATCHER.state_31__N_2788 [2]), 
            .I2(n8_adj_5192), .I3(n113), .O(n8));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'hfafe;
    SB_LUT4 i4_4_lut (.I0(n122), .I1(n8), .I2(n63), .I3(n5_adj_5234), 
            .O(n53345));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut.LUT_INIT = 16'hefcf;
    SB_LUT4 i16336_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n29106), .I3(GND_net), .O(n29858));   // verilog/coms.v(127[12] 300[6])
    defparam i16336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16337_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n29106), .I3(GND_net), .O(n29859));   // verilog/coms.v(127[12] 300[6])
    defparam i16337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16338_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n29106), .I3(GND_net), .O(n29860));   // verilog/coms.v(127[12] 300[6])
    defparam i16338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16339_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n29106), .I3(GND_net), .O(n29861));   // verilog/coms.v(127[12] 300[6])
    defparam i16339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16340_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n29106), .I3(GND_net), .O(n29862));   // verilog/coms.v(127[12] 300[6])
    defparam i16340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16341_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n29106), .I3(GND_net), .O(n29863));   // verilog/coms.v(127[12] 300[6])
    defparam i16341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16342_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n29106), .I3(GND_net), .O(n29864));   // verilog/coms.v(127[12] 300[6])
    defparam i16342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16343_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n29106), .I3(GND_net), .O(n29865));   // verilog/coms.v(127[12] 300[6])
    defparam i16343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16344_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n29106), .I3(GND_net), .O(n29866));   // verilog/coms.v(127[12] 300[6])
    defparam i16344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16345_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n29106), .I3(GND_net), .O(n29867));   // verilog/coms.v(127[12] 300[6])
    defparam i16345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16346_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n29106), .I3(GND_net), .O(n29868));   // verilog/coms.v(127[12] 300[6])
    defparam i16346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16347_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n29106), .I3(GND_net), .O(n29869));   // verilog/coms.v(127[12] 300[6])
    defparam i16347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16348_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n29106), .I3(GND_net), .O(n29870));   // verilog/coms.v(127[12] 300[6])
    defparam i16348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16349_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n29106), .I3(GND_net), .O(n29871));   // verilog/coms.v(127[12] 300[6])
    defparam i16349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16350_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n29106), .I3(GND_net), .O(n29872));   // verilog/coms.v(127[12] 300[6])
    defparam i16350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16351_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n29106), .I3(GND_net), .O(n29873));   // verilog/coms.v(127[12] 300[6])
    defparam i16351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16352_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n29106), .I3(GND_net), .O(n29874));   // verilog/coms.v(127[12] 300[6])
    defparam i16352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16353_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n29106), .I3(GND_net), .O(n29875));   // verilog/coms.v(127[12] 300[6])
    defparam i16353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16354_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n29106), .I3(GND_net), .O(n29876));   // verilog/coms.v(127[12] 300[6])
    defparam i16354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16355_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n29106), .I3(GND_net), .O(n29877));   // verilog/coms.v(127[12] 300[6])
    defparam i16355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16356_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n25095), .I3(GND_net), .O(n29878));   // verilog/coms.v(127[12] 300[6])
    defparam i16356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16357_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n25095), .I3(GND_net), .O(n29879));   // verilog/coms.v(127[12] 300[6])
    defparam i16357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16358_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n25095), .I3(GND_net), .O(n29880));   // verilog/coms.v(127[12] 300[6])
    defparam i16358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16359_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n25095), .I3(GND_net), .O(n29881));   // verilog/coms.v(127[12] 300[6])
    defparam i16359_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n6662), 
            .D(n1077), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_833_11 (.CI(n40896), .I0(n1225), 
            .I1(VCC_net), .CO(n40897));
    SB_LUT4 encoder0_position_31__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n40895), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_17 (.CI(n41121), .I0(n1819), 
            .I1(VCC_net), .CO(n41122));
    SB_LUT4 add_224_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n40431), .O(encoder1_position_scaled_23__N_75[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n40391), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_10 (.CI(n40895), .I0(n1226), 
            .I1(VCC_net), .CO(n40896));
    SB_LUT4 i16360_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n25095), .I3(GND_net), .O(n29882));   // verilog/coms.v(127[12] 300[6])
    defparam i16360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16361_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n25095), .I3(GND_net), .O(n29883));   // verilog/coms.v(127[12] 300[6])
    defparam i16361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16362_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n25095), .I3(GND_net), .O(n29884));   // verilog/coms.v(127[12] 300[6])
    defparam i16362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16363_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n25095), .I3(GND_net), .O(n29885));   // verilog/coms.v(127[12] 300[6])
    defparam i16363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n40894), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut (.I0(n45588), .I1(\FRAME_MATCHER.i_31__N_2626 ), .I2(n3684), 
            .I3(n4452), .O(n45520));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut.LUT_INIT = 16'hfafe;
    SB_LUT4 i16364_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n25095), .I3(GND_net), .O(n29886));   // verilog/coms.v(127[12] 300[6])
    defparam i16364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(n123), .I1(n45520), .I2(n63_adj_5188), .I3(GND_net), 
            .O(n7_adj_5235));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut.LUT_INIT = 16'h8c8c;
    SB_LUT4 i1_4_lut_adj_1664 (.I0(n113), .I1(n63_adj_5188), .I2(n3303), 
            .I3(n123), .O(n4_adj_5236));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1664.LUT_INIT = 16'h5551;
    SB_LUT4 i3_4_lut_adj_1665 (.I0(n4_adj_5236), .I1(n48070), .I2(n7_adj_5235), 
            .I3(n63), .O(n53344));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1665.LUT_INIT = 16'hfbff;
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n6662), 
            .D(n1078), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n6662), 
            .D(n1079), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n6662), 
            .D(n1080), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n6662), 
            .D(n1081), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n6662), 
            .D(n1082), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n6662), 
            .D(n1083), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16365_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n25095), .I3(GND_net), .O(n29887));   // verilog/coms.v(127[12] 300[6])
    defparam i16365_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n6662), 
            .D(n1084), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n6662), 
            .D(n1085), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n41120), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n6662), 
            .D(n1086), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n6662), 
            .D(n1087), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n6662), 
            .D(n1088), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16366_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n25095), .I3(GND_net), .O(n29888));   // verilog/coms.v(127[12] 300[6])
    defparam i16366_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n6662), 
            .D(n1089), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16367_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n25095), .I3(GND_net), .O(n29889));   // verilog/coms.v(127[12] 300[6])
    defparam i16367_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n6662), 
            .D(n1090), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n6662), 
            .D(n1091), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n6662), 
            .D(n1092), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n6662), 
            .D(n1093), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n6662), 
            .D(n1094), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n6662), 
            .D(n1095), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_833_9 (.CI(n40894), .I0(n1227), 
            .I1(VCC_net), .CO(n40895));
    SB_LUT4 i16368_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n25095), .I3(GND_net), .O(n29890));   // verilog/coms.v(127[12] 300[6])
    defparam i16368_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n6662), 
            .D(n1096), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n6662), 
            .D(n1097), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n6662), 
            .D(n1098), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i37324_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52807));
    defparam i37324_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n6662), 
            .D(n1099), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n6662), 
            .D(n1100), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16369_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n25095), .I3(GND_net), .O(n29891));   // verilog/coms.v(127[12] 300[6])
    defparam i16369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i31_3_lut (.I0(encoder0_position[30]), 
            .I1(n3_adj_5166), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16370_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n25095), .I3(GND_net), .O(n29892));   // verilog/coms.v(127[12] 300[6])
    defparam i16370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16371_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n25095), .I3(GND_net), .O(n29893));   // verilog/coms.v(127[12] 300[6])
    defparam i16371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16372_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n25095), .I3(GND_net), .O(n29894));   // verilog/coms.v(127[12] 300[6])
    defparam i16372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16373_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n25095), .I3(GND_net), .O(n29895));   // verilog/coms.v(127[12] 300[6])
    defparam i16373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[2]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16374_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n25095), .I3(GND_net), .O(n29896));   // verilog/coms.v(127[12] 300[6])
    defparam i16374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16375_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n25095), .I3(GND_net), .O(n29897));   // verilog/coms.v(127[12] 300[6])
    defparam i16375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[3]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16376_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n25095), .I3(GND_net), .O(n29898));   // verilog/coms.v(127[12] 300[6])
    defparam i16376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16377_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n25095), .I3(GND_net), .O(n29899));   // verilog/coms.v(127[12] 300[6])
    defparam i16377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16378_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n25095), .I3(GND_net), .O(n29900));   // verilog/coms.v(127[12] 300[6])
    defparam i16378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16379_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n25095), .I3(GND_net), .O(n29901));   // verilog/coms.v(127[12] 300[6])
    defparam i16379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16380_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n25095), .I3(GND_net), .O(n29902));   // verilog/coms.v(127[12] 300[6])
    defparam i16380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16381_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n25095), .I3(GND_net), .O(n29903));   // verilog/coms.v(127[12] 300[6])
    defparam i16381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16382_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n25095), .I3(GND_net), .O(n29904));   // verilog/coms.v(127[12] 300[6])
    defparam i16382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16383_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n25095), .I3(GND_net), .O(n29905));   // verilog/coms.v(127[12] 300[6])
    defparam i16383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16384_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n25095), .I3(GND_net), .O(n29906));   // verilog/coms.v(127[12] 300[6])
    defparam i16384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16385_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n25095), .I3(GND_net), .O(n29907));   // verilog/coms.v(127[12] 300[6])
    defparam i16385_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1235_16 (.CI(n41120), .I0(n1820), 
            .I1(VCC_net), .CO(n41121));
    SB_LUT4 i16120_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n48426), .I3(GND_net), .O(n29642));   // verilog/coms.v(127[12] 300[6])
    defparam i16120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228), 
            .I2(VCC_net), .I3(n40893), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16386_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n25095), .I3(GND_net), .O(n29908));   // verilog/coms.v(127[12] 300[6])
    defparam i16386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16121_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n48426), .I3(GND_net), .O(n29643));   // verilog/coms.v(127[12] 300[6])
    defparam i16121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16387_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n25095), .I3(GND_net), .O(n29909));   // verilog/coms.v(127[12] 300[6])
    defparam i16387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16122_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n48426), .I3(GND_net), .O(n29644));   // verilog/coms.v(127[12] 300[6])
    defparam i16122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16388_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n25095), .I3(GND_net), .O(n29910));   // verilog/coms.v(127[12] 300[6])
    defparam i16388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16389_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n25095), .I3(GND_net), .O(n29911));   // verilog/coms.v(127[12] 300[6])
    defparam i16389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16390_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n25095), .I3(GND_net), .O(n29912));   // verilog/coms.v(127[12] 300[6])
    defparam i16390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16391_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n25095), .I3(GND_net), .O(n29913));   // verilog/coms.v(127[12] 300[6])
    defparam i16391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16392_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n25095), .I3(GND_net), .O(n29914));   // verilog/coms.v(127[12] 300[6])
    defparam i16392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16123_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n48426), .I3(GND_net), .O(n29645));   // verilog/coms.v(127[12] 300[6])
    defparam i16123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16393_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n25095), .I3(GND_net), .O(n29915));   // verilog/coms.v(127[12] 300[6])
    defparam i16393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16394_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n25095), .I3(GND_net), .O(n29916));   // verilog/coms.v(127[12] 300[6])
    defparam i16394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16395_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n25095), .I3(GND_net), .O(n29917));   // verilog/coms.v(127[12] 300[6])
    defparam i16395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16396_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n25095), .I3(GND_net), .O(n29918));   // verilog/coms.v(127[12] 300[6])
    defparam i16396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16397_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n25095), .I3(GND_net), .O(n29919));   // verilog/coms.v(127[12] 300[6])
    defparam i16397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16398_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n25095), .I3(GND_net), .O(n29920));   // verilog/coms.v(127[12] 300[6])
    defparam i16398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16124_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n48426), .I3(GND_net), .O(n29646));   // verilog/coms.v(127[12] 300[6])
    defparam i16124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16399_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n25095), .I3(GND_net), .O(n29921));   // verilog/coms.v(127[12] 300[6])
    defparam i16399_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n6662), 
            .D(n1101), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16400_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n25095), .I3(GND_net), .O(n29922));   // verilog/coms.v(127[12] 300[6])
    defparam i16400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16125_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n48426), .I3(GND_net), .O(n29647));   // verilog/coms.v(127[12] 300[6])
    defparam i16125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16401_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n25095), .I3(GND_net), .O(n29923));   // verilog/coms.v(127[12] 300[6])
    defparam i16401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16402_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n25095), .I3(GND_net), .O(n29924));   // verilog/coms.v(127[12] 300[6])
    defparam i16402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16403_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n25095), .I3(GND_net), .O(n29925));   // verilog/coms.v(127[12] 300[6])
    defparam i16403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16126_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n48426), .I3(GND_net), .O(n29648));   // verilog/coms.v(127[12] 300[6])
    defparam i16126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16127_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n48426), .I3(GND_net), .O(n29649));   // verilog/coms.v(127[12] 300[6])
    defparam i16127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16128_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n48426), .I3(GND_net), .O(n29650));   // verilog/coms.v(127[12] 300[6])
    defparam i16128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16404_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n25095), 
            .I3(GND_net), .O(n29926));   // verilog/coms.v(127[12] 300[6])
    defparam i16404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16129_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n48426), .I3(GND_net), .O(n29651));   // verilog/coms.v(127[12] 300[6])
    defparam i16129_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n6662), 
            .D(n1108), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n6662), 
            .D(n1107), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n6662), 
            .D(n1106), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n6662), 
            .D(n1105), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n6662), 
            .D(n1104), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n41119), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16130_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n48426), .I3(GND_net), .O(n29652));   // verilog/coms.v(127[12] 300[6])
    defparam i16130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16131_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n48426), .I3(GND_net), .O(n29653));   // verilog/coms.v(127[12] 300[6])
    defparam i16131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[4]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16405_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n25095), 
            .I3(GND_net), .O(n29927));   // verilog/coms.v(127[12] 300[6])
    defparam i16405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16406_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n25095), 
            .I3(GND_net), .O(n29928));   // verilog/coms.v(127[12] 300[6])
    defparam i16406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16407_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n25095), 
            .I3(GND_net), .O(n29929));   // verilog/coms.v(127[12] 300[6])
    defparam i16407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16408_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n25095), 
            .I3(GND_net), .O(n29930));   // verilog/coms.v(127[12] 300[6])
    defparam i16408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16409_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n25095), 
            .I3(GND_net), .O(n29931));   // verilog/coms.v(127[12] 300[6])
    defparam i16409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16410_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n25095), 
            .I3(GND_net), .O(n29932));   // verilog/coms.v(127[12] 300[6])
    defparam i16410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16411_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n25095), 
            .I3(GND_net), .O(n29933));   // verilog/coms.v(127[12] 300[6])
    defparam i16411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16412_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n25095), 
            .I3(GND_net), .O(n29934));   // verilog/coms.v(127[12] 300[6])
    defparam i16412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16413_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n25095), 
            .I3(GND_net), .O(n29935));   // verilog/coms.v(127[12] 300[6])
    defparam i16413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16414_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n25095), 
            .I3(GND_net), .O(n29936));   // verilog/coms.v(127[12] 300[6])
    defparam i16414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16415_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n25095), 
            .I3(GND_net), .O(n29937));   // verilog/coms.v(127[12] 300[6])
    defparam i16415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16416_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n25095), 
            .I3(GND_net), .O(n29938));   // verilog/coms.v(127[12] 300[6])
    defparam i16416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16417_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n25095), 
            .I3(GND_net), .O(n29939));   // verilog/coms.v(127[12] 300[6])
    defparam i16417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16418_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n25095), 
            .I3(GND_net), .O(n29940));   // verilog/coms.v(127[12] 300[6])
    defparam i16418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16419_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n25095), 
            .I3(GND_net), .O(n29941));   // verilog/coms.v(127[12] 300[6])
    defparam i16419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16420_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n25095), 
            .I3(GND_net), .O(n29942));   // verilog/coms.v(127[12] 300[6])
    defparam i16420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16421_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n25095), 
            .I3(GND_net), .O(n29943));   // verilog/coms.v(127[12] 300[6])
    defparam i16421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16422_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n25095), 
            .I3(GND_net), .O(n29944));   // verilog/coms.v(127[12] 300[6])
    defparam i16422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16423_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n25095), 
            .I3(GND_net), .O(n29945));   // verilog/coms.v(127[12] 300[6])
    defparam i16423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16424_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n25095), 
            .I3(GND_net), .O(n29946));   // verilog/coms.v(127[12] 300[6])
    defparam i16424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16425_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n25095), 
            .I3(GND_net), .O(n29947));   // verilog/coms.v(127[12] 300[6])
    defparam i16425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16426_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n25095), 
            .I3(GND_net), .O(n29948));   // verilog/coms.v(127[12] 300[6])
    defparam i16426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16427_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n25095), 
            .I3(GND_net), .O(n29949));   // verilog/coms.v(127[12] 300[6])
    defparam i16427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16428_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n25095), .I3(GND_net), .O(n29950));   // verilog/coms.v(127[12] 300[6])
    defparam i16428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16429_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n25095), .I3(GND_net), .O(n29951));   // verilog/coms.v(127[12] 300[6])
    defparam i16429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16430_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n25095), .I3(GND_net), .O(n29952));   // verilog/coms.v(127[12] 300[6])
    defparam i16430_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1235_15 (.CI(n41119), .I0(n1821), 
            .I1(VCC_net), .CO(n41120));
    SB_LUT4 i16431_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n25095), .I3(GND_net), .O(n29953));   // verilog/coms.v(127[12] 300[6])
    defparam i16431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16432_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n25095), .I3(GND_net), .O(n29954));   // verilog/coms.v(127[12] 300[6])
    defparam i16432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16433_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n25095), .I3(GND_net), .O(n29955));   // verilog/coms.v(127[12] 300[6])
    defparam i16433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16434_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n25095), .I3(GND_net), .O(n29956));   // verilog/coms.v(127[12] 300[6])
    defparam i16434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4605_2_lut (.I0(n2_adj_5167), .I1(encoder0_position[31]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i4605_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16435_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n25095), .I3(GND_net), .O(n29957));   // verilog/coms.v(127[12] 300[6])
    defparam i16435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16436_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n25095), .I3(GND_net), .O(n29958));   // verilog/coms.v(127[12] 300[6])
    defparam i16436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16437_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n25095), .I3(GND_net), .O(n29959));   // verilog/coms.v(127[12] 300[6])
    defparam i16437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16438_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n25095), .I3(GND_net), .O(n29960));   // verilog/coms.v(127[12] 300[6])
    defparam i16438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16439_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n25095), .I3(GND_net), .O(n29961));   // verilog/coms.v(127[12] 300[6])
    defparam i16439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16440_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n25095), .I3(GND_net), .O(n29962));   // verilog/coms.v(127[12] 300[6])
    defparam i16440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16441_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n25095), .I3(GND_net), .O(n29963));   // verilog/coms.v(127[12] 300[6])
    defparam i16441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16442_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n25095), .I3(GND_net), .O(n29964));   // verilog/coms.v(127[12] 300[6])
    defparam i16442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[5]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822), 
            .I2(VCC_net), .I3(n41118), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_14 (.CI(n41118), .I0(n1822), 
            .I1(VCC_net), .CO(n41119));
    SB_LUT4 encoder0_position_31__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n41117), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_8 (.CI(n40893), .I0(n1228), 
            .I1(VCC_net), .CO(n40894));
    SB_CARRY encoder0_position_31__I_0_add_1235_13 (.CI(n41117), .I0(n1823), 
            .I1(VCC_net), .CO(n41118));
    SB_LUT4 i16443_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n25095), .I3(GND_net), .O(n29965));   // verilog/coms.v(127[12] 300[6])
    defparam i16443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16132_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n48426), .I3(GND_net), .O(n29654));   // verilog/coms.v(127[12] 300[6])
    defparam i16132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16444_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n25095), .I3(GND_net), .O(n29966));   // verilog/coms.v(127[12] 300[6])
    defparam i16444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16445_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n25095), .I3(GND_net), .O(n29967));   // verilog/coms.v(127[12] 300[6])
    defparam i16445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16446_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n25095), .I3(GND_net), .O(n29968));   // verilog/coms.v(127[12] 300[6])
    defparam i16446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16447_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n25095), .I3(GND_net), .O(n29969));   // verilog/coms.v(127[12] 300[6])
    defparam i16447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824), 
            .I2(VCC_net), .I3(n41116), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_12 (.CI(n41116), .I0(n1824), 
            .I1(VCC_net), .CO(n41117));
    SB_LUT4 encoder0_position_31__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n41115), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_11 (.CI(n41115), .I0(n1825), 
            .I1(VCC_net), .CO(n41116));
    SB_LUT4 encoder0_position_31__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n41114), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16448_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n25095), .I3(GND_net), .O(n29970));   // verilog/coms.v(127[12] 300[6])
    defparam i16448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16449_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n25095), .I3(GND_net), .O(n29971));   // verilog/coms.v(127[12] 300[6])
    defparam i16449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16450_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n25095), .I3(GND_net), .O(n29972));   // verilog/coms.v(127[12] 300[6])
    defparam i16450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16451_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n25095), .I3(GND_net), .O(n29973));   // verilog/coms.v(127[12] 300[6])
    defparam i16451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16452_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position_scaled[7]), 
            .I2(n25095), .I3(GND_net), .O(n29974));   // verilog/coms.v(127[12] 300[6])
    defparam i16452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16453_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position_scaled[6]), 
            .I2(n25095), .I3(GND_net), .O(n29975));   // verilog/coms.v(127[12] 300[6])
    defparam i16453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16454_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position_scaled[5]), 
            .I2(n25095), .I3(GND_net), .O(n29976));   // verilog/coms.v(127[12] 300[6])
    defparam i16454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16455_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position_scaled[4]), 
            .I2(n25095), .I3(GND_net), .O(n29977));   // verilog/coms.v(127[12] 300[6])
    defparam i16455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16456_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position_scaled[3]), 
            .I2(n25095), .I3(GND_net), .O(n29978));   // verilog/coms.v(127[12] 300[6])
    defparam i16456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37556_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53039));
    defparam i37556_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16457_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position_scaled[2]), 
            .I2(n25095), .I3(GND_net), .O(n29979));   // verilog/coms.v(127[12] 300[6])
    defparam i16457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16458_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position_scaled[1]), 
            .I2(n25095), .I3(GND_net), .O(n29980));   // verilog/coms.v(127[12] 300[6])
    defparam i16458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16459_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position_scaled[0]), 
            .I2(n25095), .I3(GND_net), .O(n29981));   // verilog/coms.v(127[12] 300[6])
    defparam i16459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16460_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position_scaled[15]), 
            .I2(n25095), .I3(GND_net), .O(n29982));   // verilog/coms.v(127[12] 300[6])
    defparam i16460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16461_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position_scaled[14]), 
            .I2(n25095), .I3(GND_net), .O(n29983));   // verilog/coms.v(127[12] 300[6])
    defparam i16461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16462_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position_scaled[13]), 
            .I2(n25095), .I3(GND_net), .O(n29984));   // verilog/coms.v(127[12] 300[6])
    defparam i16462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[6]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16463_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position_scaled[12]), 
            .I2(n25095), .I3(GND_net), .O(n29985));   // verilog/coms.v(127[12] 300[6])
    defparam i16463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16464_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position_scaled[11]), 
            .I2(n25095), .I3(GND_net), .O(n29986));   // verilog/coms.v(127[12] 300[6])
    defparam i16464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16465_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position_scaled[10]), 
            .I2(n25095), .I3(GND_net), .O(n29987));   // verilog/coms.v(127[12] 300[6])
    defparam i16465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16466_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position_scaled[9]), 
            .I2(n25095), .I3(GND_net), .O(n29988));   // verilog/coms.v(127[12] 300[6])
    defparam i16466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16467_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position_scaled[8]), 
            .I2(n25095), .I3(GND_net), .O(n29989));   // verilog/coms.v(127[12] 300[6])
    defparam i16467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16468_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position_scaled[23]), 
            .I2(n25095), .I3(GND_net), .O(n29990));   // verilog/coms.v(127[12] 300[6])
    defparam i16468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16469_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position_scaled[22]), 
            .I2(n25095), .I3(GND_net), .O(n29991));   // verilog/coms.v(127[12] 300[6])
    defparam i16469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16133_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n48426), .I3(GND_net), .O(n29655));   // verilog/coms.v(127[12] 300[6])
    defparam i16133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[7]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16471_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position_scaled[21]), 
            .I2(n25095), .I3(GND_net), .O(n29993));   // verilog/coms.v(127[12] 300[6])
    defparam i16471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16472_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position_scaled[20]), 
            .I2(n25095), .I3(GND_net), .O(n29994));   // verilog/coms.v(127[12] 300[6])
    defparam i16472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16473_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position_scaled[19]), 
            .I2(n25095), .I3(GND_net), .O(n29995));   // verilog/coms.v(127[12] 300[6])
    defparam i16473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5112));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16474_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position_scaled[18]), 
            .I2(n25095), .I3(GND_net), .O(n29996));   // verilog/coms.v(127[12] 300[6])
    defparam i16474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 dti_counter_2056_add_4_9_lut (.I0(n51326), .I1(n35426), .I2(dti_counter[7]), 
            .I3(n41724), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i16475_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position_scaled[17]), 
            .I2(n25095), .I3(GND_net), .O(n29997));   // verilog/coms.v(127[12] 300[6])
    defparam i16475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16476_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position_scaled[16]), 
            .I2(n25095), .I3(GND_net), .O(n29998));   // verilog/coms.v(127[12] 300[6])
    defparam i16476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[8]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16477_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n25095), .I3(GND_net), .O(n29999));   // verilog/coms.v(127[12] 300[6])
    defparam i16477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16478_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n25095), .I3(GND_net), .O(n30000));   // verilog/coms.v(127[12] 300[6])
    defparam i16478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16479_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n25095), .I3(GND_net), .O(n30001));   // verilog/coms.v(127[12] 300[6])
    defparam i16479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16480_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n25095), .I3(GND_net), .O(n30002));   // verilog/coms.v(127[12] 300[6])
    defparam i16480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16481_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n25095), .I3(GND_net), .O(n30003));   // verilog/coms.v(127[12] 300[6])
    defparam i16481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16134_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n48426), .I3(GND_net), .O(n29656));   // verilog/coms.v(127[12] 300[6])
    defparam i16134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16482_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n25095), .I3(GND_net), .O(n30004));   // verilog/coms.v(127[12] 300[6])
    defparam i16482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16483_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n25095), .I3(GND_net), .O(n30005));   // verilog/coms.v(127[12] 300[6])
    defparam i16483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16484_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n25095), .I3(GND_net), .O(n30006));   // verilog/coms.v(127[12] 300[6])
    defparam i16484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16485_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n25095), .I3(GND_net), .O(n30007));   // verilog/coms.v(127[12] 300[6])
    defparam i16485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16486_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n25095), .I3(GND_net), .O(n30008));   // verilog/coms.v(127[12] 300[6])
    defparam i16486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16135_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n48426), .I3(GND_net), .O(n29657));   // verilog/coms.v(127[12] 300[6])
    defparam i16135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16487_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n25095), .I3(GND_net), .O(n30009));   // verilog/coms.v(127[12] 300[6])
    defparam i16487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16488_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n25095), .I3(GND_net), .O(n30010));   // verilog/coms.v(127[12] 300[6])
    defparam i16488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16489_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n25095), .I3(GND_net), .O(n30011));   // verilog/coms.v(127[12] 300[6])
    defparam i16489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37560_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53043));
    defparam i37560_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position[31]), .I3(GND_net), .O(n652));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37594_1_lut (.I0(n36608), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53077));
    defparam i37594_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2196_3_lut (.I0(n3225), .I1(n3292), 
            .I2(n3237), .I3(GND_net), .O(n21_adj_5227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16490_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n25095), .I3(GND_net), .O(n30012));   // verilog/coms.v(127[12] 300[6])
    defparam i16490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2194_3_lut (.I0(n3223), .I1(n3290), 
            .I2(n3237), .I3(GND_net), .O(n25_adj_5229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2191_3_lut (.I0(n3220), .I1(n3287), 
            .I2(n3237), .I3(GND_net), .O(n31_adj_5232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16491_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n25095), .I3(GND_net), .O(n30013));   // verilog/coms.v(127[12] 300[6])
    defparam i16491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1666 (.I0(n3226), .I1(n31_adj_5232), .I2(n3293), 
            .I3(n3237), .O(n48611));
    defparam i1_4_lut_adj_1666.LUT_INIT = 16'heefc;
    SB_LUT4 dti_counter_2056_add_4_8_lut (.I0(n51325), .I1(n35426), .I2(dti_counter[6]), 
            .I3(n41723), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i16492_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n25095), .I3(GND_net), .O(n30014));   // verilog/coms.v(127[12] 300[6])
    defparam i16492_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2056_add_4_8 (.CI(n41723), .I0(n35426), .I1(dti_counter[6]), 
            .CO(n41724));
    SB_LUT4 i16493_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n25095), .I3(GND_net), .O(n30015));   // verilog/coms.v(127[12] 300[6])
    defparam i16493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1667 (.I0(n48611), .I1(n3227), .I2(n3294), .I3(n3237), 
            .O(n48617));
    defparam i1_4_lut_adj_1667.LUT_INIT = 16'heefa;
    SB_LUT4 i16494_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n25095), .I3(GND_net), .O(n30016));   // verilog/coms.v(127[12] 300[6])
    defparam i16494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16495_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n25095), .I3(GND_net), .O(n30017));   // verilog/coms.v(127[12] 300[6])
    defparam i16495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2195_3_lut (.I0(n3224), .I1(n3291), 
            .I2(n3237), .I3(GND_net), .O(n23_adj_5228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16496_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n25095), .I3(GND_net), .O(n30018));   // verilog/coms.v(127[12] 300[6])
    defparam i16496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16497_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n25095), .I3(GND_net), .O(n30019));   // verilog/coms.v(127[12] 300[6])
    defparam i16497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16498_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n25095), .I3(GND_net), .O(n30020));   // verilog/coms.v(127[12] 300[6])
    defparam i16498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16499_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n25095), .I3(GND_net), .O(n30021));   // verilog/coms.v(127[12] 300[6])
    defparam i16499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16500_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n25095), .I3(GND_net), .O(n30022));   // verilog/coms.v(127[12] 300[6])
    defparam i16500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16501_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n25095), .I3(GND_net), .O(n30023));   // verilog/coms.v(127[12] 300[6])
    defparam i16501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16502_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n25095), .I3(GND_net), .O(n30024));   // verilog/coms.v(127[12] 300[6])
    defparam i16502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 dti_counter_2056_add_4_7_lut (.I0(n51324), .I1(n35426), .I2(dti_counter[5]), 
            .I3(n41722), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i16503_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n25095), .I3(GND_net), .O(n30025));   // verilog/coms.v(127[12] 300[6])
    defparam i16503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16504_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n25095), .I3(GND_net), .O(n30026));   // verilog/coms.v(127[12] 300[6])
    defparam i16504_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2056_add_4_7 (.CI(n41722), .I0(n35426), .I1(dti_counter[5]), 
            .CO(n41723));
    SB_LUT4 dti_counter_2056_add_4_6_lut (.I0(n51323), .I1(n35426), .I2(dti_counter[4]), 
            .I3(n41721), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2056_add_4_6 (.CI(n41721), .I0(n35426), .I1(dti_counter[4]), 
            .CO(n41722));
    SB_LUT4 dti_counter_2056_add_4_5_lut (.I0(n51322), .I1(n35426), .I2(dti_counter[3]), 
            .I3(n41720), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2056_add_4_5 (.CI(n41720), .I0(n35426), .I1(dti_counter[3]), 
            .CO(n41721));
    SB_LUT4 dti_counter_2056_add_4_4_lut (.I0(n51321), .I1(n35426), .I2(dti_counter[2]), 
            .I3(n41719), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 encoder0_position_31__I_0_i2193_3_lut (.I0(n3222), .I1(n3289), 
            .I2(n3237), .I3(GND_net), .O(n27_adj_5230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2192_3_lut (.I0(n3221), .I1(n3288), 
            .I2(n3237), .I3(GND_net), .O(n29_adj_5231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16505_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n25095), .I3(GND_net), .O(n30027));   // verilog/coms.v(127[12] 300[6])
    defparam i16505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16506_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n25095), .I3(GND_net), .O(n30028));   // verilog/coms.v(127[12] 300[6])
    defparam i16506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16507_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n25095), .I3(GND_net), .O(n30029));   // verilog/coms.v(127[12] 300[6])
    defparam i16507_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2056_add_4_4 (.CI(n41719), .I0(n35426), .I1(dti_counter[2]), 
            .CO(n41720));
    SB_LUT4 dti_counter_2056_add_4_3_lut (.I0(n51320), .I1(n35426), .I2(dti_counter[1]), 
            .I3(n41718), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2056_add_4_3 (.CI(n41718), .I0(n35426), .I1(dti_counter[1]), 
            .CO(n41719));
    SB_LUT4 dti_counter_2056_add_4_2_lut (.I0(n51311), .I1(n1910), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1235_10 (.CI(n41114), .I0(n1826), 
            .I1(VCC_net), .CO(n41115));
    SB_LUT4 i16508_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n25095), .I3(GND_net), .O(n30030));   // verilog/coms.v(127[12] 300[6])
    defparam i16508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1668 (.I0(n3228), .I1(n21_adj_5227), .I2(n3295), 
            .I3(n3237), .O(n48607));
    defparam i1_4_lut_adj_1668.LUT_INIT = 16'heefc;
    SB_LUT4 i16509_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n25095), 
            .I3(GND_net), .O(n30031));   // verilog/coms.v(127[12] 300[6])
    defparam i16509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16510_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n25095), 
            .I3(GND_net), .O(n30032));   // verilog/coms.v(127[12] 300[6])
    defparam i16510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16511_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n25095), 
            .I3(GND_net), .O(n30033));   // verilog/coms.v(127[12] 300[6])
    defparam i16511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16512_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n25095), 
            .I3(GND_net), .O(n30034));   // verilog/coms.v(127[12] 300[6])
    defparam i16512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16513_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n25095), 
            .I3(GND_net), .O(n30035));   // verilog/coms.v(127[12] 300[6])
    defparam i16513_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2056_add_4_2 (.CI(VCC_net), .I0(n1910), .I1(dti_counter[0]), 
            .CO(n41718));
    SB_LUT4 i16514_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n25095), 
            .I3(GND_net), .O(n30036));   // verilog/coms.v(127[12] 300[6])
    defparam i16514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16515_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n25095), 
            .I3(GND_net), .O(n30037));   // verilog/coms.v(127[12] 300[6])
    defparam i16515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16516_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n25095), 
            .I3(GND_net), .O(n30038));   // verilog/coms.v(127[12] 300[6])
    defparam i16516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16517_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n48426), 
            .I3(GND_net), .O(n30039));   // verilog/coms.v(127[12] 300[6])
    defparam i16517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16518_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n48426), 
            .I3(GND_net), .O(n30040));   // verilog/coms.v(127[12] 300[6])
    defparam i16518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n41113), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16519_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n48426), 
            .I3(GND_net), .O(n30041));   // verilog/coms.v(127[12] 300[6])
    defparam i16519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16520_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n48426), 
            .I3(GND_net), .O(n30042));   // verilog/coms.v(127[12] 300[6])
    defparam i16520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16521_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n48426), 
            .I3(GND_net), .O(n30043));   // verilog/coms.v(127[12] 300[6])
    defparam i16521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1669 (.I0(n29_adj_5231), .I1(n27_adj_5230), .I2(n13_adj_5226), 
            .I3(n23_adj_5228), .O(n48621));
    defparam i1_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1670 (.I0(n48617), .I1(n3218), .I2(n3285), .I3(n3237), 
            .O(n48623));
    defparam i1_4_lut_adj_1670.LUT_INIT = 16'heefa;
    SB_LUT4 i1_4_lut_adj_1671 (.I0(n3219), .I1(n25_adj_5229), .I2(n3286), 
            .I3(n3237), .O(n48615));
    defparam i1_4_lut_adj_1671.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n40892), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1672 (.I0(n48615), .I1(n48623), .I2(n48621), 
            .I3(n48607), .O(n48627));
    defparam i1_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 i22664_4_lut (.I0(n652), .I1(n957), .I2(n3301), .I3(n3237), 
            .O(n36189));
    defparam i22664_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i22842_4_lut (.I0(n36189), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n36372));
    defparam i22842_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i1_4_lut_adj_1673 (.I0(n3217), .I1(n48627), .I2(n3284), .I3(n3237), 
            .O(n48629));
    defparam i1_4_lut_adj_1673.LUT_INIT = 16'heefc;
    SB_LUT4 i16522_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n48426), 
            .I3(GND_net), .O(n30044));   // verilog/coms.v(127[12] 300[6])
    defparam i16522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16523_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n48426), 
            .I3(GND_net), .O(n30045));   // verilog/coms.v(127[12] 300[6])
    defparam i16523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16524_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n48426), 
            .I3(GND_net), .O(n30046));   // verilog/coms.v(127[12] 300[6])
    defparam i16524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16525_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n48426), 
            .I3(GND_net), .O(n30047));   // verilog/coms.v(127[12] 300[6])
    defparam i16525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n51281), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5186));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i1_4_lut_adj_1674 (.I0(n3216), .I1(n48629), .I2(n3283), .I3(n3237), 
            .O(n48631));
    defparam i1_4_lut_adj_1674.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i2186_3_lut (.I0(n3215), .I1(n3282), 
            .I2(n3237), .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2186_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16526_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n48426), 
            .I3(GND_net), .O(n30048));   // verilog/coms.v(127[12] 300[6])
    defparam i16526_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22977_4_lut (.I0(n36372), .I1(n3232), .I2(n3299), .I3(n3237), 
            .O(n36510));
    defparam i22977_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i1_4_lut_adj_1675 (.I0(n36510), .I1(n41), .I2(n48631), .I3(n5_adj_5186), 
            .O(n48635));
    defparam i1_4_lut_adj_1675.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(n3214), .I1(n48635), .I2(n3281), .I3(n3237), 
            .O(n48637));
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'heefc;
    SB_LUT4 i16527_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n48426), 
            .I3(GND_net), .O(n30049));   // verilog/coms.v(127[12] 300[6])
    defparam i16527_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16528_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n48426), 
            .I3(GND_net), .O(n30050));   // verilog/coms.v(127[12] 300[6])
    defparam i16528_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1677 (.I0(n3213), .I1(n48637), .I2(n3280), .I3(n3237), 
            .O(n48639));
    defparam i1_4_lut_adj_1677.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1678 (.I0(n3212), .I1(n48639), .I2(n3279), .I3(n3237), 
            .O(n48641));
    defparam i1_4_lut_adj_1678.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1679 (.I0(n3211), .I1(n48641), .I2(n3278), .I3(n3237), 
            .O(n48643));
    defparam i1_4_lut_adj_1679.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(n3210), .I1(n48643), .I2(n3277), .I3(n3237), 
            .O(n48645));
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1681 (.I0(n3209), .I1(n48645), .I2(n3276), .I3(n3237), 
            .O(n48647));
    defparam i1_4_lut_adj_1681.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1682 (.I0(n3208), .I1(n48647), .I2(n3275), .I3(n3237), 
            .O(n48649));
    defparam i1_4_lut_adj_1682.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(n3207), .I1(n48649), .I2(n3274), .I3(n3237), 
            .O(n48651));
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i2177_3_lut (.I0(n3206), .I1(n3273), 
            .I2(n3237), .I3(GND_net), .O(n59));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2177_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1235_9 (.CI(n41113), .I0(n1827), 
            .I1(VCC_net), .CO(n41114));
    SB_LUT4 encoder0_position_31__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n41112), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16529_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n48426), 
            .I3(GND_net), .O(n30051));   // verilog/coms.v(127[12] 300[6])
    defparam i16529_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16530_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n48426), 
            .I3(GND_net), .O(n30052));   // verilog/coms.v(127[12] 300[6])
    defparam i16530_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_833_7 (.CI(n40892), .I0(n1229), 
            .I1(GND_net), .CO(n40893));
    SB_LUT4 i16531_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n48426), 
            .I3(GND_net), .O(n30053));   // verilog/coms.v(127[12] 300[6])
    defparam i16531_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i37597_4_lut (.I0(n61), .I1(n50106), .I2(n59), .I3(n48651), 
            .O(n36608));
    defparam i37597_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16532_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n48426), 
            .I3(GND_net), .O(n30054));   // verilog/coms.v(127[12] 300[6])
    defparam i16532_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16533_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n48426), 
            .I3(GND_net), .O(n30055));   // verilog/coms.v(127[12] 300[6])
    defparam i16533_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16534_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n48426), 
            .I3(GND_net), .O(n30056));   // verilog/coms.v(127[12] 300[6])
    defparam i16534_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16535_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n48426), 
            .I3(GND_net), .O(n30057));   // verilog/coms.v(127[12] 300[6])
    defparam i16535_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16536_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n48426), 
            .I3(GND_net), .O(n30058));   // verilog/coms.v(127[12] 300[6])
    defparam i16536_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16537_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n48426), 
            .I3(GND_net), .O(n30059));   // verilog/coms.v(127[12] 300[6])
    defparam i16537_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1235_8 (.CI(n41112), .I0(n1828), 
            .I1(VCC_net), .CO(n41113));
    SB_LUT4 encoder0_position_31__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16538_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n48426), 
            .I3(GND_net), .O(n30060));   // verilog/coms.v(127[12] 300[6])
    defparam i16538_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16539_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n48426), 
            .I3(GND_net), .O(n30061));   // verilog/coms.v(127[12] 300[6])
    defparam i16539_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n41111), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16540_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n48426), 
            .I3(GND_net), .O(n30062));   // verilog/coms.v(127[12] 300[6])
    defparam i16540_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16541_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n48426), 
            .I3(GND_net), .O(n30063));   // verilog/coms.v(127[12] 300[6])
    defparam i16541_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230), 
            .I2(GND_net), .I3(n40891), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_7 (.CI(n41111), .I0(n1829), 
            .I1(GND_net), .CO(n41112));
    SB_LUT4 encoder0_position_31__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n41110), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16542_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n48426), 
            .I3(GND_net), .O(n30064));   // verilog/coms.v(127[12] 300[6])
    defparam i16542_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16543_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n48426), 
            .I3(GND_net), .O(n30065));   // verilog/coms.v(127[12] 300[6])
    defparam i16543_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16544_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n48426), 
            .I3(GND_net), .O(n30066));   // verilog/coms.v(127[12] 300[6])
    defparam i16544_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16545_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n48426), 
            .I3(GND_net), .O(n30067));   // verilog/coms.v(127[12] 300[6])
    defparam i16545_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16546_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n48426), 
            .I3(GND_net), .O(n30068));   // verilog/coms.v(127[12] 300[6])
    defparam i16546_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i2_3_lut (.I0(encoder0_position[1]), 
            .I1(n32), .I2(encoder0_position[31]), .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16547_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30069));   // verilog/coms.v(127[12] 300[6])
    defparam i16547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16548_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30070));   // verilog/coms.v(127[12] 300[6])
    defparam i16548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n3221), .I1(n3225), .I2(GND_net), .I3(GND_net), 
            .O(n49225));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16549_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30071));   // verilog/coms.v(127[12] 300[6])
    defparam i16549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16550_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30072));   // verilog/coms.v(127[12] 300[6])
    defparam i16550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16551_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30073));   // verilog/coms.v(127[12] 300[6])
    defparam i16551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n3222), .I1(n3226), .I2(n3223), .I3(n3224), 
            .O(n49231));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n3227), .I1(n49231), .I2(n49225), .I3(n3219), 
            .O(n49235));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 i16552_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30074));   // verilog/coms.v(127[12] 300[6])
    defparam i16552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16553_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30075));   // verilog/coms.v(127[12] 300[6])
    defparam i16553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16554_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30076));   // verilog/coms.v(127[12] 300[6])
    defparam i16554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16555_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30077));   // verilog/coms.v(127[12] 300[6])
    defparam i16555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n3217), .I1(n3218), .I2(n3220), .I3(n3228), 
            .O(n49237));
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'hfffe;
    SB_LUT4 i22846_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n36376));
    defparam i22846_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n3215), .I1(n3216), .I2(n49237), .I3(n49235), 
            .O(n49243));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(n3229), .I1(n36376), .I2(n3230), .I3(n3231), 
            .O(n46818));
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1689 (.I0(n3213), .I1(n3214), .I2(n46818), .I3(n49243), 
            .O(n49249));
    defparam i1_4_lut_adj_1689.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n3210), .I1(n3211), .I2(n3212), .I3(n49249), 
            .O(n49255));
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1691 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n49255), 
            .O(n49261));
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 i37593_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n49261), 
            .O(n3237));
    defparam i37593_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16556_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30078));   // verilog/coms.v(127[12] 300[6])
    defparam i16556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16557_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30079));   // verilog/coms.v(127[12] 300[6])
    defparam i16557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16558_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30080));   // verilog/coms.v(127[12] 300[6])
    defparam i16558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16559_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30081));   // verilog/coms.v(127[12] 300[6])
    defparam i16559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16560_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30082));   // verilog/coms.v(127[12] 300[6])
    defparam i16560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16561_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30083));   // verilog/coms.v(127[12] 300[6])
    defparam i16561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16562_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30084));   // verilog/coms.v(127[12] 300[6])
    defparam i16562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16563_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30085));   // verilog/coms.v(127[12] 300[6])
    defparam i16563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16564_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30086));   // verilog/coms.v(127[12] 300[6])
    defparam i16564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16565_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30087));   // verilog/coms.v(127[12] 300[6])
    defparam i16565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16566_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30088));   // verilog/coms.v(127[12] 300[6])
    defparam i16566_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i3_3_lut (.I0(encoder0_position[2]), 
            .I1(n31), .I2(encoder0_position[31]), .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16567_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30089));   // verilog/coms.v(127[12] 300[6])
    defparam i16567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16568_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30090));   // verilog/coms.v(127[12] 300[6])
    defparam i16568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16569_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30091));   // verilog/coms.v(127[12] 300[6])
    defparam i16569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16570_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30092));   // verilog/coms.v(127[12] 300[6])
    defparam i16570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16571_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30093));   // verilog/coms.v(127[12] 300[6])
    defparam i16571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16572_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30094));   // verilog/coms.v(127[12] 300[6])
    defparam i16572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16573_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30095));   // verilog/coms.v(127[12] 300[6])
    defparam i16573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16574_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30096));   // verilog/coms.v(127[12] 300[6])
    defparam i16574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16575_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30097));   // verilog/coms.v(127[12] 300[6])
    defparam i16575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16576_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30098));   // verilog/coms.v(127[12] 300[6])
    defparam i16576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16577_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30099));   // verilog/coms.v(127[12] 300[6])
    defparam i16577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16578_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n48426), .I3(GND_net), .O(n30100));   // verilog/coms.v(127[12] 300[6])
    defparam i16578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16579_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n48426), .I3(GND_net), .O(n30101));   // verilog/coms.v(127[12] 300[6])
    defparam i16579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16580_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n48426), .I3(GND_net), .O(n30102));   // verilog/coms.v(127[12] 300[6])
    defparam i16580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16581_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n48426), .I3(GND_net), .O(n30103));   // verilog/coms.v(127[12] 300[6])
    defparam i16581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16582_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n48426), .I3(GND_net), .O(n30104));   // verilog/coms.v(127[12] 300[6])
    defparam i16582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16583_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n48426), .I3(GND_net), .O(n30105));   // verilog/coms.v(127[12] 300[6])
    defparam i16583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16584_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n48426), .I3(GND_net), .O(n30106));   // verilog/coms.v(127[12] 300[6])
    defparam i16584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16585_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n48426), .I3(GND_net), .O(n30107));   // verilog/coms.v(127[12] 300[6])
    defparam i16585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n6662), 
            .D(n1103), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1235_6 (.CI(n41110), .I0(n1830), 
            .I1(GND_net), .CO(n41111));
    SB_LUT4 encoder0_position_31__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n41109), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_5 (.CI(n41109), .I0(n1831), 
            .I1(VCC_net), .CO(n41110));
    SB_LUT4 encoder0_position_31__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n41108), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_22 (.CI(n40431), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n40432));
    SB_CARRY encoder0_position_31__I_0_add_1235_4 (.CI(n41108), .I0(n1832), 
            .I1(GND_net), .CO(n41109));
    SB_LUT4 add_224_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n40430), .O(encoder1_position_scaled_23__N_75[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_6 (.CI(n40891), .I0(n1230), 
            .I1(GND_net), .CO(n40892));
    SB_LUT4 i16586_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n48426), .I3(GND_net), .O(n30108));   // verilog/coms.v(127[12] 300[6])
    defparam i16586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231), 
            .I2(VCC_net), .I3(n40890), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_5 (.CI(n40890), .I0(n1231), 
            .I1(VCC_net), .CO(n40891));
    SB_LUT4 i16587_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n48426), .I3(GND_net), .O(n30109));   // verilog/coms.v(127[12] 300[6])
    defparam i16587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16588_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n48426), .I3(GND_net), .O(n30110));   // verilog/coms.v(127[12] 300[6])
    defparam i16588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16589_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n48426), .I3(GND_net), .O(n30111));   // verilog/coms.v(127[12] 300[6])
    defparam i16589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1692 (.I0(n3121), .I1(n3126), .I2(GND_net), .I3(GND_net), 
            .O(n48699));
    defparam i1_2_lut_adj_1692.LUT_INIT = 16'heeee;
    SB_LUT4 i16590_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n48426), .I3(GND_net), .O(n30112));   // verilog/coms.v(127[12] 300[6])
    defparam i16590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1693 (.I0(n3125), .I1(n3122), .I2(n3128), .I3(n3127), 
            .O(n48707));
    defparam i1_4_lut_adj_1693.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1694 (.I0(n3118), .I1(n3119), .I2(n3120), .I3(GND_net), 
            .O(n48711));
    defparam i1_3_lut_adj_1694.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n3123), .I1(n48707), .I2(n48699), .I3(n3124), 
            .O(n48713));
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'hfffe;
    SB_LUT4 i16591_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n48426), .I3(GND_net), .O(n30113));   // verilog/coms.v(127[12] 300[6])
    defparam i16591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n41107), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_21 (.CI(n40430), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n40431));
    SB_CARRY encoder0_position_31__I_0_add_1235_3 (.CI(n41107), .I0(n1833), 
            .I1(VCC_net), .CO(n41108));
    SB_LUT4 add_224_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n40429), .O(encoder1_position_scaled_23__N_75[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22848_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n36378));
    defparam i22848_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i16592_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n48426), .I3(GND_net), .O(n30114));   // verilog/coms.v(127[12] 300[6])
    defparam i16592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_setpoint__i0 (.Q(pwm_setpoint[0]), .C(CLK_c), .D(pwm_setpoint_23__N_191[0]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_CARRY encoder0_position_31__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n41107));
    SB_LUT4 add_2455_25_lut (.I0(n52491), .I1(n2_adj_5194), .I2(n1059), 
            .I3(n41708), .O(encoder0_position_scaled_23__N_51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_25_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_224_8 (.CI(n40417), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n40418));
    SB_LUT4 encoder0_position_31__I_0_add_1168_17_lut (.I0(n52615), .I1(n1719), 
            .I2(VCC_net), .I3(n41106), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1696 (.I0(n3116), .I1(n3117), .I2(n48713), .I3(n48711), 
            .O(n48719));
    defparam i1_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 i16593_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n48426), .I3(GND_net), .O(n30115));   // verilog/coms.v(127[12] 300[6])
    defparam i16593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16594_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n48426), .I3(GND_net), .O(n30116));   // verilog/coms.v(127[12] 300[6])
    defparam i16594_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1697 (.I0(n3129), .I1(n36378), .I2(n3130), .I3(n3131), 
            .O(n46774));
    defparam i1_4_lut_adj_1697.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1698 (.I0(n3114), .I1(n46774), .I2(n3115), .I3(n48719), 
            .O(n48725));
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1699 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n48725), 
            .O(n48731));
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n41105), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_24_lut (.I0(n52505), .I1(n2_adj_5194), .I2(n1158), 
            .I3(n41707), .O(encoder0_position_scaled_23__N_51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n48731), 
            .O(n48737));
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'hfffe;
    SB_CARRY add_2455_24 (.CI(n41707), .I0(n2_adj_5194), .I1(n1158), .CO(n41708));
    SB_LUT4 add_2455_23_lut (.I0(n52520), .I1(n2_adj_5194), .I2(n1257), 
            .I3(n41706), .O(encoder0_position_scaled_23__N_51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i37559_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n48737), 
            .O(n3138));
    defparam i37559_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 add_224_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n40416), .O(encoder1_position_scaled_23__N_75[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2455_23 (.CI(n41706), .I0(n2_adj_5194), .I1(n1257), .CO(n41707));
    SB_LUT4 encoder0_position_31__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2455_22_lut (.I0(n52524), .I1(n2_adj_5194), .I2(n1356), 
            .I3(n41705), .O(encoder0_position_scaled_23__N_51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16595_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n48426), .I3(GND_net), .O(n30117));   // verilog/coms.v(127[12] 300[6])
    defparam i16595_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2455_22 (.CI(n41705), .I0(n2_adj_5194), .I1(n1356), .CO(n41706));
    SB_LUT4 encoder0_position_31__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16596_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n48426), .I3(GND_net), .O(n30118));   // verilog/coms.v(127[12] 300[6])
    defparam i16596_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2455_21_lut (.I0(n52553), .I1(n2_adj_5194), .I2(n1455), 
            .I3(n41704), .O(encoder0_position_scaled_23__N_51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i16597_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n48426), .I3(GND_net), .O(n30119));   // verilog/coms.v(127[12] 300[6])
    defparam i16597_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2455_21 (.CI(n41704), .I0(n2_adj_5194), .I1(n1455), .CO(n41705));
    SB_LUT4 add_2455_20_lut (.I0(n52571), .I1(n2_adj_5194), .I2(n1554), 
            .I3(n41703), .O(encoder0_position_scaled_23__N_51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2455_20 (.CI(n41703), .I0(n2_adj_5194), .I1(n1554), .CO(n41704));
    SB_LUT4 i16598_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n48426), .I3(GND_net), .O(n30120));   // verilog/coms.v(127[12] 300[6])
    defparam i16598_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31064_3_lut (.I0(n5_adj_5164), .I1(n7285), .I2(n46394), .I3(GND_net), 
            .O(n46425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2455_19_lut (.I0(n52590), .I1(n2_adj_5194), .I2(n1653_adj_5183), 
            .I3(n41702), .O(encoder0_position_scaled_23__N_51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_224_20 (.CI(n40429), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n40430));
    SB_LUT4 i16599_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n48426), .I3(GND_net), .O(n30121));   // verilog/coms.v(127[12] 300[6])
    defparam i16599_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2455_19 (.CI(n41702), .I0(n2_adj_5194), .I1(n1653_adj_5183), 
            .CO(n41703));
    SB_LUT4 encoder0_position_31__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2455_18_lut (.I0(n52615), .I1(n2_adj_5194), .I2(n1752), 
            .I3(n41701), .O(encoder0_position_scaled_23__N_51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_18 (.CI(n41701), .I0(n2_adj_5194), .I1(n1752), .CO(n41702));
    SB_LUT4 add_2455_17_lut (.I0(n52641), .I1(n2_adj_5194), .I2(n1851), 
            .I3(n41700), .O(encoder0_position_scaled_23__N_51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_17 (.CI(n41700), .I0(n2_adj_5194), .I1(n1851), .CO(n41701));
    SB_LUT4 i16600_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n48426), .I3(GND_net), .O(n30122));   // verilog/coms.v(127[12] 300[6])
    defparam i16600_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2455_16_lut (.I0(n52665), .I1(n2_adj_5194), .I2(n1950), 
            .I3(n41699), .O(encoder0_position_scaled_23__N_51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2455_16 (.CI(n41699), .I0(n2_adj_5194), .I1(n1950), .CO(n41700));
    SB_LUT4 encoder0_position_31__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16072_3_lut (.I0(n29186), .I1(\ID_READOUT_FSM.state [0]), .I2(n6970), 
            .I3(GND_net), .O(n29594));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16072_3_lut.LUT_INIT = 16'h4646;
    SB_LUT4 add_2455_15_lut (.I0(n52689), .I1(n2_adj_5194), .I2(n2049), 
            .I3(n41698), .O(encoder0_position_scaled_23__N_51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2455_15 (.CI(n41698), .I0(n2_adj_5194), .I1(n2049), .CO(n41699));
    SB_LUT4 encoder0_position_31__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2455_14_lut (.I0(n52719), .I1(n2_adj_5194), .I2(n2148), 
            .I3(n41697), .O(encoder0_position_scaled_23__N_51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i4_3_lut (.I0(encoder0_position[3]), 
            .I1(n30), .I2(encoder0_position[31]), .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2455_14 (.CI(n41697), .I0(n2_adj_5194), .I1(n2148), .CO(n41698));
    SB_LUT4 encoder0_position_31__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232), 
            .I2(GND_net), .I3(n40889), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_13_lut (.I0(n52752), .I1(n2_adj_5194), .I2(n2247), 
            .I3(n41696), .O(encoder0_position_scaled_23__N_51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2455_13 (.CI(n41696), .I0(n2_adj_5194), .I1(n2247), .CO(n41697));
    SB_LUT4 encoder0_position_31__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2455_12_lut (.I0(n52784), .I1(n2_adj_5194), .I2(n2346), 
            .I3(n41695), .O(encoder0_position_scaled_23__N_51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_12 (.CI(n41695), .I0(n2_adj_5194), .I1(n2346), .CO(n41696));
    SB_LUT4 add_2455_11_lut (.I0(n52807), .I1(n2_adj_5194), .I2(n2445), 
            .I3(n41694), .O(encoder0_position_scaled_23__N_51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_16 (.CI(n41105), .I0(n1720), 
            .I1(VCC_net), .CO(n41106));
    SB_LUT4 add_224_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n40428), .O(encoder1_position_scaled_23__N_75[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n41104), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2455_11 (.CI(n41694), .I0(n2_adj_5194), .I1(n2445), .CO(n41695));
    SB_LUT4 add_2455_10_lut (.I0(n52846), .I1(n2_adj_5194), .I2(n2544), 
            .I3(n41693), .O(encoder0_position_scaled_23__N_51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_10 (.CI(n41693), .I0(n2_adj_5194), .I1(n2544), .CO(n41694));
    SB_LUT4 i16603_4_lut (.I0(state_7__N_4103[3]), .I1(data[2]), .I2(n4_adj_5120), 
            .I3(n27911), .O(n30125));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16603_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2455_9_lut (.I0(n52874), .I1(n2_adj_5194), .I2(n2643), 
            .I3(n41692), .O(encoder0_position_scaled_23__N_51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i16060_4_lut (.I0(n29175), .I1(r_Bit_Index[0]), .I2(n45526), 
            .I3(r_SM_Main[1]), .O(n29582));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16060_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 i16056_4_lut (.I0(n29165), .I1(r_Bit_Index_adj_5307[0]), .I2(n45528), 
            .I3(r_SM_Main_adj_5305[1]), .O(n29578));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i16056_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 encoder0_position_31__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1701 (.I0(n6970), .I1(n21721), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n46392));
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'heaee;
    SB_LUT4 i2_4_lut_adj_1702 (.I0(\ID_READOUT_FSM.state [0]), .I1(n35272), 
            .I2(\ID_READOUT_FSM.state [1]), .I3(n46392), .O(n29186));
    defparam i2_4_lut_adj_1702.LUT_INIT = 16'h4c00;
    SB_CARRY add_2455_9 (.CI(n41692), .I0(n2_adj_5194), .I1(n2643), .CO(n41693));
    SB_LUT4 add_2455_8_lut (.I0(n52908), .I1(n2_adj_5194), .I2(n2742), 
            .I3(n41691), .O(encoder0_position_scaled_23__N_51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_8 (.CI(n41691), .I0(n2_adj_5194), .I1(n2742), .CO(n41692));
    SB_CARRY encoder0_position_31__I_0_add_833_4 (.CI(n40889), .I0(n1232), 
            .I1(GND_net), .CO(n40890));
    SB_LUT4 add_2455_7_lut (.I0(n52940), .I1(n2_adj_5194), .I2(n2841), 
            .I3(n41690), .O(encoder0_position_scaled_23__N_51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_224_7 (.CI(n40416), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n40417));
    SB_LUT4 add_224_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n40415), .O(encoder1_position_scaled_23__N_75[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2455_7 (.CI(n41690), .I0(n2_adj_5194), .I1(n2841), .CO(n41691));
    SB_LUT4 add_2455_6_lut (.I0(n52972), .I1(n2_adj_5194), .I2(n2940), 
            .I3(n41689), .O(encoder0_position_scaled_23__N_51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6970), .I2(n29186), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n44751));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(h3), .I1(commutation_state[1]), .I2(h2), 
            .I3(h1), .O(n45417));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'hd054;
    SB_CARRY add_2455_6 (.CI(n41689), .I0(n2_adj_5194), .I1(n2940), .CO(n41690));
    SB_LUT4 i37522_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53005));
    defparam i37522_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n3024), .I1(n3023), .I2(n3021), .I3(n3025), 
            .O(n49187));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n3022), .I1(n3026), .I2(n3027), .I3(n3019), 
            .O(n49185));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1706 (.I0(n49187), .I1(n3020), .I2(n3028), .I3(GND_net), 
            .O(n49189));
    defparam i1_3_lut_adj_1706.LUT_INIT = 16'hfefe;
    SB_LUT4 i22851_3_lut (.I0(n955), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n36382));
    defparam i22851_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233), 
            .I2(VCC_net), .I3(n40888), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_5_lut (.I0(n53005), .I1(n2_adj_5194), .I2(n3039), 
            .I3(n41688), .O(encoder0_position_scaled_23__N_51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_5 (.CI(n41688), .I0(n2_adj_5194), .I1(n3039), .CO(n41689));
    SB_LUT4 add_2455_4_lut (.I0(n53039), .I1(n2_adj_5194), .I2(n3138), 
            .I3(n41687), .O(encoder0_position_scaled_23__N_51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_4 (.CI(n41687), .I0(n2_adj_5194), .I1(n3138), .CO(n41688));
    SB_LUT4 add_2455_3_lut (.I0(n53043), .I1(n2_adj_5194), .I2(n3237), 
            .I3(n41686), .O(encoder0_position_scaled_23__N_51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_3 (.CI(n41686), .I0(n2_adj_5194), .I1(n3237), .CO(n41687));
    SB_LUT4 add_2455_2_lut (.I0(n53077), .I1(n2_adj_5194), .I2(n36608), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_2 (.CI(VCC_net), .I0(n2_adj_5194), .I1(n36608), 
            .CO(n41686));
    SB_LUT4 encoder0_position_31__I_0_add_2173_33_lut (.I0(n53043), .I1(n3204), 
            .I2(VCC_net), .I3(n41685), .O(n50106)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n41684), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_32 (.CI(n41684), .I0(n3205), 
            .I1(VCC_net), .CO(n41685));
    SB_LUT4 encoder0_position_31__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n41683), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_31 (.CI(n41683), .I0(n3206), 
            .I1(VCC_net), .CO(n41684));
    SB_LUT4 encoder0_position_31__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n41682), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_30 (.CI(n41682), .I0(n3207), 
            .I1(VCC_net), .CO(n41683));
    SB_LUT4 encoder0_position_31__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n41681), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_29 (.CI(n41681), .I0(n3208), 
            .I1(VCC_net), .CO(n41682));
    SB_LUT4 encoder0_position_31__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n41680), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_28 (.CI(n41680), .I0(n3209), 
            .I1(VCC_net), .CO(n41681));
    SB_LUT4 encoder0_position_31__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n41679), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_15 (.CI(n41104), .I0(n1721), 
            .I1(VCC_net), .CO(n41105));
    SB_LUT4 i1_4_lut_adj_1707 (.I0(n3017), .I1(n3018), .I2(n49189), .I3(n49185), 
            .O(n49195));
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1708 (.I0(n3029), .I1(n36382), .I2(n3030), .I3(n3031), 
            .O(n46814));
    defparam i1_4_lut_adj_1708.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n3015), .I1(n46814), .I2(n3016), .I3(n49195), 
            .O(n49201));
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1710 (.I0(n3012), .I1(n3013), .I2(n3014), .I3(n49201), 
            .O(n49207));
    defparam i1_4_lut_adj_1710.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_2173_27 (.CI(n41679), .I0(n3210), 
            .I1(VCC_net), .CO(n41680));
    SB_LUT4 encoder0_position_31__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n41678), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n49207), 
            .O(n49213));
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_2173_26 (.CI(n41678), .I0(n3211), 
            .I1(VCC_net), .CO(n41679));
    SB_LUT4 encoder0_position_31__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n41677), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37363_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52846));
    defparam i37363_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37525_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n49213), 
            .O(n3039));
    defparam i37525_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_25 (.CI(n41677), .I0(n3212), 
            .I1(VCC_net), .CO(n41678));
    SB_LUT4 encoder0_position_31__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n41103), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n41676), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_24 (.CI(n41676), .I0(n3213), 
            .I1(VCC_net), .CO(n41677));
    SB_LUT4 i37391_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52874));
    defparam i37391_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n41675), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_23 (.CI(n41675), .I0(n3214), 
            .I1(VCC_net), .CO(n41676));
    SB_LUT4 encoder0_position_31__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n41674), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_22 (.CI(n41674), .I0(n3215), 
            .I1(VCC_net), .CO(n41675));
    SB_LUT4 encoder0_position_31__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n41673), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_21 (.CI(n41673), .I0(n3216), 
            .I1(VCC_net), .CO(n41674));
    SB_CARRY encoder0_position_31__I_0_add_833_3 (.CI(n40888), .I0(n1233), 
            .I1(VCC_net), .CO(n40889));
    SB_LUT4 encoder0_position_31__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n41672), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_20 (.CI(n41672), .I0(n3217), 
            .I1(VCC_net), .CO(n41673));
    SB_LUT4 encoder0_position_31__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n41671), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n40888));
    SB_CARRY encoder0_position_31__I_0_add_2173_19 (.CI(n41671), .I0(n3218), 
            .I1(VCC_net), .CO(n41672));
    SB_LUT4 encoder0_position_31__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n41670), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[16]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_18 (.CI(n41670), .I0(n3219), 
            .I1(VCC_net), .CO(n41671));
    SB_LUT4 encoder0_position_31__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n41669), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_add_2173_17 (.CI(n41669), .I0(n3220), 
            .I1(VCC_net), .CO(n41670));
    SB_LUT4 encoder0_position_31__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n41668), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_16 (.CI(n41668), .I0(n3221), 
            .I1(VCC_net), .CO(n41669));
    SB_LUT4 encoder0_position_31__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n41667), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_15 (.CI(n41667), .I0(n3222), 
            .I1(VCC_net), .CO(n41668));
    SB_LUT4 encoder0_position_31__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n41666), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_14 (.CI(n41666), .I0(n3223), 
            .I1(VCC_net), .CO(n41667));
    SB_LUT4 encoder0_position_31__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_224_19 (.CI(n40428), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n40429));
    SB_LUT4 encoder0_position_31__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n41665), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i5_3_lut (.I0(encoder0_position[4]), 
            .I1(n29), .I2(encoder0_position[31]), .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_13 (.CI(n41665), .I0(n3224), 
            .I1(VCC_net), .CO(n41666));
    SB_LUT4 encoder0_position_31__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n41664), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37489_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52972));
    defparam i37489_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1712 (.I0(n2920), .I1(n2926), .I2(GND_net), .I3(GND_net), 
            .O(n49083));
    defparam i1_2_lut_adj_1712.LUT_INIT = 16'heeee;
    SB_LUT4 i22853_3_lut (.I0(n954), .I1(n2932), .I2(n2933), .I3(GND_net), 
            .O(n36384));
    defparam i22853_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(n2927), .I1(n2928), .I2(n2923), .I3(n2925), 
            .O(n48673));
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1714 (.I0(n2918), .I1(n49083), .I2(n2919), .I3(n2922), 
            .O(n49089));
    defparam i1_4_lut_adj_1714.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1715 (.I0(n2929), .I1(n36384), .I2(n2930), .I3(n2931), 
            .O(n46765));
    defparam i1_4_lut_adj_1715.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n2916), .I1(n48673), .I2(n2921), .I3(n2924), 
            .O(n48677));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_2173_12 (.CI(n41664), .I0(n3225), 
            .I1(VCC_net), .CO(n41665));
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n2917), .I1(n48677), .I2(n46765), .I3(n49089), 
            .O(n48679));
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n41663), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_11 (.CI(n41663), .I0(n3226), 
            .I1(VCC_net), .CO(n41664));
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n2913), .I1(n2914), .I2(n48679), .I3(n2915), 
            .O(n48685));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'hfffe;
    SB_LUT4 add_224_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n40427), .O(encoder1_position_scaled_23__N_75[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31065_3_lut (.I0(encoder0_position[28]), .I1(n46425), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1719 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n48685), 
            .O(n48691));
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'hfffe;
    SB_LUT4 i37492_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n48691), 
            .O(n2940));
    defparam i37492_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n41662), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_10 (.CI(n41662), .I0(n3227), 
            .I1(VCC_net), .CO(n41663));
    SB_LUT4 encoder0_position_31__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n41661), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_9 (.CI(n41661), .I0(n3228), 
            .I1(VCC_net), .CO(n41662));
    SB_LUT4 encoder0_position_31__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n41660), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_8 (.CI(n41660), .I0(n3229), 
            .I1(GND_net), .CO(n41661));
    SB_LUT4 encoder0_position_31__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i6_3_lut (.I0(encoder0_position[5]), 
            .I1(n28), .I2(encoder0_position[31]), .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36494_3_lut (.I0(n2624), .I1(n2691), .I2(n2643), .I3(GND_net), 
            .O(n2723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36494_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36495_3_lut (.I0(n2723), .I1(n2790), .I2(n2742), .I3(GND_net), 
            .O(n2822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36495_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36498_3_lut (.I0(n2627), .I1(n2694), .I2(n2643), .I3(GND_net), 
            .O(n2726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36498_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36499_3_lut (.I0(n2726), .I1(n2793), .I2(n2742), .I3(GND_net), 
            .O(n2825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36499_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36496_3_lut (.I0(n2626), .I1(n2693), .I2(n2643), .I3(GND_net), 
            .O(n2725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36496_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36497_3_lut (.I0(n2725), .I1(n2792), .I2(n2742), .I3(GND_net), 
            .O(n2824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36497_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36500_3_lut (.I0(n2628), .I1(n2695), .I2(n2643), .I3(GND_net), 
            .O(n2727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36500_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36501_3_lut (.I0(n2727), .I1(n2794), .I2(n2742), .I3(GND_net), 
            .O(n2826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36501_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i37457_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52940));
    defparam i37457_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16065_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_5101), 
            .I3(n27903), .O(n29587));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16065_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n2826), .I1(n2823), .I2(n2821), .I3(n2828), 
            .O(n49103));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1721 (.I0(n49103), .I1(n2822), .I2(n2827), .I3(GND_net), 
            .O(n49105));
    defparam i1_3_lut_adj_1721.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n2819), .I1(n2824), .I2(n2825), .I3(n2820), 
            .O(n49107));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'hfffe;
    SB_LUT4 i22987_4_lut (.I0(n953), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n36520));
    defparam i22987_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(n2817), .I1(n2818), .I2(n49107), .I3(n49105), 
            .O(n49113));
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n2829), .I1(n49113), .I2(n36520), .I3(n2830), 
            .O(n49115));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n2814), .I1(n2815), .I2(n2816), .I3(n49115), 
            .O(n49121));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n41659), .O(n51281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n49121), 
            .O(n49127));
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 i37460_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n49127), 
            .O(n2841));
    defparam i37460_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_7 (.CI(n41659), .I0(n3230), 
            .I1(GND_net), .CO(n41660));
    SB_LUT4 encoder0_position_31__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n41658), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_6 (.CI(n41658), .I0(n3231), 
            .I1(VCC_net), .CO(n41659));
    SB_LUT4 encoder0_position_31__I_0_add_2173_5_lut (.I0(GND_net), .I1(n3232), 
            .I2(GND_net), .I3(n41657), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_5 (.CI(n41657), .I0(n3232), 
            .I1(GND_net), .CO(n41658));
    SB_LUT4 encoder0_position_31__I_0_add_2173_4_lut (.I0(GND_net), .I1(n3233), 
            .I2(VCC_net), .I3(n41656), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_4 (.CI(n41656), .I0(n3233), 
            .I1(VCC_net), .CO(n41657));
    SB_LUT4 encoder0_position_31__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14_3_lut (.I0(h2), .I1(h3), .I2(h1), .I3(GND_net), .O(n6_adj_5189));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1727 (.I0(h3), .I1(h2), .I2(h1), .I3(GND_net), 
            .O(commutation_state_7__N_216[0]));   // verilog/TinyFPGA_B.v(148[4] 150[7])
    defparam i1_3_lut_adj_1727.LUT_INIT = 16'h1414;
    SB_LUT4 encoder0_position_31__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i7_3_lut (.I0(encoder0_position[6]), 
            .I1(n27), .I2(encoder0_position[31]), .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n41655), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_3 (.CI(n41655), .I0(n957), 
            .I1(GND_net), .CO(n41656));
    SB_CARRY encoder0_position_31__I_0_add_2173_2 (.CI(VCC_net), .I0(n652), 
            .I1(VCC_net), .CO(n41655));
    SB_LUT4 encoder0_position_31__I_0_add_2106_31_lut (.I0(n53039), .I1(n3105), 
            .I2(VCC_net), .I3(n41654), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n41653), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_30 (.CI(n41653), .I0(n3106), 
            .I1(VCC_net), .CO(n41654));
    SB_LUT4 encoder0_position_31__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n41652), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_29 (.CI(n41652), .I0(n3107), 
            .I1(VCC_net), .CO(n41653));
    SB_LUT4 encoder0_position_31__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n41651), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_28 (.CI(n41651), .I0(n3108), 
            .I1(VCC_net), .CO(n41652));
    SB_LUT4 encoder0_position_31__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n41650), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_27 (.CI(n41650), .I0(n3109), 
            .I1(VCC_net), .CO(n41651));
    SB_CARRY encoder0_position_31__I_0_add_1168_14 (.CI(n41103), .I0(n1722), 
            .I1(VCC_net), .CO(n41104));
    SB_LUT4 encoder0_position_31__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n41649), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36769_3_lut (.I0(n2522), .I1(n2589), .I2(n2544), .I3(GND_net), 
            .O(n2621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36769_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_26 (.CI(n41649), .I0(n3110), 
            .I1(VCC_net), .CO(n41650));
    SB_LUT4 i36711_3_lut (.I0(n2621), .I1(n2688), .I2(n2643), .I3(GND_net), 
            .O(n2720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n41648), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_25 (.CI(n41648), .I0(n3111), 
            .I1(VCC_net), .CO(n41649));
    SB_CARRY add_224_18 (.CI(n40427), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n40428));
    SB_LUT4 i36767_3_lut (.I0(n2524), .I1(n2591), .I2(n2544), .I3(GND_net), 
            .O(n2623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36767_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36713_3_lut (.I0(n2623), .I1(n2690), .I2(n2643), .I3(GND_net), 
            .O(n2722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n41647), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i37425_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52908));
    defparam i37425_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1728 (.I0(n2727), .I1(n2725), .I2(GND_net), .I3(GND_net), 
            .O(n48815));
    defparam i1_2_lut_adj_1728.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(n2724), .I1(n2721), .I2(n2722), .I3(n2728), 
            .O(n48817));
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(n2723), .I1(n2720), .I2(n48815), .I3(n2726), 
            .O(n48821));
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'hfffe;
    SB_LUT4 i22989_4_lut (.I0(n952), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n36522));
    defparam i22989_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1731 (.I0(n2718), .I1(n2719), .I2(n48821), .I3(n48817), 
            .O(n48827));
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n2729), .I1(n48827), .I2(n36522), .I3(n2730), 
            .O(n48829));
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1733 (.I0(n2715), .I1(n2716), .I2(n48829), .I3(n2717), 
            .O(n48835));
    defparam i1_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1734 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n48835), 
            .O(n48841));
    defparam i1_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i37429_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n48841), 
            .O(n2742));
    defparam i37429_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY add_145_13 (.CI(n40391), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n40392));
    SB_LUT4 encoder0_position_31__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n41102), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_24 (.CI(n41647), .I0(n3112), 
            .I1(VCC_net), .CO(n41648));
    SB_LUT4 encoder0_position_31__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n41646), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_23 (.CI(n41646), .I0(n3113), 
            .I1(VCC_net), .CO(n41647));
    SB_LUT4 encoder0_position_31__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_13 (.CI(n41102), .I0(n1723), 
            .I1(VCC_net), .CO(n41103));
    SB_LUT4 i16136_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n48426), .I3(GND_net), .O(n29658));   // verilog/coms.v(127[12] 300[6])
    defparam i16136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n41645), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_22 (.CI(n41645), .I0(n3114), 
            .I1(VCC_net), .CO(n41646));
    SB_LUT4 encoder0_position_31__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n41644), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16137_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n48426), .I3(GND_net), .O(n29659));   // verilog/coms.v(127[12] 300[6])
    defparam i16137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_21 (.CI(n41644), .I0(n3115), 
            .I1(VCC_net), .CO(n41645));
    SB_LUT4 encoder0_position_31__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n41101), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_12 (.CI(n41101), .I0(n1724), 
            .I1(VCC_net), .CO(n41102));
    SB_LUT4 encoder0_position_31__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n41643), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5111));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2106_20 (.CI(n41643), .I0(n3116), 
            .I1(VCC_net), .CO(n41644));
    SB_LUT4 encoder0_position_31__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i17_3_lut (.I0(encoder0_position[16]), 
            .I1(n17), .I2(encoder0_position[31]), .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n41100), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n41642), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_19 (.CI(n41642), .I0(n3117), 
            .I1(VCC_net), .CO(n41643));
    SB_CARRY encoder0_position_31__I_0_add_1168_11 (.CI(n41100), .I0(n1725), 
            .I1(VCC_net), .CO(n41101));
    SB_LUT4 encoder0_position_31__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n41641), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n41099), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_10 (.CI(n41099), .I0(n1726), 
            .I1(VCC_net), .CO(n41100));
    SB_LUT4 encoder0_position_31__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n40426), .O(encoder1_position_scaled_23__N_75[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36655_3_lut (.I0(n51971), .I1(n2490), .I2(n2445), .I3(GND_net), 
            .O(n2522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36655_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_18 (.CI(n41641), .I0(n3118), 
            .I1(VCC_net), .CO(n41642));
    SB_LUT4 encoder0_position_31__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n41640), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_17 (.CI(n40426), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n40427));
    SB_LUT4 encoder0_position_31__I_0_i1721_rep_18_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1721_rep_18_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_17 (.CI(n41640), .I0(n3119), 
            .I1(VCC_net), .CO(n41641));
    SB_LUT4 encoder0_position_31__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n41639), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_16 (.CI(n41639), .I0(n3120), 
            .I1(VCC_net), .CO(n41640));
    SB_LUT4 add_224_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n40425), .O(encoder1_position_scaled_23__N_75[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n41638), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_15 (.CI(n41638), .I0(n3121), 
            .I1(VCC_net), .CO(n41639));
    SB_LUT4 encoder0_position_31__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n41098), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n41637), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_14 (.CI(n41637), .I0(n3122), 
            .I1(VCC_net), .CO(n41638));
    SB_CARRY add_224_16 (.CI(n40425), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n40426));
    SB_LUT4 encoder0_position_31__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n41636), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_13 (.CI(n41636), .I0(n3123), 
            .I1(VCC_net), .CO(n41637));
    SB_CARRY add_224_6 (.CI(n40415), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n40416));
    SB_LUT4 add_224_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n40424), .O(encoder1_position_scaled_23__N_75[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n41635), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_12 (.CI(n41635), .I0(n3124), 
            .I1(VCC_net), .CO(n41636));
    SB_LUT4 encoder0_position_31__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n40414), .O(encoder1_position_scaled_23__N_75[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_9 (.CI(n41098), .I0(n1727), 
            .I1(VCC_net), .CO(n41099));
    SB_LUT4 encoder0_position_31__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i8_3_lut (.I0(encoder0_position[7]), 
            .I1(n26), .I2(encoder0_position[31]), .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1718_rep_19_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1718_rep_19_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n41634), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1720_rep_11_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1720_rep_11_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n6662), 
            .D(n1102), .R(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_2106_11 (.CI(n41634), .I0(n3125), 
            .I1(VCC_net), .CO(n41635));
    SB_LUT4 encoder0_position_31__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n41633), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_10 (.CI(n41633), .I0(n3126), 
            .I1(VCC_net), .CO(n41634));
    SB_LUT4 i36653_3_lut (.I0(n51973), .I1(n2492), .I2(n2445), .I3(GND_net), 
            .O(n2524));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n41632), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_9 (.CI(n41632), .I0(n3127), 
            .I1(VCC_net), .CO(n41633));
    SB_LUT4 encoder0_position_31__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n41631), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_8 (.CI(n41631), .I0(n3128), 
            .I1(VCC_net), .CO(n41632));
    SB_LUT4 encoder0_position_31__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n41630), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1735 (.I0(n2626), .I1(n2625), .I2(GND_net), .I3(GND_net), 
            .O(n49135));
    defparam i1_2_lut_adj_1735.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(n2623), .I1(n2624), .I2(n2622), .I3(n2627), 
            .O(n49143));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_2106_7 (.CI(n41630), .I0(n3129), 
            .I1(GND_net), .CO(n41631));
    SB_LUT4 encoder0_position_31__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n41629), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_5 (.CI(n40414), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n40415));
    SB_LUT4 add_224_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n40413), .O(encoder1_position_scaled_23__N_75[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n2628), .I1(n49143), .I2(n49135), .I3(n2621), 
            .O(n49145));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hfffe;
    SB_CARRY add_224_15 (.CI(n40424), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n40425));
    SB_LUT4 i22866_3_lut (.I0(n951), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n36398));
    defparam i22866_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_31__I_0_add_2106_6 (.CI(n41629), .I0(n3130), 
            .I1(GND_net), .CO(n41630));
    SB_CARRY add_224_4 (.CI(n40413), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n40414));
    SB_LUT4 i1_4_lut_adj_1738 (.I0(n2618), .I1(n2619), .I2(n49145), .I3(n2620), 
            .O(n49151));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n41628), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1739 (.I0(n2629), .I1(n36398), .I2(n2630), .I3(n2631), 
            .O(n46786));
    defparam i1_4_lut_adj_1739.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_add_766_11_lut (.I0(n52505), .I1(n1125), 
            .I2(VCC_net), .I3(n40788), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n41097), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1740 (.I0(n2616), .I1(n2617), .I2(n46786), .I3(n49151), 
            .O(n49157));
    defparam i1_4_lut_adj_1740.LUT_INIT = 16'hfffe;
    SB_LUT4 add_224_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n40412), .O(encoder1_position_scaled_23__N_75[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1741 (.I0(n2613), .I1(n2614), .I2(n2615), .I3(n49157), 
            .O(n49163));
    defparam i1_4_lut_adj_1741.LUT_INIT = 16'hfffe;
    SB_LUT4 i37399_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n49163), 
            .O(n2643));
    defparam i37399_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_8 (.CI(n41097), .I0(n1728), 
            .I1(VCC_net), .CO(n41098));
    SB_CARRY encoder0_position_31__I_0_add_2106_5 (.CI(n41628), .I0(n3131), 
            .I1(VCC_net), .CO(n41629));
    SB_LUT4 encoder0_position_31__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n40787), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_766_10 (.CI(n40787), .I0(n1126), 
            .I1(VCC_net), .CO(n40788));
    SB_CARRY add_224_3 (.CI(n40412), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n40413));
    SB_LUT4 encoder0_position_31__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n41627), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_4 (.CI(n41627), .I0(n3132), 
            .I1(GND_net), .CO(n41628));
    SB_LUT4 encoder0_position_31__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n41096), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_7 (.CI(n41096), .I0(n1729), 
            .I1(GND_net), .CO(n41097));
    SB_LUT4 add_224_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n40423), .O(encoder1_position_scaled_23__N_75[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_14_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n41626), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_3 (.CI(n41626), .I0(n3133), 
            .I1(VCC_net), .CO(n41627));
    SB_LUT4 encoder0_position_31__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n41095), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n40786), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n41626));
    SB_LUT4 encoder0_position_31__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_766_9 (.CI(n40786), .I0(n1127), 
            .I1(VCC_net), .CO(n40787));
    SB_LUT4 encoder0_position_31__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n40785), .O(n1195_adj_5182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_6 (.CI(n41095), .I0(n1730), 
            .I1(GND_net), .CO(n41096));
    SB_LUT4 encoder0_position_31__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i9_3_lut (.I0(encoder0_position[8]), 
            .I1(n25), .I2(encoder0_position[31]), .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2), .I3(n40695), .O(displacement_23__N_99[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1451_rep_64_3_lut (.I0(n2195), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n50236));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1451_rep_64_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1518_rep_48_3_lut (.I0(n50236), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n50220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1518_rep_48_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_30_lut (.I0(n53005), .I1(n3006), 
            .I2(VCC_net), .I3(n41625), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i36340_3_lut (.I0(n2346), .I1(n2247), .I2(n2148), .I3(GND_net), 
            .O(n51822));
    defparam i36340_3_lut.LUT_INIT = 16'h7f7f;
    SB_LUT4 encoder0_position_31__I_0_i1449_rep_56_3_lut (.I0(n2193), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n50228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1449_rep_56_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n41624), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_29 (.CI(n41624), .I0(n3007), 
            .I1(VCC_net), .CO(n41625));
    SB_LUT4 encoder0_position_31__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n41623), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_28 (.CI(n41623), .I0(n3008), 
            .I1(VCC_net), .CO(n41624));
    SB_LUT4 encoder0_position_31__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n41622), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_27 (.CI(n41622), .I0(n3009), 
            .I1(VCC_net), .CO(n41623));
    SB_LUT4 encoder0_position_31__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n41621), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_26 (.CI(n41621), .I0(n3010), 
            .I1(VCC_net), .CO(n41622));
    SB_LUT4 encoder0_position_31__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n41620), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_25 (.CI(n41620), .I0(n3011), 
            .I1(VCC_net), .CO(n41621));
    SB_LUT4 encoder0_position_31__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n41094), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n41619), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_24 (.CI(n41619), .I0(n3012), 
            .I1(VCC_net), .CO(n41620));
    SB_CARRY encoder0_position_31__I_0_add_1168_5 (.CI(n41094), .I0(n1731), 
            .I1(VCC_net), .CO(n41095));
    SB_LUT4 encoder0_position_31__I_0_i1516_rep_40_3_lut (.I0(n50228), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n50212));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1516_rep_40_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n41618), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_23 (.CI(n41618), .I0(n3013), 
            .I1(VCC_net), .CO(n41619));
    SB_LUT4 encoder0_position_31__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n41617), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36488_3_lut (.I0(n50212), .I1(n2126), .I2(n51822), .I3(GND_net), 
            .O(n51971));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36488_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_22 (.CI(n41617), .I0(n3014), 
            .I1(VCC_net), .CO(n41618));
    SB_LUT4 encoder0_position_31__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n41616), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_21 (.CI(n41616), .I0(n3015), 
            .I1(VCC_net), .CO(n41617));
    SB_LUT4 encoder0_position_31__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n41615), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_20 (.CI(n41615), .I0(n3016), 
            .I1(VCC_net), .CO(n41616));
    SB_LUT4 encoder0_position_31__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n41093), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36490_3_lut (.I0(n50220), .I1(n2128), .I2(n51822), .I3(GND_net), 
            .O(n51973));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36490_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n41614), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_8 (.CI(n40785), .I0(n1128), 
            .I1(VCC_net), .CO(n40786));
    SB_CARRY encoder0_position_31__I_0_add_1168_4 (.CI(n41093), .I0(n1732), 
            .I1(GND_net), .CO(n41094));
    SB_LUT4 encoder0_position_31__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_19 (.CI(n41614), .I0(n3017), 
            .I1(VCC_net), .CO(n41615));
    SB_LUT4 i36771_3_lut (.I0(n2325), .I1(n2392), .I2(n2346), .I3(GND_net), 
            .O(n2424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5148), .I3(n40694), .O(displacement_23__N_99[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36709_3_lut (.I0(n2424), .I1(n2491), .I2(n2445), .I3(GND_net), 
            .O(n2523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n41613), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_5110));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2039_18 (.CI(n41613), .I0(n3018), 
            .I1(VCC_net), .CO(n41614));
    SB_LUT4 encoder0_position_31__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n41612), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36275_3_lut (.I0(n2426), .I1(n2493), .I2(n2445), .I3(GND_net), 
            .O(n2525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36275_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_17 (.CI(n41612), .I0(n3019), 
            .I1(VCC_net), .CO(n41613));
    SB_LUT4 i36492_3_lut (.I0(n2328), .I1(n2395), .I2(n2346), .I3(GND_net), 
            .O(n2427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36492_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n41611), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36493_3_lut (.I0(n2427), .I1(n2494), .I2(n2445), .I3(GND_net), 
            .O(n2526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36493_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1742 (.I0(n2526), .I1(n2525), .I2(n2523), .I3(n2528), 
            .O(n48581));
    defparam i1_4_lut_adj_1742.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1743 (.I0(n2524), .I1(n2521), .I2(n2527), .I3(n2522), 
            .O(n48583));
    defparam i1_4_lut_adj_1743.LUT_INIT = 16'hfffe;
    SB_LUT4 i22870_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n36402));
    defparam i22870_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n40784), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(n2519), .I1(n2520), .I2(n48583), .I3(n48581), 
            .O(n48589));
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1745 (.I0(n2529), .I1(n36402), .I2(n2530), .I3(n2531), 
            .O(n46745));
    defparam i1_4_lut_adj_1745.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1746 (.I0(n2517), .I1(n46745), .I2(n2518), .I3(n48589), 
            .O(n48595));
    defparam i1_4_lut_adj_1746.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_2039_16 (.CI(n41611), .I0(n3020), 
            .I1(VCC_net), .CO(n41612));
    SB_LUT4 encoder0_position_31__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n41610), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_15 (.CI(n41610), .I0(n3021), 
            .I1(VCC_net), .CO(n41611));
    SB_LUT4 encoder0_position_31__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n41609), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1747 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n48595), 
            .O(n48601));
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'hfffe;
    SB_LUT4 i37366_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n48601), 
            .O(n2544));
    defparam i37366_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_2039_14 (.CI(n41609), .I0(n3022), 
            .I1(VCC_net), .CO(n41610));
    SB_LUT4 encoder0_position_31__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n41608), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_13 (.CI(n41608), .I0(n3023), 
            .I1(VCC_net), .CO(n41609));
    SB_LUT4 encoder0_position_31__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n41607), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_12 (.CI(n41607), .I0(n3024), 
            .I1(VCC_net), .CO(n41608));
    SB_LUT4 encoder0_position_31__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n41606), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_11 (.CI(n41606), .I0(n3025), 
            .I1(VCC_net), .CO(n41607));
    SB_LUT4 encoder0_position_31__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n41605), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_10 (.CI(n41605), .I0(n3026), 
            .I1(VCC_net), .CO(n41606));
    SB_LUT4 encoder0_position_31__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n41604), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_9 (.CI(n41604), .I0(n3027), 
            .I1(VCC_net), .CO(n41605));
    SB_LUT4 encoder0_position_31__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n41603), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_8 (.CI(n41603), .I0(n3028), 
            .I1(VCC_net), .CO(n41604));
    SB_LUT4 encoder0_position_31__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n41602), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_7 (.CI(n41602), .I0(n3029), 
            .I1(GND_net), .CO(n41603));
    SB_LUT4 encoder0_position_31__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n41601), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_224_14 (.CI(n40423), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n40424));
    SB_LUT4 encoder0_position_31__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_6 (.CI(n41601), .I0(n3030), 
            .I1(GND_net), .CO(n41602));
    SB_LUT4 encoder0_position_31__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n41600), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_5 (.CI(n41600), .I0(n3031), 
            .I1(VCC_net), .CO(n41601));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i10_3_lut (.I0(encoder0_position[9]), 
            .I1(n24), .I2(encoder0_position[31]), .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1519_rep_51_3_lut (.I0(n2295), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n50223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1519_rep_51_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1588_rep_35_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1588_rep_35_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n41599), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_4 (.CI(n41599), .I0(n3032), 
            .I1(GND_net), .CO(n41600));
    SB_LUT4 encoder0_position_31__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n41598), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_3 (.CI(n41598), .I0(n3033), 
            .I1(VCC_net), .CO(n41599));
    SB_LUT4 encoder0_position_31__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n41092), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_3 (.CI(n41092), .I0(n1733), 
            .I1(VCC_net), .CO(n41093));
    SB_CARRY encoder0_position_31__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n41598));
    SB_LUT4 encoder0_position_31__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n40422), .O(encoder1_position_scaled_23__N_75[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_13 (.CI(n40422), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n40423));
    SB_LUT4 encoder0_position_31__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_7 (.CI(n40784), .I0(n1129), 
            .I1(GND_net), .CO(n40785));
    SB_LUT4 add_224_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_279), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n40694), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5148), .CO(n40695));
    SB_LUT4 i36659_3_lut (.I0(n2225), .I1(n2292), .I2(n2247), .I3(GND_net), 
            .O(n2324));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5109));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36611_3_lut (.I0(n2324), .I1(n2391), .I2(n2346), .I3(GND_net), 
            .O(n2423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36611_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5147), .I3(n40693), .O(displacement_23__N_99[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36657_3_lut (.I0(n2227), .I1(n2294), .I2(n2247), .I3(GND_net), 
            .O(n2326));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36615_3_lut (.I0(n2326), .I1(n2393), .I2(n2346), .I3(GND_net), 
            .O(n2425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36615_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_DFFSR pwm_setpoint__i23 (.Q(pwm_setpoint[23]), .C(CLK_c), .D(pwm_setpoint_23__N_191[23]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 i1_4_lut_adj_1748 (.I0(n2423), .I1(n2424), .I2(n2426), .I3(n2428), 
            .O(n49053));
    defparam i1_4_lut_adj_1748.LUT_INIT = 16'hfffe;
    SB_CARRY add_224_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_279), 
            .CO(n40412));
    SB_LUT4 i1_4_lut_adj_1749 (.I0(n2427), .I1(n49053), .I2(n2422), .I3(n2425), 
            .O(n49055));
    defparam i1_4_lut_adj_1749.LUT_INIT = 16'hfffe;
    SB_LUT4 i22997_4_lut (.I0(n949), .I1(n2431), .I2(n2432), .I3(n2433), 
            .O(n36530));
    defparam i22997_4_lut.LUT_INIT = 16'hfcec;
    SB_DFFSR pwm_setpoint__i22 (.Q(pwm_setpoint[22]), .C(CLK_c), .D(pwm_setpoint_23__N_191[22]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i21 (.Q(pwm_setpoint[21]), .C(CLK_c), .D(pwm_setpoint_23__N_191[21]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i20 (.Q(pwm_setpoint[20]), .C(CLK_c), .D(pwm_setpoint_23__N_191[20]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i19 (.Q(pwm_setpoint[19]), .C(CLK_c), .D(pwm_setpoint_23__N_191[19]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i18 (.Q(pwm_setpoint[18]), .C(CLK_c), .D(pwm_setpoint_23__N_191[18]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i17 (.Q(pwm_setpoint[17]), .C(CLK_c), .D(pwm_setpoint_23__N_191[17]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i16 (.Q(pwm_setpoint[16]), .C(CLK_c), .D(pwm_setpoint_23__N_191[16]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i15 (.Q(pwm_setpoint[15]), .C(CLK_c), .D(pwm_setpoint_23__N_191[15]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i14 (.Q(pwm_setpoint[14]), .C(CLK_c), .D(pwm_setpoint_23__N_191[14]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i13 (.Q(pwm_setpoint[13]), .C(CLK_c), .D(pwm_setpoint_23__N_191[13]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i12 (.Q(pwm_setpoint[12]), .C(CLK_c), .D(pwm_setpoint_23__N_191[12]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i11 (.Q(pwm_setpoint[11]), .C(CLK_c), .D(pwm_setpoint_23__N_191[11]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i10 (.Q(pwm_setpoint[10]), .C(CLK_c), .D(pwm_setpoint_23__N_191[10]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i9 (.Q(pwm_setpoint[9]), .C(CLK_c), .D(pwm_setpoint_23__N_191[9]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i8 (.Q(pwm_setpoint[8]), .C(CLK_c), .D(pwm_setpoint_23__N_191[8]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i7 (.Q(pwm_setpoint[7]), .C(CLK_c), .D(pwm_setpoint_23__N_191[7]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i6 (.Q(pwm_setpoint[6]), .C(CLK_c), .D(pwm_setpoint_23__N_191[6]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i5 (.Q(pwm_setpoint[5]), .C(CLK_c), .D(pwm_setpoint_23__N_191[5]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i4 (.Q(pwm_setpoint[4]), .C(CLK_c), .D(pwm_setpoint_23__N_191[4]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i3 (.Q(pwm_setpoint[3]), .C(CLK_c), .D(pwm_setpoint_23__N_191[3]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i2 (.Q(pwm_setpoint[2]), .C(CLK_c), .D(pwm_setpoint_23__N_191[2]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i1 (.Q(pwm_setpoint[1]), .C(CLK_c), .D(pwm_setpoint_23__N_191[1]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 i1_4_lut_adj_1750 (.I0(n2419), .I1(n2420), .I2(n49055), .I3(n2421), 
            .O(n49061));
    defparam i1_4_lut_adj_1750.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1751 (.I0(n2429), .I1(n2430), .I2(GND_net), .I3(GND_net), 
            .O(n49269));
    defparam i1_2_lut_adj_1751.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n40418), .O(encoder1_position_scaled_23__N_75[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1752 (.I0(n2418), .I1(n49269), .I2(n49061), .I3(n36530), 
            .O(n49065));
    defparam i1_4_lut_adj_1752.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n49065), 
            .O(n49071));
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'hfffe;
    SB_LUT4 i37041_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52524));
    defparam i37041_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37336_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n49071), 
            .O(n2445));
    defparam i37336_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n41092));
    SB_LUT4 encoder0_position_31__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1515_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHC_184 (.Q(GHC), .C(CLK_c), .E(n29048), .D(GHC_N_403), 
            .R(n29375));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_mux_3_i11_3_lut (.I0(encoder0_position[10]), 
            .I1(n23), .I2(encoder0_position[31]), .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36347_3_lut (.I0(n2247), .I1(n2148), .I2(n2049), .I3(GND_net), 
            .O(n51830));
    defparam i36347_3_lut.LUT_INIT = 16'h7f7f;
    SB_LUT4 encoder0_position_31__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n40783), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n40693), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5147), .CO(n40694));
    SB_LUT4 add_145_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n40411), .O(n1077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1383_rep_71_3_lut (.I0(n2095), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n50243));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1383_rep_71_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1450_rep_67_3_lut (.I0(n50243), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n50239));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1450_rep_67_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1517_3_lut (.I0(n50239), .I1(n2028), 
            .I2(n51830), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i37301_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52784));
    defparam i37301_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n2326), .I1(n2324), .I2(n2327), .I3(n2325), 
            .O(n48853));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1755 (.I0(n2322), .I1(n2328), .I2(n2323), .I3(GND_net), 
            .O(n48855));
    defparam i1_3_lut_adj_1755.LUT_INIT = 16'hfefe;
    SB_LUT4 i22999_4_lut (.I0(n948), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n36532));
    defparam i22999_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1756 (.I0(n2320), .I1(n2321), .I2(n48855), .I3(n48853), 
            .O(n48861));
    defparam i1_4_lut_adj_1756.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1757 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n49043));
    defparam i1_2_lut_adj_1757.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n49043), .I1(n2319), .I2(n48861), .I3(n36532), 
            .O(n48865));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n48865), 
            .O(n48871));
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 i37305_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n48871), 
            .O(n2346));
    defparam i37305_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_238_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[9]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n40421), .O(encoder1_position_scaled_23__N_75[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16138_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n48426), .I3(GND_net), .O(n29660));   // verilog/coms.v(127[12] 300[6])
    defparam i16138_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5146), .I3(n40692), .O(displacement_23__N_99[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n40410), .O(n1078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_766_6 (.CI(n40783), .I0(n1130), 
            .I1(GND_net), .CO(n40784));
    SB_LUT4 encoder0_position_31__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5108));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHB_182 (.Q(GHB), .C(CLK_c), .E(n29048), .D(GHB_N_389), 
            .R(n29375));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36608_3_lut (.I0(n2028), .I1(n2095), .I2(n2049), .I3(GND_net), 
            .O(n2127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36608_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36609_3_lut (.I0(n2127), .I1(n2194), .I2(n2148), .I3(GND_net), 
            .O(n2226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36609_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_224_12 (.CI(n40421), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n40422));
    SB_LUT4 encoder0_position_31__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i12_3_lut (.I0(encoder0_position[11]), 
            .I1(n22), .I2(encoder0_position[31]), .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37269_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52752));
    defparam i37269_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(n2228), .I1(n2226), .I2(n2225), .I3(n2227), 
            .O(n49021));
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 i22880_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n36412));
    defparam i22880_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n2222), .I1(n49021), .I2(n2223), .I3(n2224), 
            .O(n49025));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n2229), .I1(n36412), .I2(n2230), .I3(n2231), 
            .O(n46756));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n2220), .I1(n46756), .I2(n2221), .I3(n49025), 
            .O(n49031));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n2217), .I1(n2218), .I2(n2219), .I3(n49031), 
            .O(n49037));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hfffe;
    SB_LUT4 i37273_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n49037), 
            .O(n2247));
    defparam i37273_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n40782), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_215), 
            .I3(n40457), .O(pwm_setpoint_23__N_191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n40420), .O(encoder1_position_scaled_23__N_75[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n40692), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5146), .CO(n40693));
    SB_LUT4 encoder0_position_31__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5145), .I3(n40691), .O(displacement_23__N_99[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n40691), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5145), .CO(n40692));
    SB_CARRY add_224_11 (.CI(n40420), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n40421));
    SB_LUT4 encoder0_position_31__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1382_rep_83_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1382_rep_83_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5144), .I3(n40690), .O(displacement_23__N_99[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n40690), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5144), .CO(n40691));
    SB_LUT4 encoder0_position_31__I_0_i1384_rep_77_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1384_rep_77_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1179_rep_97_3_lut (.I0(n1795), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n50269));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1179_rep_97_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36070_2_lut (.I0(n1851), .I1(n1752), .I2(GND_net), .I3(GND_net), 
            .O(n51552));
    defparam i36070_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 encoder0_position_31__I_0_i1246_rep_93_3_lut (.I0(n50269), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n50265));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1246_rep_93_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_766_5 (.CI(n40782), .I0(n1131), 
            .I1(VCC_net), .CO(n40783));
    SB_LUT4 i36606_4_lut (.I0(n50265), .I1(n1728), .I2(n1950), .I3(n51552), 
            .O(n52089));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36606_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5143), .I3(n40689), .O(displacement_23__N_99[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n40781), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_32 (.CI(n40410), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n40411));
    SB_CARRY add_224_9 (.CI(n40418), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n40419));
    SB_LUT4 i36607_3_lut (.I0(n52089), .I1(n2092), .I2(n2049), .I3(GND_net), 
            .O(n2124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36607_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_mux_3_i13_3_lut (.I0(encoder0_position[12]), 
            .I1(n21), .I2(encoder0_position[31]), .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n3), 
            .I3(n40456), .O(pwm_setpoint_23__N_191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_29_lut (.I0(n52972), .I1(n2907), 
            .I2(VCC_net), .I3(n41550), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n40689), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5143), .CO(n40690));
    SB_LUT4 encoder0_position_31__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n41549), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_24 (.CI(n40456), .I0(GND_net), .I1(n3), 
            .CO(n40457));
    SB_LUT4 add_145_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n40409), .O(n1079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_4 (.CI(n40781), .I0(n1132), 
            .I1(GND_net), .CO(n40782));
    SB_CARRY encoder0_position_31__I_0_add_1972_28 (.CI(n41549), .I0(n2908), 
            .I1(VCC_net), .CO(n41550));
    SB_LUT4 i37236_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52719));
    defparam i37236_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_224_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n40419), .O(encoder1_position_scaled_23__N_75[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1765 (.I0(n2125), .I1(n2124), .I2(n2128), .I3(GND_net), 
            .O(n48787));
    defparam i1_3_lut_adj_1765.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n40780), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1766 (.I0(n2123), .I1(n2127), .I2(n2126), .I3(GND_net), 
            .O(n48789));
    defparam i1_3_lut_adj_1766.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n41548), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5141), .I3(n40688), .O(displacement_23__N_99[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_27 (.CI(n41548), .I0(n2909), 
            .I1(VCC_net), .CO(n41549));
    SB_LUT4 encoder0_position_31__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n41547), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23003_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n36536));
    defparam i23003_4_lut.LUT_INIT = 16'hfcec;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_10_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n4_adj_5102), 
            .I3(n40455), .O(pwm_setpoint_23__N_191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n40688), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5141), .CO(n40689));
    SB_CARRY encoder0_position_31__I_0_add_1972_26 (.CI(n41547), .I0(n2910), 
            .I1(VCC_net), .CO(n41548));
    SB_LUT4 i1_4_lut_adj_1767 (.I0(n2121), .I1(n2122), .I2(n48789), .I3(n48787), 
            .O(n48795));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n41546), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_25 (.CI(n41546), .I0(n2911), 
            .I1(VCC_net), .CO(n41547));
    SB_LUT4 encoder0_position_31__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n41545), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(n2129), .I1(n48795), .I2(n36536), .I3(n2130), 
            .O(n48797));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'heccc;
    SB_CARRY encoder0_position_31__I_0_add_1972_24 (.CI(n41545), .I0(n2912), 
            .I1(VCC_net), .CO(n41546));
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n2118), .I1(n2119), .I2(n48797), .I3(n2120), 
            .O(n48803));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n41544), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_23 (.CI(n41544), .I0(n2913), 
            .I1(VCC_net), .CO(n41545));
    SB_LUT4 encoder0_position_31__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n41543), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37241_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n48803), 
            .O(n2148));
    defparam i37241_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_1972_22 (.CI(n41543), .I0(n2914), 
            .I1(VCC_net), .CO(n41544));
    SB_LUT4 encoder0_position_31__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n41542), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_21 (.CI(n41542), .I0(n2915), 
            .I1(VCC_net), .CO(n41543));
    SB_LUT4 encoder0_position_31__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n41541), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_20 (.CI(n41541), .I0(n2916), 
            .I1(VCC_net), .CO(n41542));
    SB_LUT4 encoder0_position_31__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n41540), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_19 (.CI(n41540), .I0(n2917), 
            .I1(VCC_net), .CO(n41541));
    SB_LUT4 i36519_3_lut (.I0(n1827), .I1(n1894), .I2(n1851), .I3(GND_net), 
            .O(n1926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n41539), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_18 (.CI(n41539), .I0(n2918), 
            .I1(VCC_net), .CO(n41540));
    SB_LUT4 i36483_3_lut (.I0(n1926), .I1(n1993), .I2(n1950), .I3(GND_net), 
            .O(n2025));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36483_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n41538), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_17 (.CI(n41538), .I0(n2919), 
            .I1(VCC_net), .CO(n41539));
    SB_CARRY encoder0_position_31__I_0_add_766_3 (.CI(n40780), .I0(n1133), 
            .I1(VCC_net), .CO(n40781));
    SB_LUT4 encoder0_position_31__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n41537), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36521_3_lut (.I0(n1826), .I1(n1893), .I2(n1851), .I3(GND_net), 
            .O(n1925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5140), .I3(n40687), .O(displacement_23__N_99[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_16 (.CI(n41537), .I0(n2920), 
            .I1(VCC_net), .CO(n41538));
    SB_LUT4 encoder0_position_31__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n41536), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n40687), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5140), .CO(n40688));
    SB_CARRY encoder0_position_31__I_0_add_1972_15 (.CI(n41536), .I0(n2921), 
            .I1(VCC_net), .CO(n41537));
    SB_LUT4 encoder0_position_31__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n41535), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_14 (.CI(n41535), .I0(n2922), 
            .I1(VCC_net), .CO(n41536));
    SB_LUT4 encoder0_position_31__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n41534), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_31 (.CI(n40409), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n40410));
    SB_CARRY encoder0_position_31__I_0_add_1972_13 (.CI(n41534), .I0(n2923), 
            .I1(VCC_net), .CO(n41535));
    SB_LUT4 encoder0_position_31__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n41533), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_12 (.CI(n41533), .I0(n2924), 
            .I1(VCC_net), .CO(n41534));
    SB_LUT4 encoder0_position_31__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n41532), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_11 (.CI(n41532), .I0(n2925), 
            .I1(VCC_net), .CO(n41533));
    SB_CARRY unary_minus_10_add_3_23 (.CI(n40455), .I0(GND_net), .I1(n4_adj_5102), 
            .CO(n40456));
    SB_LUT4 encoder0_position_31__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n41531), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5139), .I3(n40686), .O(displacement_23__N_99[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_10 (.CI(n41531), .I0(n2926), 
            .I1(VCC_net), .CO(n41532));
    SB_LUT4 encoder0_position_31__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i771_3_lut (.I0(n1128), .I1(n1195_adj_5182), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i777_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22713_3_lut (.I0(n937), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n36240));
    defparam i22713_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1770 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n48915));
    defparam i1_3_lut_adj_1770.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(n1229), .I1(n36240), .I2(n1230), .I3(n1231), 
            .O(n46666));
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'ha080;
    SB_LUT4 i36481_3_lut (.I0(n1925), .I1(n1992), .I2(n1950), .I3(GND_net), 
            .O(n2024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36481_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n41530), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_9 (.CI(n41530), .I0(n2927), 
            .I1(VCC_net), .CO(n41531));
    SB_LUT4 encoder0_position_31__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n41529), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1316_rep_89_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1316_rep_89_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_8 (.CI(n41529), .I0(n2928), 
            .I1(VCC_net), .CO(n41530));
    SB_LUT4 encoder0_position_31__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n41528), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_7 (.CI(n41528), .I0(n2929), 
            .I1(GND_net), .CO(n41529));
    SB_LUT4 encoder0_position_31__I_0_add_766_2_lut (.I0(GND_net), .I1(n936), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n41527), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_2 (.CI(VCC_net), .I0(n936), 
            .I1(GND_net), .CO(n40780));
    SB_LUT4 add_145_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n40390), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_6 (.CI(n41527), .I0(n2930), 
            .I1(GND_net), .CO(n41528));
    SB_LUT4 encoder0_position_31__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n41526), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_5 (.CI(n41526), .I0(n2931), 
            .I1(VCC_net), .CO(n41527));
    SB_LUT4 encoder0_position_31__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n41525), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_4 (.CI(n41525), .I0(n2932), 
            .I1(GND_net), .CO(n41526));
    SB_LUT4 encoder0_position_31__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n41524), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_3 (.CI(n41524), .I0(n2933), 
            .I1(VCC_net), .CO(n41525));
    SB_LUT4 encoder0_position_31__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n41524));
    SB_LUT4 i36602_3_lut (.I0(n1828), .I1(n1895), .I2(n1851), .I3(GND_net), 
            .O(n1927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36602_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36603_3_lut (.I0(n1927), .I1(n1994), .I2(n1950), .I3(GND_net), 
            .O(n2026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36603_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5107));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n40686), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5139), .CO(n40687));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5138), .I3(n40685), .O(displacement_23__N_99[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n40685), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5138), .CO(n40686));
    SB_LUT4 encoder0_position_31__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i14_3_lut (.I0(encoder0_position[13]), 
            .I1(n20), .I2(encoder0_position[31]), .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37206_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52689));
    defparam i37206_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22717_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n36244));
    defparam i22717_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1772 (.I0(n2026), .I1(n2027), .I2(GND_net), .I3(GND_net), 
            .O(n48989));
    defparam i1_2_lut_adj_1772.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n2028), .I1(n48989), .I2(n2024), .I3(n2025), 
            .O(n48993));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n2029), .I1(n36244), .I2(n2030), .I3(n2031), 
            .O(n46749));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n48993), 
            .O(n48999));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5137), .I3(n40684), .O(displacement_23__N_99[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n2019), .I1(n2020), .I2(n48999), .I3(n46749), 
            .O(n49005));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'hfffe;
    SB_LUT4 i37210_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n49005), 
            .O(n2049));
    defparam i37210_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_10_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5106));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n40684), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5137), .CO(n40685));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5136), .I3(n40683), .O(displacement_23__N_99[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_16_lut (.I0(n52590), .I1(n1620), 
            .I2(VCC_net), .I3(n41081), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n41080), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_15 (.CI(n41080), .I0(n1621), 
            .I1(VCC_net), .CO(n41081));
    SB_LUT4 encoder0_position_31__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n41079), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_14 (.CI(n41079), .I0(n1622), 
            .I1(VCC_net), .CO(n41080));
    SB_LUT4 i16139_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n48426), .I3(GND_net), .O(n29661));   // verilog/coms.v(127[12] 300[6])
    defparam i16139_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHA_180 (.Q(GHA), .C(CLK_c), .E(n29048), .D(GHA_N_367), 
            .R(n29375));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n41078), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_13 (.CI(n41078), .I0(n1623), 
            .I1(VCC_net), .CO(n41079));
    SB_LUT4 encoder0_position_31__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1241_3_lut (.I0(n1822), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1243_3_lut (.I0(n1824), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n40683), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5136), .CO(n40684));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5135), .I3(n40682), .O(displacement_23__N_99[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n41077), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_12 (.CI(n41077), .I0(n1624), 
            .I1(VCC_net), .CO(n41078));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i15_3_lut (.I0(encoder0_position[14]), 
            .I1(n19), .I2(encoder0_position[31]), .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n41076), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n5), 
            .I3(n40454), .O(pwm_setpoint_23__N_191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_11 (.CI(n41076), .I0(n1625), 
            .I1(VCC_net), .CO(n41077));
    SB_LUT4 i37182_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52665));
    defparam i37182_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n40769), .O(n1093_adj_5173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_10 (.CI(n40419), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n40420));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n40682), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5135), .CO(n40683));
    SB_LUT4 encoder0_position_31__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n41075), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_10 (.CI(n41075), .I0(n1626), 
            .I1(VCC_net), .CO(n41076));
    SB_LUT4 encoder0_position_31__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n41074), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n40768), .O(n1094_adj_5174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n1927), .I1(n1926), .I2(n1925), .I3(n1928), 
            .O(n48765));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_LUT4 i22719_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n36246));
    defparam i22719_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_31__I_0_add_699_9 (.CI(n40768), .I0(n1027), 
            .I1(VCC_net), .CO(n40769));
    SB_LUT4 i1_4_lut_adj_1778 (.I0(n1922), .I1(n1923), .I2(n48765), .I3(n1924), 
            .O(n48771));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n1929), .I1(n36246), .I2(n1930), .I3(n1931), 
            .O(n46713));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1780 (.I0(n1920), .I1(n46713), .I2(n1921), .I3(n48771), 
            .O(n48777));
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 i37185_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n48777), 
            .O(n1950));
    defparam i37185_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i37158_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52641));
    defparam i37158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1781 (.I0(n1825), .I1(n1827), .I2(n1826), .I3(n1828), 
            .O(n48965));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'hfffe;
    SB_LUT4 i22723_3_lut (.I0(n943), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n36250));
    defparam i22723_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1782 (.I0(n1823), .I1(n1824), .I2(n48965), .I3(GND_net), 
            .O(n48969));
    defparam i1_3_lut_adj_1782.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1783 (.I0(n1829), .I1(n36250), .I2(n1830), .I3(n1831), 
            .O(n46728));
    defparam i1_4_lut_adj_1783.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1784 (.I0(n1821), .I1(n1822), .I2(n46728), .I3(n48969), 
            .O(n48975));
    defparam i1_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n40767), .O(n1095_adj_5175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37161_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n48975), 
            .O(n1851));
    defparam i37161_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_1101_9 (.CI(n41074), .I0(n1627), 
            .I1(VCC_net), .CO(n41075));
    SB_LUT4 i16140_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n48426), .I3(GND_net), .O(n29662));   // verilog/coms.v(127[12] 300[6])
    defparam i16140_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_699_8 (.CI(n40767), .I0(n1028), 
            .I1(VCC_net), .CO(n40768));
    SB_LUT4 i37132_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52615));
    defparam i37132_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n41073), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_8 (.CI(n41073), .I0(n1628), 
            .I1(VCC_net), .CO(n41074));
    SB_LUT4 i37107_1_lut (.I0(n1653_adj_5183), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n52590));
    defparam i37107_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37088_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52571));
    defparam i37088_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5134), .I3(n40681), .O(displacement_23__N_99[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n41072), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_7 (.CI(n41072), .I0(n1629), 
            .I1(GND_net), .CO(n41073));
    SB_LUT4 i37040_4_lut (.I0(n1225), .I1(n1224), .I2(n46666), .I3(n48915), 
            .O(n1257));
    defparam i37040_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(244[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37070_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52553));
    defparam i37070_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(CLK_c), .D(displacement_23__N_99[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i37037_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52520));
    defparam i37037_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37022_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52505));
    defparam i37022_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(CLK_c), .D(displacement_23__N_99[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n41071), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n40766), .O(n1096_adj_5176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_6 (.CI(n41071), .I0(n1630), 
            .I1(GND_net), .CO(n41072));
    SB_CARRY unary_minus_10_add_3_22 (.CI(n40454), .I0(GND_net), .I1(n5), 
            .CO(n40455));
    SB_LUT4 add_145_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n40408), .O(n1080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_7 (.CI(n40766), .I0(n1029), 
            .I1(GND_net), .CO(n40767));
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(CLK_c), .D(displacement_23__N_99[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(CLK_c), .D(displacement_23__N_99[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(CLK_c), .D(displacement_23__N_99[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(CLK_c), .D(displacement_23__N_99[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(CLK_c), .D(displacement_23__N_99[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(CLK_c), .D(displacement_23__N_99[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(CLK_c), .D(displacement_23__N_99[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(CLK_c), .D(displacement_23__N_99[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(CLK_c), .D(displacement_23__N_99[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(CLK_c), .D(displacement_23__N_99[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(CLK_c), .D(displacement_23__N_99[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(CLK_c), .D(displacement_23__N_99[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(CLK_c), .D(displacement_23__N_99[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(CLK_c), .D(displacement_23__N_99[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(CLK_c), .D(displacement_23__N_99[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(CLK_c), .D(displacement_23__N_99[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(CLK_c), .D(displacement_23__N_99[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(CLK_c), .D(displacement_23__N_99[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(CLK_c), .D(displacement_23__N_99[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(CLK_c), .D(displacement_23__N_99[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(CLK_c), .D(displacement_23__N_99[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i37008_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52491));
    defparam i37008_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5194));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i22_3_lut (.I0(encoder0_position[21]), 
            .I1(n12_adj_5151), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n937));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n41070), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n6), 
            .I3(n40453), .O(pwm_setpoint_23__N_191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i16_3_lut (.I0(encoder0_position[15]), 
            .I1(n18), .I2(encoder0_position[31]), .I3(GND_net), .O(n943));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[10]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_145_12 (.CI(n40390), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n40391));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n40681), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5134), .CO(n40682));
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_CARRY encoder0_position_31__I_0_add_1101_5 (.CI(n41070), .I0(n1631), 
            .I1(VCC_net), .CO(n41071));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5133), .I3(n40680), .O(displacement_23__N_99[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF dti_counter_2056__i0 (.Q(dti_counter[0]), .C(CLK_c), .D(n55));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_LUT4 encoder0_position_31__I_0_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n40765), .O(n1097_adj_5177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n40389), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n40680), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5133), .CO(n40681));
    SB_LUT4 encoder0_position_31__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n41069), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_238_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[11]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_1101_4 (.CI(n41069), .I0(n1632), 
            .I1(GND_net), .CO(n41070));
    SB_LUT4 encoder0_position_31__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n41068), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_3 (.CI(n41068), .I0(n1633), 
            .I1(VCC_net), .CO(n41069));
    SB_CARRY encoder0_position_31__I_0_add_699_6 (.CI(n40765), .I0(n1030), 
            .I1(GND_net), .CO(n40766));
    SB_CARRY add_145_30 (.CI(n40408), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n40409));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5132), .I3(n40679), .O(displacement_23__N_99[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_21 (.CI(n40453), .I0(GND_net), .I1(n6), 
            .CO(n40454));
    SB_LUT4 encoder0_position_31__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n40764), .O(n1098_adj_5178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n40407), .O(n1081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n41068));
    SB_LUT4 encoder0_position_31__I_0_add_1034_15_lut (.I0(n52571), .I1(n1521), 
            .I2(VCC_net), .I3(n41067), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n41066), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_14 (.CI(n41066), .I0(n1522), 
            .I1(VCC_net), .CO(n41067));
    SB_CARRY encoder0_position_31__I_0_add_699_5 (.CI(n40764), .I0(n1031), 
            .I1(VCC_net), .CO(n40765));
    SB_LUT4 encoder0_position_31__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n41065), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22787_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n36316));
    defparam i22787_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_CARRY encoder0_position_31__I_0_add_1034_13 (.CI(n41065), .I0(n1523), 
            .I1(VCC_net), .CO(n41066));
    SB_LUT4 encoder0_position_31__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n41064), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_12 (.CI(n41064), .I0(n1524), 
            .I1(VCC_net), .CO(n41065));
    SB_LUT4 encoder0_position_31__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n41063), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_11 (.CI(n41063), .I0(n1525), 
            .I1(VCC_net), .CO(n41064));
    SB_LUT4 encoder0_position_31__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n41062), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_10 (.CI(n41062), .I0(n1526), 
            .I1(VCC_net), .CO(n41063));
    SB_LUT4 encoder0_position_31__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n41061), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_9 (.CI(n41061), .I0(n1527), 
            .I1(VCC_net), .CO(n41062));
    SB_LUT4 encoder0_position_31__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n41060), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_8 (.CI(n41060), .I0(n1528), 
            .I1(VCC_net), .CO(n41061));
    SB_LUT4 encoder0_position_31__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n41059), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n7), 
            .I3(n40452), .O(pwm_setpoint_23__N_191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n40679), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5132), .CO(n40680));
    SB_CARRY encoder0_position_31__I_0_add_1034_7 (.CI(n41059), .I0(n1529), 
            .I1(GND_net), .CO(n41060));
    SB_LUT4 add_145_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n40383), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5105));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_145_29 (.CI(n40407), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n40408));
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(CLK_c), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(CLK_c), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_mux_3_i26_3_lut (.I0(encoder0_position[25]), 
            .I1(n8_adj_5161), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n834));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n41058), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31070_3_lut (.I0(n7_adj_5162), .I1(n7287), .I2(n46394), .I3(GND_net), 
            .O(n46432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n48661));
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'hfffe;
    SB_LUT4 i31071_3_lut (.I0(encoder0_position[26]), .I1(n46432), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n40763), .O(n1099_adj_5179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_4 (.CI(n40763), .I0(n1032), 
            .I1(GND_net), .CO(n40764));
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n1329), .I1(n36316), .I2(n1330), .I3(n1331), 
            .O(n46663));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n40762), .O(n1100_adj_5180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31072_3_lut (.I0(n6_adj_5163), .I1(n7286), .I2(n46394), .I3(GND_net), 
            .O(n46434));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31073_3_lut (.I0(encoder0_position[27]), .I1(n46434), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1034_6 (.CI(n41058), .I0(n1530), 
            .I1(GND_net), .CO(n41059));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5131), .I3(n40678), .O(displacement_23__N_99[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_20 (.CI(n40452), .I0(GND_net), .I1(n7), 
            .CO(n40453));
    SB_LUT4 encoder0_position_31__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n41057), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_3 (.CI(n40762), .I0(n1033), 
            .I1(VCC_net), .CO(n40763));
    SB_LUT4 unary_minus_10_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n8_adj_5103), 
            .I3(n40451), .O(pwm_setpoint_23__N_191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n40678), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5131), .CO(n40679));
    SB_LUT4 encoder0_position_31__I_0_add_699_2_lut (.I0(GND_net), .I1(n935), 
            .I2(GND_net), .I3(VCC_net), .O(n1101_adj_5181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5130), .I3(n40677), .O(displacement_23__N_99[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_5 (.CI(n41057), .I0(n1531), 
            .I1(VCC_net), .CO(n41058));
    SB_CARRY encoder0_position_31__I_0_add_699_2 (.CI(VCC_net), .I0(n935), 
            .I1(GND_net), .CO(n40762));
    SB_CARRY add_145_5 (.CI(n40383), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n40384));
    SB_LUT4 encoder0_position_31__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n41056), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_19 (.CI(n40451), .I0(GND_net), .I1(n8_adj_5103), 
            .CO(n40452));
    SB_LUT4 encoder0_position_31__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n40761), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n40760), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_11 (.CI(n40389), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n40390));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n40677), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5130), .CO(n40678));
    SB_CARRY encoder0_position_31__I_0_add_632_8 (.CI(n40760), .I0(n928), 
            .I1(VCC_net), .CO(n40761));
    SB_CARRY encoder0_position_31__I_0_add_1034_4 (.CI(n41056), .I0(n1532), 
            .I1(GND_net), .CO(n41057));
    SB_LUT4 encoder0_position_31__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n40759), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n40388), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5129), .I3(n40676), .O(displacement_23__N_99[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_7 (.CI(n40759), .I0(n929), 
            .I1(GND_net), .CO(n40760));
    SB_LUT4 encoder0_position_31__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n41055), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_3 (.CI(n41055), .I0(n1533), 
            .I1(VCC_net), .CO(n41056));
    SB_LUT4 add_145_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n40406), .O(n1082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n40758), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_145_28 (.CI(n40406), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n40407));
    SB_CARRY encoder0_position_31__I_0_add_632_6 (.CI(n40758), .I0(n930), 
            .I1(GND_net), .CO(n40759));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n40676), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5129), .CO(n40677));
    SB_CARRY encoder0_position_31__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n41055));
    SB_LUT4 encoder0_position_31__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n40757), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5128), .I3(n40675), .O(displacement_23__N_99[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n40675), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5128), .CO(n40676));
    SB_CARRY encoder0_position_31__I_0_add_632_5 (.CI(n40757), .I0(n931), 
            .I1(VCC_net), .CO(n40758));
    SB_LUT4 unary_minus_10_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n9), 
            .I3(n40450), .O(pwm_setpoint_23__N_191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5127), .I3(n40674), .O(displacement_23__N_99[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n40405), .O(n1083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n40756), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n40674), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5127), .CO(n40675));
    SB_CARRY unary_minus_10_add_3_18 (.CI(n40450), .I0(GND_net), .I1(n9), 
            .CO(n40451));
    SB_LUT4 unary_minus_10_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n10_adj_5104), 
            .I3(n40449), .O(pwm_setpoint_23__N_191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_27 (.CI(n40405), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n40406));
    SB_LUT4 add_145_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n40404), .O(n1084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_4 (.CI(n40756), .I0(n932), 
            .I1(GND_net), .CO(n40757));
    SB_CARRY add_145_26 (.CI(n40404), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n40405));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5126), .I3(n40673), .O(displacement_23__N_99[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n40403), .O(n1085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n40673), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5126), .CO(n40674));
    SB_CARRY add_145_25 (.CI(n40403), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n40404));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5125), .I3(VCC_net), .O(displacement_23__N_99[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5125), .CO(n40673));
    SB_LUT4 encoder0_position_31__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n40755), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_632_3 (.CI(n40755), .I0(n933), 
            .I1(VCC_net), .CO(n40756));
    SB_CARRY unary_minus_10_add_3_17 (.CI(n40449), .I0(GND_net), .I1(n10_adj_5104), 
            .CO(n40450));
    SB_LUT4 i16073_4_lut (.I0(state_7__N_4103[3]), .I1(data[7]), .I2(n35513), 
            .I3(n27954), .O(n29595));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16073_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16074_4_lut (.I0(state_7__N_4103[3]), .I1(data[6]), .I2(n35513), 
            .I3(n27911), .O(n29596));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16074_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16075_4_lut (.I0(state_7__N_4103[3]), .I1(data[5]), .I2(n4_adj_5097), 
            .I3(n27954), .O(n29597));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16075_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16076_4_lut (.I0(state_7__N_4103[3]), .I1(data[4]), .I2(n4_adj_5097), 
            .I3(n27911), .O(n29598));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16076_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_967_14_lut (.I0(n52553), .I1(n1422), 
            .I2(VCC_net), .I3(n41054), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_145_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n40402), .O(n1086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_28_lut (.I0(n52940), .I1(n2808), 
            .I2(VCC_net), .I3(n41428), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n41427), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_27 (.CI(n41427), .I0(n2809), 
            .I1(VCC_net), .CO(n41428));
    SB_LUT4 encoder0_position_31__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n41426), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_26 (.CI(n41426), .I0(n2810), 
            .I1(VCC_net), .CO(n41427));
    SB_LUT4 i1_3_lut_adj_1787 (.I0(n5_adj_5123), .I1(n3_adj_5166), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n48985));
    defparam i1_3_lut_adj_1787.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_31__I_0_i500_4_lut (.I0(n2_adj_5167), .I1(n7282), 
            .I2(n48985), .I3(encoder0_position[31]), .O(n828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 encoder0_position_31__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n41425), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_25 (.CI(n41425), .I0(n2811), 
            .I1(VCC_net), .CO(n41426));
    SB_LUT4 encoder0_position_31__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n41424), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_10 (.CI(n40388), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n40389));
    SB_LUT4 encoder0_position_31__I_0_add_632_2_lut (.I0(GND_net), .I1(n934), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_24 (.CI(n41424), .I0(n2812), 
            .I1(VCC_net), .CO(n41425));
    SB_CARRY encoder0_position_31__I_0_add_632_2 (.CI(VCC_net), .I0(n934), 
            .I1(GND_net), .CO(n40755));
    SB_LUT4 encoder0_position_31__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n41423), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_23 (.CI(n41423), .I0(n2813), 
            .I1(VCC_net), .CO(n41424));
    SB_LUT4 encoder0_position_31__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n41422), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_22 (.CI(n41422), .I0(n2814), 
            .I1(VCC_net), .CO(n41423));
    SB_LUT4 encoder0_position_31__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n41421), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n40754), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n41053), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_21 (.CI(n41421), .I0(n2815), 
            .I1(VCC_net), .CO(n41422));
    SB_LUT4 encoder0_position_31__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n41420), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_20 (.CI(n41420), .I0(n2816), 
            .I1(VCC_net), .CO(n41421));
    SB_LUT4 encoder0_position_31__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n41419), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_19 (.CI(n41419), .I0(n2817), 
            .I1(VCC_net), .CO(n41420));
    SB_LUT4 encoder0_position_31__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n41418), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n40753), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_18 (.CI(n41418), .I0(n2818), 
            .I1(VCC_net), .CO(n41419));
    SB_LUT4 encoder0_position_31__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n41417), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_17 (.CI(n41417), .I0(n2819), 
            .I1(VCC_net), .CO(n41418));
    SB_LUT4 encoder0_position_31__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n41416), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_16 (.CI(n41416), .I0(n2820), 
            .I1(VCC_net), .CO(n41417));
    SB_LUT4 encoder0_position_31__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n41415), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_15 (.CI(n41415), .I0(n2821), 
            .I1(VCC_net), .CO(n41416));
    SB_LUT4 encoder0_position_31__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n41414), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_14 (.CI(n41414), .I0(n2822), 
            .I1(VCC_net), .CO(n41415));
    SB_LUT4 encoder0_position_31__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n41413), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_13 (.CI(n41413), .I0(n2823), 
            .I1(VCC_net), .CO(n41414));
    SB_LUT4 encoder0_position_31__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n41412), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_12 (.CI(n41412), .I0(n2824), 
            .I1(VCC_net), .CO(n41413));
    SB_LUT4 encoder0_position_31__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n41411), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_11 (.CI(n41411), .I0(n2825), 
            .I1(VCC_net), .CO(n41412));
    SB_LUT4 encoder0_position_31__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n41410), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_10 (.CI(n41410), .I0(n2826), 
            .I1(VCC_net), .CO(n41411));
    SB_LUT4 encoder0_position_31__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n41409), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_9 (.CI(n41409), .I0(n2827), 
            .I1(VCC_net), .CO(n41410));
    SB_LUT4 encoder0_position_31__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n41408), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_8 (.CI(n41408), .I0(n2828), 
            .I1(VCC_net), .CO(n41409));
    SB_LUT4 encoder0_position_31__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n41407), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_7 (.CI(n41407), .I0(n2829), 
            .I1(GND_net), .CO(n41408));
    SB_LUT4 encoder0_position_31__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n41406), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_6 (.CI(n41406), .I0(n2830), 
            .I1(GND_net), .CO(n41407));
    SB_LUT4 encoder0_position_31__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n41405), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37056_4_lut (.I0(n46663), .I1(n1323), .I2(n1324), .I3(n48661), 
            .O(n1356));
    defparam i37056_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_1905_5 (.CI(n41405), .I0(n2831), 
            .I1(VCC_net), .CO(n41406));
    SB_LUT4 encoder0_position_31__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n41404), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_4 (.CI(n41404), .I0(n2832), 
            .I1(GND_net), .CO(n41405));
    SB_LUT4 encoder0_position_31__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n41403), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i573_3_lut (.I0(n834), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_3 (.CI(n41403), .I0(n2833), 
            .I1(VCC_net), .CO(n41404));
    SB_LUT4 encoder0_position_31__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n41403));
    SB_LUT4 encoder0_position_31__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i25_3_lut (.I0(encoder0_position[24]), 
            .I1(n9_adj_5158), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n934));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_967_13 (.CI(n41053), .I0(n1423), 
            .I1(VCC_net), .CO(n41054));
    SB_CARRY encoder0_position_31__I_0_add_565_7 (.CI(n40753), .I0(n829), 
            .I1(GND_net), .CO(n40754));
    SB_LUT4 unary_minus_10_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11), 
            .I3(n40448), .O(pwm_setpoint_23__N_191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_16 (.CI(n40448), .I0(GND_net), .I1(n11), 
            .CO(n40449));
    SB_LUT4 encoder0_position_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n40752), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12), 
            .I3(n40447), .O(pwm_setpoint_23__N_191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_6 (.CI(n40752), .I0(n830), 
            .I1(GND_net), .CO(n40753));
    SB_CARRY add_145_24 (.CI(n40402), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n40403));
    SB_LUT4 add_145_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n40401), .O(n1087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n40751), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n41052), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_5 (.CI(n40751), .I0(n831), 
            .I1(VCC_net), .CO(n40752));
    SB_CARRY encoder0_position_31__I_0_add_967_12 (.CI(n41052), .I0(n1424), 
            .I1(VCC_net), .CO(n41053));
    SB_LUT4 encoder0_position_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n40750), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n41051), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_4 (.CI(n40750), .I0(n832), 
            .I1(GND_net), .CO(n40751));
    SB_LUT4 encoder0_position_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n40749), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5125));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_565_3 (.CI(n40749), .I0(n833), 
            .I1(VCC_net), .CO(n40750));
    SB_LUT4 encoder0_position_31__I_0_add_565_2_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_2 (.CI(VCC_net), .I0(n834), 
            .I1(GND_net), .CO(n40749));
    SB_CARRY encoder0_position_31__I_0_add_967_11 (.CI(n41051), .I0(n1425), 
            .I1(VCC_net), .CO(n41052));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5126));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_10_add_3_15 (.CI(n40447), .I0(GND_net), .I1(n12), 
            .CO(n40448));
    SB_LUT4 unary_minus_10_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n13_adj_5105), 
            .I3(n40446), .O(pwm_setpoint_23__N_191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n41050), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_10 (.CI(n41050), .I0(n1426), 
            .I1(VCC_net), .CO(n41051));
    SB_LUT4 encoder0_position_31__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_23 (.CI(n40401), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n40402));
    SB_LUT4 unary_minus_10_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5104));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16141_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n48426), .I3(GND_net), .O(n29663));   // verilog/coms.v(127[12] 300[6])
    defparam i16141_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[12]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_145_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n40400), .O(n1088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n41049), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n40382), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n40387), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_9 (.CI(n41049), .I0(n1427), 
            .I1(VCC_net), .CO(n41050));
    SB_LUT4 i16142_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n48426), .I3(GND_net), .O(n29664));   // verilog/coms.v(127[12] 300[6])
    defparam i16142_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1180_rep_100_3_lut (.I0(n1729), .I1(n1796), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1180_rep_100_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5127));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i21_3_lut (.I0(encoder0_position[20]), 
            .I1(n13), .I2(encoder0_position[31]), .I3(GND_net), .O(n938));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16143_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n48426), .I3(GND_net), .O(n29665));   // verilog/coms.v(127[12] 300[6])
    defparam i16143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16144_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n48426), .I3(GND_net), .O(n29666));   // verilog/coms.v(127[12] 300[6])
    defparam i16144_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n41048), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5128));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16145_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n48426), .I3(GND_net), .O(n29667));   // verilog/coms.v(127[12] 300[6])
    defparam i16145_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_8 (.CI(n41048), .I0(n1428), 
            .I1(VCC_net), .CO(n41049));
    SB_LUT4 encoder0_position_31__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n41047), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_14 (.CI(n40446), .I0(GND_net), .I1(n13_adj_5105), 
            .CO(n40447));
    SB_LUT4 unary_minus_10_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5106), 
            .I3(n40445), .O(pwm_setpoint_23__N_191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_7 (.CI(n41047), .I0(n1429), 
            .I1(GND_net), .CO(n41048));
    SB_CARRY add_145_22 (.CI(n40400), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n40401));
    SB_LUT4 i16146_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n48426), .I3(GND_net), .O(n29668));   // verilog/coms.v(127[12] 300[6])
    defparam i16146_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21913_2_lut (.I0(n25316), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n35426));
    defparam i21913_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_238_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[18]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16147_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n48426), .I3(GND_net), .O(n29669));   // verilog/coms.v(127[12] 300[6])
    defparam i16147_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5129));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[19]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY unary_minus_10_add_3_13 (.CI(n40445), .I0(GND_net), .I1(n14_adj_5106), 
            .CO(n40446));
    SB_LUT4 unary_minus_10_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5107), 
            .I3(n40444), .O(pwm_setpoint_23__N_191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n40399), .O(n1089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1178_3_lut (.I0(n1727), .I1(n1794), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1176_3_lut (.I0(n1725), .I1(n1792), 
            .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1174_3_lut (.I0(n1723), .I1(n1790), 
            .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_9 (.CI(n40387), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n40388));
    SB_LUT4 encoder0_position_31__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16148_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n48426), .I3(GND_net), .O(n29670));   // verilog/coms.v(127[12] 300[6])
    defparam i16148_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n41046), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_12 (.CI(n40444), .I0(GND_net), .I1(n15_adj_5107), 
            .CO(n40445));
    SB_CARRY encoder0_position_31__I_0_add_967_6 (.CI(n41046), .I0(n1430), 
            .I1(GND_net), .CO(n41047));
    SB_CARRY add_145_21 (.CI(n40399), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n40400));
    SB_LUT4 encoder0_position_31__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n41045), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_238_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[20]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_967_5 (.CI(n41045), .I0(n1431), 
            .I1(VCC_net), .CO(n41046));
    SB_LUT4 encoder0_position_31__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n41044), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_4 (.CI(n41044), .I0(n1432), 
            .I1(GND_net), .CO(n41045));
    SB_LUT4 encoder0_position_31__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n41043), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6643_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_403));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6643_3_lut_4_lut.LUT_INIT = 16'haa1c;
    SB_LUT4 i6645_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_412));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6645_3_lut_4_lut.LUT_INIT = 16'h1caa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5130));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5103));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5131));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5108), 
            .I3(n40443), .O(pwm_setpoint_23__N_191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_3 (.CI(n41043), .I0(n1433), 
            .I1(VCC_net), .CO(n41044));
    SB_LUT4 mux_238_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[21]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_145_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n40386), .O(n1102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i20_3_lut (.I0(encoder0_position[19]), 
            .I1(n14_adj_5099), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n939));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6639_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHB_N_389));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6639_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_CARRY unary_minus_10_add_3_11 (.CI(n40443), .I0(GND_net), .I1(n16_adj_5108), 
            .CO(n40444));
    SB_LUT4 mux_238_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[22]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i6641_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLB_N_398));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6641_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 mux_238_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[23]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n41043));
    SB_LUT4 encoder0_position_31__I_0_add_900_13_lut (.I0(n52524), .I1(n1323), 
            .I2(VCC_net), .I3(n41042), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_10_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5109), 
            .I3(n40442), .O(pwm_setpoint_23__N_191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n41041), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_12 (.CI(n41041), .I0(n1324), 
            .I1(VCC_net), .CO(n41042));
    SB_LUT4 encoder0_position_31__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n41040), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_11 (.CI(n41040), .I0(n1325), 
            .I1(VCC_net), .CO(n41041));
    SB_LUT4 add_145_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n40398), .O(n1090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n41039), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_10 (.CI(n40442), .I0(GND_net), .I1(n17_adj_5109), 
            .CO(n40443));
    SB_CARRY encoder0_position_31__I_0_add_900_10 (.CI(n41039), .I0(n1326), 
            .I1(VCC_net), .CO(n41040));
    SB_LUT4 encoder0_position_31__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n41038), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_9 (.CI(n41038), .I0(n1327), 
            .I1(VCC_net), .CO(n41039));
    SB_LUT4 encoder0_position_31__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n41037), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5117));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5110), 
            .I3(n40441), .O(pwm_setpoint_23__N_191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22772_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n36300));
    defparam i22772_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1788 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n48925));
    defparam i1_2_lut_adj_1788.LUT_INIT = 16'heeee;
    SB_LUT4 unary_minus_10_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_5116));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_900_8 (.CI(n41037), .I0(n1328), 
            .I1(VCC_net), .CO(n41038));
    SB_CARRY add_145_20 (.CI(n40398), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n40399));
    SB_LUT4 encoder0_position_31__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n41036), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_27_lut (.I0(n52908), .I1(n2709), 
            .I2(VCC_net), .I3(n41321), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_900_7 (.CI(n41036), .I0(n1329), 
            .I1(GND_net), .CO(n41037));
    SB_LUT4 encoder0_position_31__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n41035), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n41320), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_26 (.CI(n41320), .I0(n2710), 
            .I1(VCC_net), .CO(n41321));
    SB_CARRY encoder0_position_31__I_0_add_900_6 (.CI(n41035), .I0(n1330), 
            .I1(GND_net), .CO(n41036));
    SB_LUT4 encoder0_position_31__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n41319), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1838_25 (.CI(n41319), .I0(n2711), 
            .I1(VCC_net), .CO(n41320));
    SB_LUT4 encoder0_position_31__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n41318), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_10_add_3_9 (.CI(n40441), .I0(GND_net), .I1(n18_adj_5110), 
            .CO(n40442));
    SB_LUT4 encoder0_position_31__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n41034), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_24 (.CI(n41318), .I0(n2712), 
            .I1(VCC_net), .CO(n41319));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5111), 
            .I3(n40440), .O(pwm_setpoint_23__N_191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5115));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5214));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5213));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5212));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n1429), .I1(n36300), .I2(n1430), .I3(n1431), 
            .O(n46682));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_900_5 (.CI(n41034), .I0(n1331), 
            .I1(VCC_net), .CO(n41035));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5211));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5210));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5209));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5208));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n41317), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_23 (.CI(n41317), .I0(n2713), 
            .I1(VCC_net), .CO(n41318));
    SB_LUT4 encoder0_position_31__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n41033), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5207));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n41316), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5206));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1838_22 (.CI(n41316), .I0(n2714), 
            .I1(VCC_net), .CO(n41317));
    SB_CARRY encoder0_position_31__I_0_add_900_4 (.CI(n41033), .I0(n1332), 
            .I1(GND_net), .CO(n41034));
    SB_LUT4 encoder0_position_31__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n41315), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_21 (.CI(n41315), .I0(n2715), 
            .I1(VCC_net), .CO(n41316));
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n48925), 
            .O(n48931));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n41314), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(CLK_c), 
            .E(n6_adj_5189), .D(commutation_state_7__N_216[0]), .S(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1838_20 (.CI(n41314), .I0(n2716), 
            .I1(VCC_net), .CO(n41315));
    SB_LUT4 encoder0_position_31__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n41313), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_19 (.CI(n41313), .I0(n2717), 
            .I1(VCC_net), .CO(n41314));
    SB_LUT4 encoder0_position_31__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n41312), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_18 (.CI(n41312), .I0(n2718), 
            .I1(VCC_net), .CO(n41313));
    SB_LUT4 encoder0_position_31__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n41311), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLA_181 (.Q(INLA_c_0), .C(CLK_c), .E(n29048), .D(GLA_N_384), 
            .R(n29375));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5205));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_DFF dti_counter_2056__i1 (.Q(dti_counter[1]), .C(CLK_c), .D(n54));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_CARRY encoder0_position_31__I_0_add_1838_17 (.CI(n41311), .I0(n2719), 
            .I1(VCC_net), .CO(n41312));
    SB_LUT4 encoder0_position_31__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n41032), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n41310), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5204));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1838_16 (.CI(n41310), .I0(n2720), 
            .I1(VCC_net), .CO(n41311));
    SB_LUT4 encoder0_position_31__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n41309), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_8 (.CI(n40440), .I0(GND_net), .I1(n19_adj_5111), 
            .CO(n40441));
    SB_CARRY encoder0_position_31__I_0_add_1838_15 (.CI(n41309), .I0(n2721), 
            .I1(VCC_net), .CO(n41310));
    SB_LUT4 encoder0_position_31__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n41308), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_14 (.CI(n41308), .I0(n2722), 
            .I1(VCC_net), .CO(n41309));
    SB_CARRY encoder0_position_31__I_0_add_900_3 (.CI(n41032), .I0(n1333), 
            .I1(VCC_net), .CO(n41033));
    SB_LUT4 encoder0_position_31__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n41307), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_13 (.CI(n41307), .I0(n2723), 
            .I1(VCC_net), .CO(n41308));
    SB_LUT4 encoder0_position_31__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n41032));
    SB_LUT4 encoder0_position_31__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n41306), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_12 (.CI(n41306), .I0(n2724), 
            .I1(VCC_net), .CO(n41307));
    SB_LUT4 encoder0_position_31__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n41305), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_11 (.CI(n41305), .I0(n2725), 
            .I1(VCC_net), .CO(n41306));
    SB_LUT4 i37073_4_lut (.I0(n1423), .I1(n1422), .I2(n48931), .I3(n46682), 
            .O(n1455));
    defparam i37073_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1172_3_lut (.I0(n1721), .I1(n1788), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[13]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_238_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[14]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5203));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[15]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5202));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5190));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(delay_counter[28]), .I1(n12_adj_5190), .I2(delay_counter[25]), 
            .I3(delay_counter[30]), .O(n27787));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22956_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n36488));
    defparam i22956_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5201));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_adj_1791 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n27784));
    defparam i2_3_lut_adj_1791.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5200));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1792 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15));
    defparam i6_4_lut_adj_1792.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5199));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(delay_counter[2]), .I2(n14), .I3(delay_counter[6]), 
            .O(n27790));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4275_4_lut (.I0(n27790), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5185));
    defparam i4275_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1793 (.I0(n24_adj_5185), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n47661));
    defparam i2_4_lut_adj_1793.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1794 (.I0(n47661), .I1(delay_counter[18]), .I2(n27784), 
            .I3(GND_net), .O(n47281));
    defparam i2_3_lut_adj_1794.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1795 (.I0(n47281), .I1(delay_counter[23]), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5187));
    defparam i2_4_lut_adj_1795.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5198));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_4_lut_adj_1796 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_5122));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i4_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5197));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_4_lut_adj_1797 (.I0(n7_adj_5187), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n27787), .O(n62));
    defparam i4_4_lut_adj_1797.LUT_INIT = 16'hfffe;
    SB_LUT4 i8273_3_lut (.I0(n62), .I1(\ID_READOUT_FSM.state [0]), .I2(delay_counter[31]), 
            .I3(GND_net), .O(n21721));
    defparam i8273_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i1_2_lut_adj_1798 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5121));
    defparam i1_2_lut_adj_1798.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5196));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut_adj_1799 (.I0(delay_counter[9]), .I1(n4_adj_5121), 
            .I2(delay_counter[10]), .I3(n27790), .O(n47488));
    defparam i2_4_lut_adj_1799.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1800 (.I0(n47488), .I1(n27784), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n47921));
    defparam i2_4_lut_adj_1800.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5237));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5195));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut_adj_1801 (.I0(delay_counter[22]), .I1(n47921), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5238));
    defparam i2_4_lut_adj_1801.LUT_INIT = 16'ha8a0;
    SB_LUT4 i22054_4_lut (.I0(n7_adj_5238), .I1(delay_counter[31]), .I2(n27787), 
            .I3(n8_adj_5237), .O(n1195));   // verilog/TinyFPGA_B.v(378[14:38])
    defparam i22054_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_2_lut (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5119));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1802 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_5118));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i6_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(ID[3]), .I1(n14_adj_5118), .I2(n10_adj_5119), 
            .I3(ID[6]), .O(n27761));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15955_4_lut (.I0(n6662), .I1(n1195), .I2(n21721), .I3(n27762), 
            .O(n29394));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15955_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 encoder0_position_31__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n41304), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_10 (.CI(n41304), .I0(n2726), 
            .I1(VCC_net), .CO(n41305));
    SB_LUT4 encoder0_position_31__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n41303), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_9 (.CI(n41303), .I0(n2727), 
            .I1(VCC_net), .CO(n41304));
    SB_LUT4 encoder0_position_31__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n41302), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_8 (.CI(n41302), .I0(n2728), 
            .I1(VCC_net), .CO(n41303));
    SB_LUT4 encoder0_position_31__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n41301), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_7 (.CI(n41301), .I0(n2729), 
            .I1(GND_net), .CO(n41302));
    SB_LUT4 encoder0_position_31__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n41300), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_6 (.CI(n41300), .I0(n2730), 
            .I1(GND_net), .CO(n41301));
    SB_LUT4 encoder0_position_31__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n41299), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_5 (.CI(n41299), .I0(n2731), 
            .I1(VCC_net), .CO(n41300));
    SB_LUT4 encoder0_position_31__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n41298), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_4 (.CI(n41298), .I0(n2732), 
            .I1(GND_net), .CO(n41299));
    SB_LUT4 encoder0_position_31__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n41297), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_3 (.CI(n41297), .I0(n2733), 
            .I1(VCC_net), .CO(n41298));
    SB_LUT4 i1_2_lut_adj_1803 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n48883));
    defparam i1_2_lut_adj_1803.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n41297));
    SB_LUT4 encoder0_position_31__I_0_add_1771_26_lut (.I0(n52874), .I1(n2610), 
            .I2(VCC_net), .I3(n41296), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i22910_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n36442));
    defparam i22910_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n41295), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1804 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n48883), 
            .O(n48889));
    defparam i1_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1771_25 (.CI(n41295), .I0(n2611), 
            .I1(VCC_net), .CO(n41296));
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n1529), .I1(n48889), .I2(n36442), .I3(n1530), 
            .O(n48891));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_31__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n41294), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_24 (.CI(n41294), .I0(n2612), 
            .I1(VCC_net), .CO(n41295));
    SB_LUT4 encoder0_position_31__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n41293), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37091_4_lut (.I0(n1522), .I1(n1521), .I2(n48891), .I3(n1523), 
            .O(n1554));
    defparam i37091_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_1771_23 (.CI(n41293), .I0(n2613), 
            .I1(VCC_net), .CO(n41294));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i19_3_lut (.I0(encoder0_position[18]), 
            .I1(n15_adj_5098), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n940));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n41292), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_22 (.CI(n41292), .I0(n2614), 
            .I1(VCC_net), .CO(n41293));
    SB_LUT4 encoder0_position_31__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n41291), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_21 (.CI(n41291), .I0(n2615), 
            .I1(VCC_net), .CO(n41292));
    SB_LUT4 encoder0_position_31__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n41290), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_20 (.CI(n41290), .I0(n2616), 
            .I1(VCC_net), .CO(n41291));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i18_3_lut (.I0(encoder0_position[17]), 
            .I1(n16), .I2(encoder0_position[31]), .I3(GND_net), .O(n941));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n41289), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_19 (.CI(n41289), .I0(n2617), 
            .I1(VCC_net), .CO(n41290));
    SB_LUT4 i22729_3_lut (.I0(n941), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n36256));
    defparam i22729_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n41288), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_18 (.CI(n41288), .I0(n2618), 
            .I1(VCC_net), .CO(n41289));
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n1625), .I1(n1627), .I2(n1626), .I3(n1628), 
            .O(n48943));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n41287), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_17 (.CI(n41287), .I0(n2619), 
            .I1(VCC_net), .CO(n41288));
    SB_LUT4 encoder0_position_31__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n41286), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1807 (.I0(n1629), .I1(n36256), .I2(n1630), .I3(n1631), 
            .O(n46691));
    defparam i1_4_lut_adj_1807.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_1771_16 (.CI(n41286), .I0(n2620), 
            .I1(VCC_net), .CO(n41287));
    SB_LUT4 encoder0_position_31__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n41285), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_15 (.CI(n41285), .I0(n2621), 
            .I1(VCC_net), .CO(n41286));
    SB_DFFESR GLB_183 (.Q(INLB_c_0), .C(CLK_c), .E(n29048), .D(GLB_N_398), 
            .R(n29375));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n1623), .I1(n46691), .I2(n1624), .I3(n48943), 
            .O(n48949));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n41284), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_14 (.CI(n41284), .I0(n2622), 
            .I1(VCC_net), .CO(n41285));
    SB_LUT4 i37110_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n48949), 
            .O(n1653_adj_5183));
    defparam i37110_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n41283), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_13 (.CI(n41283), .I0(n2623), 
            .I1(VCC_net), .CO(n41284));
    SB_LUT4 encoder0_position_31__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n41282), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_12 (.CI(n41282), .I0(n2624), 
            .I1(VCC_net), .CO(n41283));
    SB_LUT4 encoder0_position_31__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n41281), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_11 (.CI(n41281), .I0(n2625), 
            .I1(VCC_net), .CO(n41282));
    SB_LUT4 encoder0_position_31__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n41280), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_10 (.CI(n41280), .I0(n2626), 
            .I1(VCC_net), .CO(n41281));
    SB_LUT4 encoder0_position_31__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n41279), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_9 (.CI(n41279), .I0(n2627), 
            .I1(VCC_net), .CO(n41280));
    SB_LUT4 encoder0_position_31__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n41278), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_8 (.CI(n41278), .I0(n2628), 
            .I1(VCC_net), .CO(n41279));
    SB_LUT4 encoder0_position_31__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n41277), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_7 (.CI(n41277), .I0(n2629), 
            .I1(GND_net), .CO(n41278));
    SB_LUT4 encoder0_position_31__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n41276), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_6 (.CI(n41276), .I0(n2630), 
            .I1(GND_net), .CO(n41277));
    SB_LUT4 i5_3_lut_adj_1809 (.I0(control_mode[6]), .I1(n10_adj_5122), 
            .I2(control_mode[2]), .I3(GND_net), .O(n27946));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i5_3_lut_adj_1809.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n41275), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1810 (.I0(n1728), .I1(n1726), .I2(n1727), .I3(GND_net), 
            .O(n48745));
    defparam i1_3_lut_adj_1810.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_31__I_0_add_1771_5 (.CI(n41275), .I0(n2631), 
            .I1(VCC_net), .CO(n41276));
    SB_LUT4 encoder0_position_31__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n41274), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22898_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n36430));
    defparam i22898_4_lut.LUT_INIT = 16'hfcec;
    SB_CARRY encoder0_position_31__I_0_add_1771_4 (.CI(n41274), .I0(n2632), 
            .I1(GND_net), .CO(n41275));
    SB_LUT4 encoder0_position_31__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n41273), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_3 (.CI(n41273), .I0(n2633), 
            .I1(VCC_net), .CO(n41274));
    SB_LUT4 encoder0_position_31__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n41273));
    SB_LUT4 i1_4_lut_adj_1811 (.I0(n1723), .I1(n1724), .I2(n48745), .I3(n1725), 
            .O(n48751));
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1704_25_lut (.I0(n52846), .I1(n2511), 
            .I2(VCC_net), .I3(n41272), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n41271), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_24 (.CI(n41271), .I0(n2512), 
            .I1(VCC_net), .CO(n41272));
    SB_LUT4 encoder0_position_31__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n41270), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(CLK_c), .D(n45417));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n44751));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
           .D(n29594));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1704_23 (.CI(n41270), .I0(n2513), 
            .I1(VCC_net), .CO(n41271));
    SB_LUT4 unary_minus_10_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_5114));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n41269), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5112), 
            .I3(n40439), .O(pwm_setpoint_23__N_191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_22 (.CI(n41269), .I0(n2514), 
            .I1(VCC_net), .CO(n41270));
    SB_LUT4 encoder0_position_31__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n41268), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_21 (.CI(n41268), .I0(n2515), 
            .I1(VCC_net), .CO(n41269));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i28_3_lut (.I0(encoder0_position[27]), 
            .I1(n6_adj_5163), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n41267), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1812 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n48955));
    defparam i1_2_lut_adj_1812.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_31__I_0_add_1704_20 (.CI(n41267), .I0(n2516), 
            .I1(VCC_net), .CO(n41268));
    SB_LUT4 add_2393_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n40552), 
            .O(n7282)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2393_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n41266), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_19 (.CI(n41266), .I0(n2517), 
            .I1(VCC_net), .CO(n41267));
    SB_LUT4 i1_2_lut_adj_1813 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n48901));
    defparam i1_2_lut_adj_1813.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n41265), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1814 (.I0(n927), .I1(n48901), .I2(n928), .I3(n36488), 
            .O(n960));
    defparam i1_4_lut_adj_1814.LUT_INIT = 16'hfefa;
    SB_CARRY encoder0_position_31__I_0_add_1704_18 (.CI(n41265), .I0(n2518), 
            .I1(VCC_net), .CO(n41266));
    SB_LUT4 encoder0_position_31__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n41264), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_17 (.CI(n41264), .I0(n2519), 
            .I1(VCC_net), .CO(n41265));
    SB_LUT4 encoder0_position_31__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n41263), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1704_16 (.CI(n41263), .I0(n2520), 
            .I1(VCC_net), .CO(n41264));
    SB_LUT4 encoder0_position_31__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n41262), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_15 (.CI(n41262), .I0(n2521), 
            .I1(VCC_net), .CO(n41263));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i24_3_lut (.I0(encoder0_position[23]), 
            .I1(n10_adj_5155), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n935));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n41261), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_14 (.CI(n41261), .I0(n2522), 
            .I1(VCC_net), .CO(n41262));
    SB_LUT4 encoder0_position_31__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n41260), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22793_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n36322));
    defparam i22793_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_31__I_0_add_1704_13 (.CI(n41260), .I0(n2523), 
            .I1(VCC_net), .CO(n41261));
    SB_LUT4 encoder0_position_31__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n41259), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1815 (.I0(n1029), .I1(n36322), .I2(n1030), .I3(n1031), 
            .O(n46671));
    defparam i1_4_lut_adj_1815.LUT_INIT = 16'ha080;
    SB_LUT4 i37011_4_lut (.I0(n1026), .I1(n46671), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i37011_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_adj_1816 (.I0(n27765), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5150));   // verilog/TinyFPGA_B.v(268[5:22])
    defparam i1_2_lut_adj_1816.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_31__I_0_i641_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1704_12 (.CI(n41259), .I0(n2524), 
            .I1(VCC_net), .CO(n41260));
    SB_LUT4 encoder0_position_31__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n41258), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i709_3_lut (.I0(n935), .I1(n1101_adj_5181), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_11 (.CI(n41258), .I0(n2525), 
            .I1(VCC_net), .CO(n41259));
    SB_LUT4 encoder0_position_31__I_0_i708_3_lut (.I0(n1033), .I1(n1100_adj_5180), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n41257), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_10 (.CI(n41257), .I0(n2526), 
            .I1(VCC_net), .CO(n41258));
    SB_LUT4 encoder0_position_31__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n41256), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i707_3_lut (.I0(n1032), .I1(n1099_adj_5179), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_9 (.CI(n41256), .I0(n2527), 
            .I1(VCC_net), .CO(n41257));
    SB_LUT4 encoder0_position_31__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n41255), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_8 (.CI(n41255), .I0(n2528), 
            .I1(VCC_net), .CO(n41256));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i23_3_lut (.I0(encoder0_position[22]), 
            .I1(n11_adj_5154), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n936));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1817 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n27946), .I3(GND_net), .O(n15_adj_5124));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i2_3_lut_adj_1817.LUT_INIT = 16'hfdfd;
    SB_LUT4 i22952_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n36484));
    defparam i22952_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1818 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n48879));
    defparam i1_3_lut_adj_1818.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n41254), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1819 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n48911));
    defparam i1_2_lut_adj_1819.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_31__I_0_add_1704_7 (.CI(n41254), .I0(n2529), 
            .I1(GND_net), .CO(n41255));
    SB_LUT4 encoder0_position_31__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n41253), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2393_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n40551), 
            .O(n7283)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2393_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37025_4_lut (.I0(n48911), .I1(n1125), .I2(n48879), .I3(n36484), 
            .O(n1158));
    defparam i37025_4_lut.LUT_INIT = 16'h0103;
    SB_CARRY encoder0_position_31__I_0_add_1704_6 (.CI(n41253), .I0(n2530), 
            .I1(GND_net), .CO(n41254));
    SB_LUT4 encoder0_position_31__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n41252), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i702_3_lut (.I0(n1027), .I1(n1094_adj_5174), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_5 (.CI(n41252), .I0(n2531), 
            .I1(VCC_net), .CO(n41253));
    SB_LUT4 encoder0_position_31__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n41251), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_4 (.CI(n41251), .I0(n2532), 
            .I1(GND_net), .CO(n41252));
    SB_LUT4 encoder0_position_31__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[17]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n41250), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_3 (.CI(n41250), .I0(n2533), 
            .I1(VCC_net), .CO(n41251));
    SB_LUT4 encoder0_position_31__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n41250));
    SB_LUT4 encoder0_position_31__I_0_add_1637_24_lut (.I0(n52807), .I1(n2412), 
            .I2(VCC_net), .I3(n41249), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n41248), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_23 (.CI(n41248), .I0(n2413), 
            .I1(VCC_net), .CO(n41249));
    SB_LUT4 encoder0_position_31__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n41247), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_22 (.CI(n41247), .I0(n2414), 
            .I1(VCC_net), .CO(n41248));
    SB_LUT4 encoder0_position_31__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n41246), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_21 (.CI(n41246), .I0(n2415), 
            .I1(VCC_net), .CO(n41247));
    SB_LUT4 encoder0_position_31__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n41245), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_20 (.CI(n41245), .I0(n2416), 
            .I1(VCC_net), .CO(n41246));
    SB_LUT4 encoder0_position_31__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n41244), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_19 (.CI(n41244), .I0(n2417), 
            .I1(VCC_net), .CO(n41245));
    SB_LUT4 encoder0_position_31__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n41243), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_18 (.CI(n41243), .I0(n2418), 
            .I1(VCC_net), .CO(n41244));
    SB_LUT4 encoder0_position_31__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n41242), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_17 (.CI(n41242), .I0(n2419), 
            .I1(VCC_net), .CO(n41243));
    SB_LUT4 encoder0_position_31__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n41241), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_16 (.CI(n41241), .I0(n2420), 
            .I1(VCC_net), .CO(n41242));
    SB_LUT4 encoder0_position_31__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n41240), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_15 (.CI(n41240), .I0(n2421), 
            .I1(VCC_net), .CO(n41241));
    SB_LUT4 encoder0_position_31__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n41239), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_14 (.CI(n41239), .I0(n2422), 
            .I1(VCC_net), .CO(n41240));
    SB_LUT4 encoder0_position_31__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n41238), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_13 (.CI(n41238), .I0(n2423), 
            .I1(VCC_net), .CO(n41239));
    SB_LUT4 encoder0_position_31__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n41237), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_12 (.CI(n41237), .I0(n2424), 
            .I1(VCC_net), .CO(n41238));
    SB_LUT4 encoder0_position_31__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n41236), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_11 (.CI(n41236), .I0(n2425), 
            .I1(VCC_net), .CO(n41237));
    SB_LUT4 encoder0_position_31__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n41235), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_10 (.CI(n41235), .I0(n2426), 
            .I1(VCC_net), .CO(n41236));
    SB_LUT4 encoder0_position_31__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n41234), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_9 (.CI(n41234), .I0(n2427), 
            .I1(VCC_net), .CO(n41235));
    SB_LUT4 encoder0_position_31__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n41233), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_8 (.CI(n41233), .I0(n2428), 
            .I1(VCC_net), .CO(n41234));
    SB_LUT4 encoder0_position_31__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n41232), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_7 (.CI(n41232), .I0(n2429), 
            .I1(GND_net), .CO(n41233));
    SB_LUT4 encoder0_position_31__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n41231), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_6 (.CI(n41231), .I0(n2430), 
            .I1(GND_net), .CO(n41232));
    SB_LUT4 encoder0_position_31__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n41230), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_5 (.CI(n41230), .I0(n2431), 
            .I1(VCC_net), .CO(n41231));
    SB_LUT4 encoder0_position_31__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n41229), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_4 (.CI(n41229), .I0(n2432), 
            .I1(GND_net), .CO(n41230));
    SB_LUT4 encoder0_position_31__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n41228), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n29854));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n29853));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n29852));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n29851));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n29850));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n29849));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n29848));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(CLK_c), .D(n46452));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1637_3 (.CI(n41228), .I0(n2433), 
            .I1(VCC_net), .CO(n41229));
    SB_LUT4 encoder0_position_31__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n41228));
    SB_CARRY add_2393_6 (.CI(n40551), .I0(n622), .I1(GND_net), .CO(n40552));
    SB_LUT4 encoder0_position_31__I_0_add_1570_23_lut (.I0(n52784), .I1(n2313), 
            .I2(VCC_net), .I3(n41227), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n41226), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_22 (.CI(n41226), .I0(n2314), 
            .I1(VCC_net), .CO(n41227));
    SB_LUT4 unary_minus_10_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5113));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n41225), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF dti_counter_2056__i2 (.Q(dti_counter[2]), .C(CLK_c), .D(n53));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2056__i3 (.Q(dti_counter[3]), .C(CLK_c), .D(n52));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2056__i4 (.Q(dti_counter[4]), .C(CLK_c), .D(n51));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2056__i5 (.Q(dti_counter[5]), .C(CLK_c), .D(n50));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2056__i6 (.Q(dti_counter[6]), .C(CLK_c), .D(n49));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2056__i7 (.Q(dti_counter[7]), .C(CLK_c), .D(n48));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF read_189 (.Q(read), .C(CLK_c), .D(n48551));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n29567));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_mux_3_i29_3_lut (.I0(encoder0_position[28]), 
            .I1(n5_adj_5164), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n516));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dir_175 (.Q(dir), .C(CLK_c), .D(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_CARRY encoder0_position_31__I_0_add_1570_21 (.CI(n41225), .I0(n2315), 
            .I1(VCC_net), .CO(n41226));
    SB_LUT4 add_2393_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n40550), 
            .O(n7284)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2393_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n41224), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_20 (.CI(n41224), .I0(n2316), 
            .I1(VCC_net), .CO(n41225));
    SB_LUT4 encoder0_position_31__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n41223), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_7 (.CI(n40439), .I0(GND_net), .I1(n20_adj_5112), 
            .CO(n40440));
    SB_CARRY encoder0_position_31__I_0_add_1570_19 (.CI(n41223), .I0(n2317), 
            .I1(VCC_net), .CO(n41224));
    SB_LUT4 encoder0_position_31__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n41222), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_18 (.CI(n41222), .I0(n2318), 
            .I1(VCC_net), .CO(n41223));
    SB_CARRY add_2393_5 (.CI(n40550), .I0(n623), .I1(VCC_net), .CO(n40551));
    SB_LUT4 add_2393_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n40549), 
            .O(n7285)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2393_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n41221), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_17 (.CI(n41221), .I0(n2319), 
            .I1(VCC_net), .CO(n41222));
    SB_LUT4 encoder0_position_31__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n41220), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_16 (.CI(n41220), .I0(n2320), 
            .I1(VCC_net), .CO(n41221));
    SB_LUT4 unary_minus_10_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5113), 
            .I3(n40438), .O(pwm_setpoint_23__N_191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n41219), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_15 (.CI(n41219), .I0(n2321), 
            .I1(VCC_net), .CO(n41220));
    SB_CARRY unary_minus_10_add_3_6 (.CI(n40438), .I0(GND_net), .I1(n21_adj_5113), 
            .CO(n40439));
    SB_LUT4 encoder0_position_31__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n41218), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n40397), .O(n1091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_14 (.CI(n41218), .I0(n2322), 
            .I1(VCC_net), .CO(n41219));
    SB_LUT4 encoder0_position_31__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n41217), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_13 (.CI(n41217), .I0(n2323), 
            .I1(VCC_net), .CO(n41218));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i30_3_lut (.I0(encoder0_position[29]), 
            .I1(n4_adj_5165), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_145_19 (.CI(n40397), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n40398));
    SB_LUT4 encoder0_position_31__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n41216), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_12 (.CI(n41216), .I0(n2324), 
            .I1(VCC_net), .CO(n41217));
    SB_CARRY add_145_4 (.CI(n40382), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n40383));
    SB_LUT4 i16016_4_lut (.I0(state_7__N_4103[3]), .I1(data[1]), .I2(n10_adj_5233), 
            .I3(n27954), .O(n29538));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16016_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n41215), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_11 (.CI(n41215), .I0(n2325), 
            .I1(VCC_net), .CO(n41216));
    SB_LUT4 encoder0_position_31__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n41214), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_10 (.CI(n41214), .I0(n2326), 
            .I1(VCC_net), .CO(n41215));
    SB_CARRY add_2393_4 (.CI(n40549), .I0(n516), .I1(GND_net), .CO(n40550));
    SB_LUT4 add_2393_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n40548), 
            .O(n7286)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2393_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2393_3 (.CI(n40548), .I0(n625), .I1(VCC_net), .CO(n40549));
    SB_LUT4 encoder0_position_31__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n41213), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_9 (.CI(n41213), .I0(n2327), 
            .I1(VCC_net), .CO(n41214));
    SB_LUT4 encoder0_position_31__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n41212), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1820 (.I0(n48955), .I1(n1722), .I2(n48751), .I3(n36430), 
            .O(n48755));
    defparam i1_4_lut_adj_1820.LUT_INIT = 16'hfefc;
    SB_LUT4 add_2393_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n7287)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2393_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2393_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n40548));
    SB_CARRY encoder0_position_31__I_0_add_1570_8 (.CI(n41212), .I0(n2328), 
            .I1(VCC_net), .CO(n41213));
    SB_LUT4 encoder0_position_31__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n41211), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_7 (.CI(n41211), .I0(n2329), 
            .I1(GND_net), .CO(n41212));
    SB_LUT4 encoder0_position_31__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n41210), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_6 (.CI(n41210), .I0(n2330), 
            .I1(GND_net), .CO(n41211));
    SB_LUT4 unary_minus_10_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5114), 
            .I3(n40437), .O(pwm_setpoint_23__N_191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n41209), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_5 (.CI(n41209), .I0(n2331), 
            .I1(VCC_net), .CO(n41210));
    SB_LUT4 encoder0_position_31__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n41208), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n40396), .O(n1092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_4 (.CI(n41208), .I0(n2332), 
            .I1(GND_net), .CO(n41209));
    SB_LUT4 encoder0_position_31__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n41207), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_3 (.CI(n41207), .I0(n2333), 
            .I1(VCC_net), .CO(n41208));
    SB_LUT4 encoder0_position_31__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n41207));
    SB_LUT4 encoder0_position_31__I_0_add_1503_22_lut (.I0(n52752), .I1(n2214), 
            .I2(VCC_net), .I3(n41206), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n41205), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_21 (.CI(n41205), .I0(n2215), 
            .I1(VCC_net), .CO(n41206));
    SB_CARRY unary_minus_10_add_3_5 (.CI(n40437), .I0(GND_net), .I1(n22_adj_5114), 
            .CO(n40438));
    SB_LUT4 encoder0_position_31__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n41204), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_20 (.CI(n41204), .I0(n2216), 
            .I1(VCC_net), .CO(n41205));
    SB_LUT4 encoder0_position_31__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n41203), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_19 (.CI(n41203), .I0(n2217), 
            .I1(VCC_net), .CO(n41204));
    SB_LUT4 encoder0_position_31__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n41202), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_18 (.CI(n41202), .I0(n2218), 
            .I1(VCC_net), .CO(n41203));
    SB_LUT4 encoder0_position_31__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n41201), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_8 (.CI(n40386), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n40387));
    SB_CARRY encoder0_position_31__I_0_add_1503_17 (.CI(n41201), .I0(n2219), 
            .I1(VCC_net), .CO(n41202));
    SB_LUT4 encoder0_position_31__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n41200), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_16 (.CI(n41200), .I0(n2220), 
            .I1(VCC_net), .CO(n41201));
    SB_LUT4 encoder0_position_31__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n41199), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5194), .I3(n41931), .O(n2_adj_5167)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5195), .I3(n41930), .O(n3_adj_5166)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_15 (.CI(n41199), .I0(n2221), 
            .I1(VCC_net), .CO(n41200));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_32 (.CI(n41930), 
            .I0(GND_net), .I1(n3_adj_5195), .CO(n41931));
    SB_LUT4 encoder0_position_31__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n41198), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_14 (.CI(n41198), .I0(n2222), 
            .I1(VCC_net), .CO(n41199));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5196), .I3(n41929), .O(n4_adj_5165)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n41197), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_13 (.CI(n41197), .I0(n2223), 
            .I1(VCC_net), .CO(n41198));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_31 (.CI(n41929), 
            .I0(GND_net), .I1(n4_adj_5196), .CO(n41930));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5197), .I3(n41928), .O(n5_adj_5164)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n41196), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_12 (.CI(n41196), .I0(n2224), 
            .I1(VCC_net), .CO(n41197));
    SB_LUT4 encoder0_position_31__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n41195), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_30 (.CI(n41928), 
            .I0(GND_net), .I1(n5_adj_5197), .CO(n41929));
    SB_CARRY encoder0_position_31__I_0_add_1503_11 (.CI(n41195), .I0(n2225), 
            .I1(VCC_net), .CO(n41196));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5198), .I3(n41927), .O(n6_adj_5163)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_29 (.CI(n41927), 
            .I0(GND_net), .I1(n6_adj_5198), .CO(n41928));
    SB_LUT4 encoder0_position_31__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n41194), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5199), .I3(n41926), .O(n7_adj_5162)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_28 (.CI(n41926), 
            .I0(GND_net), .I1(n7_adj_5199), .CO(n41927));
    SB_LUT4 add_145_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n40385), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5200), .I3(n41925), .O(n8_adj_5161)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_10 (.CI(n41194), .I0(n2226), 
            .I1(VCC_net), .CO(n41195));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_27 (.CI(n41925), 
            .I0(GND_net), .I1(n8_adj_5200), .CO(n41926));
    SB_LUT4 encoder0_position_31__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n41193), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5201), .I3(n41924), .O(n9_adj_5158)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_26 (.CI(n41924), 
            .I0(GND_net), .I1(n9_adj_5201), .CO(n41925));
    SB_CARRY encoder0_position_31__I_0_add_1503_9 (.CI(n41193), .I0(n2227), 
            .I1(VCC_net), .CO(n41194));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5202), .I3(n41923), .O(n10_adj_5155)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n41192), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_25 (.CI(n41923), 
            .I0(GND_net), .I1(n10_adj_5202), .CO(n41924));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5203), .I3(n41922), .O(n11_adj_5154)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_24 (.CI(n41922), 
            .I0(GND_net), .I1(n11_adj_5203), .CO(n41923));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5204), .I3(n41921), .O(n12_adj_5151)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_23 (.CI(n41921), 
            .I0(GND_net), .I1(n12_adj_5204), .CO(n41922));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5205), .I3(n41920), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_8 (.CI(n41192), .I0(n2228), 
            .I1(VCC_net), .CO(n41193));
    SB_LUT4 encoder0_position_31__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n41191), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_22 (.CI(n41920), 
            .I0(GND_net), .I1(n13_adj_5205), .CO(n41921));
    SB_CARRY encoder0_position_31__I_0_add_1503_7 (.CI(n41191), .I0(n2229), 
            .I1(GND_net), .CO(n41192));
    SB_LUT4 encoder0_position_31__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n41190), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_6 (.CI(n41190), .I0(n2230), 
            .I1(GND_net), .CO(n41191));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5206), .I3(n41919), .O(n14_adj_5099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n41189), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_21 (.CI(n41919), 
            .I0(GND_net), .I1(n14_adj_5206), .CO(n41920));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5207), .I3(n41918), .O(n15_adj_5098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_20 (.CI(n41918), 
            .I0(GND_net), .I1(n15_adj_5207), .CO(n41919));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5208), .I3(n41917), .O(n16)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_5 (.CI(n41189), .I0(n2231), 
            .I1(VCC_net), .CO(n41190));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_19 (.CI(n41917), 
            .I0(GND_net), .I1(n16_adj_5208), .CO(n41918));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5209), .I3(n41916), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_18 (.CI(n41916), 
            .I0(GND_net), .I1(n17_adj_5209), .CO(n41917));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5210), .I3(n41915), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_17 (.CI(n41915), 
            .I0(GND_net), .I1(n18_adj_5210), .CO(n41916));
    SB_LUT4 encoder0_position_31__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n41188), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5211), .I3(n41914), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_16 (.CI(n41914), 
            .I0(GND_net), .I1(n19_adj_5211), .CO(n41915));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5212), .I3(n41913), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_15 (.CI(n41913), 
            .I0(GND_net), .I1(n20_adj_5212), .CO(n41914));
    SB_CARRY encoder0_position_31__I_0_add_1503_4 (.CI(n41188), .I0(n2232), 
            .I1(GND_net), .CO(n41189));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5213), .I3(n41912), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_14 (.CI(n41912), 
            .I0(GND_net), .I1(n21_adj_5213), .CO(n41913));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5214), .I3(n41911), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5115), 
            .I3(n40436), .O(pwm_setpoint_23__N_191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_13 (.CI(n41911), 
            .I0(GND_net), .I1(n22_adj_5214), .CO(n41912));
    SB_LUT4 encoder0_position_31__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n41187), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_3 (.CI(n41187), .I0(n2233), 
            .I1(VCC_net), .CO(n41188));
    SB_LUT4 encoder0_position_31__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5215), .I3(n41910), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n41187));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_12 (.CI(n41910), 
            .I0(GND_net), .I1(n23_adj_5215), .CO(n41911));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5216), .I3(n41909), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_11 (.CI(n41909), 
            .I0(GND_net), .I1(n24_adj_5216), .CO(n41910));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5217), .I3(n41908), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_10 (.CI(n41908), 
            .I0(GND_net), .I1(n25_adj_5217), .CO(n41909));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5218), .I3(n41907), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_18 (.CI(n40396), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n40397));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_9 (.CI(n41907), 
            .I0(GND_net), .I1(n26_adj_5218), .CO(n41908));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5219), .I3(n41906), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_8 (.CI(n41906), 
            .I0(GND_net), .I1(n27_adj_5219), .CO(n41907));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5220), .I3(n41905), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_7 (.CI(n41905), 
            .I0(GND_net), .I1(n28_adj_5220), .CO(n41906));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5221), .I3(n41904), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_6 (.CI(n41904), 
            .I0(GND_net), .I1(n29_adj_5221), .CO(n41905));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5222), .I3(n41903), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_5 (.CI(n41903), 
            .I0(GND_net), .I1(n30_adj_5222), .CO(n41904));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5223), .I3(n41902), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_4 (.CI(n41902), 
            .I0(GND_net), .I1(n31_adj_5223), .CO(n41903));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5224), .I3(n41901), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_3 (.CI(n41901), 
            .I0(GND_net), .I1(n32_adj_5224), .CO(n41902));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5225), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5225), .CO(n41901));
    SB_CARRY unary_minus_10_add_3_4 (.CI(n40436), .I0(GND_net), .I1(n23_adj_5115), 
            .CO(n40437));
    SB_LUT4 add_145_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n40381), .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5116), 
            .I3(n40435), .O(pwm_setpoint_23__N_191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_3 (.CI(n40435), .I0(GND_net), .I1(n24_adj_5116), 
            .CO(n40436));
    SB_LUT4 encoder0_position_31__I_0_add_1436_21_lut (.I0(n52719), .I1(n2115), 
            .I2(VCC_net), .I3(n41176), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n41175), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n40417), .O(encoder1_position_scaled_23__N_75[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_20 (.CI(n41175), .I0(n2116), 
            .I1(VCC_net), .CO(n41176));
    SB_LUT4 encoder0_position_31__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n41174), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_19 (.CI(n41174), .I0(n2117), 
            .I1(VCC_net), .CO(n41175));
    SB_CARRY add_145_7 (.CI(n40385), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n40386));
    SB_LUT4 encoder0_position_31__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n41173), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_18 (.CI(n41173), .I0(n2118), 
            .I1(VCC_net), .CO(n41174));
    SB_LUT4 unary_minus_10_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n25_adj_5117), 
            .I3(VCC_net), .O(pwm_setpoint_23__N_191[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n41172), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_17 (.CI(n41172), .I0(n2119), 
            .I1(VCC_net), .CO(n41173));
    SB_LUT4 encoder0_position_31__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n41171), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n40395), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_16 (.CI(n41171), .I0(n2120), 
            .I1(VCC_net), .CO(n41172));
    SB_LUT4 encoder0_position_31__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n41170), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_15 (.CI(n41170), .I0(n2121), 
            .I1(VCC_net), .CO(n41171));
    SB_LUT4 encoder0_position_31__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n41169), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_14 (.CI(n41169), .I0(n2122), 
            .I1(VCC_net), .CO(n41170));
    SB_LUT4 encoder0_position_31__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n41168), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_17 (.CI(n40395), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n40396));
    SB_CARRY encoder0_position_31__I_0_add_1436_13 (.CI(n41168), .I0(n2123), 
            .I1(VCC_net), .CO(n41169));
    SB_LUT4 i37135_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n48755), 
            .O(n1752));
    defparam i37135_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n41167), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_12 (.CI(n41167), .I0(n2124), 
            .I1(VCC_net), .CO(n41168));
    SB_LUT4 encoder0_position_31__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n41166), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_CARRY encoder0_position_31__I_0_add_1436_11 (.CI(n41166), .I0(n2125), 
            .I1(VCC_net), .CO(n41167));
    SB_LUT4 encoder0_position_31__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n41165), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_10 (.CI(n41165), .I0(n2126), 
            .I1(VCC_net), .CO(n41166));
    SB_LUT4 encoder0_position_31__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653_adj_5183), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n41164), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_9 (.CI(n41164), .I0(n2127), 
            .I1(VCC_net), .CO(n41165));
    SB_LUT4 encoder0_position_31__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n41163), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5117), 
            .CO(n40435));
    SB_CARRY encoder0_position_31__I_0_add_1436_8 (.CI(n41163), .I0(n2128), 
            .I1(VCC_net), .CO(n41164));
    SB_LUT4 encoder0_position_31__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n41162), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_7 (.CI(n41162), .I0(n2129), 
            .I1(GND_net), .CO(n41163));
    SB_LUT4 encoder0_position_31__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n41161), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_6 (.CI(n41161), .I0(n2130), 
            .I1(GND_net), .CO(n41162));
    SB_LUT4 encoder0_position_31__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n41160), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_5 (.CI(n41160), .I0(n2131), 
            .I1(VCC_net), .CO(n41161));
    SB_LUT4 encoder0_position_31__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n41159), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_4 (.CI(n41159), .I0(n2132), 
            .I1(GND_net), .CO(n41160));
    SB_LUT4 encoder0_position_31__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n41158), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_3 (.CI(n41158), .I0(n2133), 
            .I1(VCC_net), .CO(n41159));
    SB_LUT4 encoder0_position_31__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n40394), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_3 (.CI(n40381), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n40382));
    SB_CARRY encoder0_position_31__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n41158));
    SB_LUT4 encoder0_position_31__I_0_add_1369_20_lut (.I0(n52689), .I1(n2016), 
            .I2(VCC_net), .I3(n41157), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n41156), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_19 (.CI(n41156), .I0(n2017), 
            .I1(VCC_net), .CO(n41157));
    SB_DFFESR GLC_185 (.Q(INLC_c_0), .C(CLK_c), .E(n29048), .D(GLC_N_412), 
            .R(n29375));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n41155), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_18 (.CI(n41155), .I0(n2018), 
            .I1(VCC_net), .CO(n41156));
    SB_LUT4 encoder0_position_31__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n41154), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n40384), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n40434), .O(encoder1_position_scaled_23__N_75[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_16 (.CI(n40394), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n40395));
    SB_LUT4 add_145_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_17 (.CI(n41154), .I0(n2019), 
            .I1(VCC_net), .CO(n41155));
    SB_LUT4 add_145_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n40393), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_15 (.CI(n40393), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n40394));
    SB_LUT4 encoder0_position_31__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n41153), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_16 (.CI(n41153), .I0(n2020), 
            .I1(VCC_net), .CO(n41154));
    SB_LUT4 encoder0_position_31__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n41152), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n40392), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_15 (.CI(n41152), .I0(n2021), 
            .I1(VCC_net), .CO(n41153));
    SB_LUT4 encoder0_position_31__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n41151), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_6 (.CI(n40384), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n40385));
    SB_CARRY encoder0_position_31__I_0_add_1369_14 (.CI(n41151), .I0(n2022), 
            .I1(VCC_net), .CO(n41152));
    SB_LUT4 add_224_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n40433), .O(encoder1_position_scaled_23__N_75[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n41150), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_13 (.CI(n41150), .I0(n2023), 
            .I1(VCC_net), .CO(n41151));
    SB_LUT4 encoder0_position_31__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n41149), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_12 (.CI(n41149), .I0(n2024), 
            .I1(VCC_net), .CO(n41150));
    SB_LUT4 encoder0_position_31__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n41148), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_11 (.CI(n41148), .I0(n2025), 
            .I1(VCC_net), .CO(n41149));
    SB_LUT4 encoder0_position_31__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n41147), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_10 (.CI(n41147), .I0(n2026), 
            .I1(VCC_net), .CO(n41148));
    SB_LUT4 encoder0_position_31__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n41146), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_9 (.CI(n41146), .I0(n2027), 
            .I1(VCC_net), .CO(n41147));
    SB_LUT4 encoder0_position_31__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n41145), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_8 (.CI(n41145), .I0(n2028), 
            .I1(VCC_net), .CO(n41146));
    SB_LUT4 encoder0_position_31__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n41144), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_7 (.CI(n41144), .I0(n2029), 
            .I1(GND_net), .CO(n41145));
    SB_LUT4 encoder0_position_31__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n41143), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_6 (.CI(n41143), .I0(n2030), 
            .I1(GND_net), .CO(n41144));
    SB_LUT4 encoder0_position_31__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n41142), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_5 (.CI(n41142), .I0(n2031), 
            .I1(VCC_net), .CO(n41143));
    SB_LUT4 encoder0_position_31__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n41141), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1369_4 (.CI(n41141), .I0(n2032), 
            .I1(GND_net), .CO(n41142));
    SB_LUT4 encoder0_position_31__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n41140), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_3 (.CI(n41140), .I0(n2033), 
            .I1(VCC_net), .CO(n41141));
    SB_LUT4 encoder0_position_31__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n41140));
    SB_LUT4 encoder0_position_31__I_0_add_1302_19_lut (.I0(n52665), .I1(n1917), 
            .I2(VCC_net), .I3(n41139), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n41138), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_18 (.CI(n41138), .I0(n1918), 
            .I1(VCC_net), .CO(n41139));
    SB_LUT4 encoder0_position_31__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n41137), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_24 (.CI(n40433), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n40434));
    SB_CARRY encoder0_position_31__I_0_add_1302_17 (.CI(n41137), .I0(n1919), 
            .I1(VCC_net), .CO(n41138));
    SB_LUT4 encoder0_position_31__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n41136), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_14 (.CI(n40392), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n40393));
    SB_CARRY encoder0_position_31__I_0_add_1302_16 (.CI(n41136), .I0(n1920), 
            .I1(VCC_net), .CO(n41137));
    SB_LUT4 encoder0_position_31__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n41135), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n40432), .O(encoder1_position_scaled_23__N_75[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_15 (.CI(n41135), .I0(n1921), 
            .I1(VCC_net), .CO(n41136));
    SB_LUT4 encoder0_position_31__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n41134), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_14 (.CI(n41134), .I0(n1922), 
            .I1(VCC_net), .CO(n41135));
    SB_LUT4 encoder0_position_31__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n41133), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_13 (.CI(n41133), .I0(n1923), 
            .I1(VCC_net), .CO(n41134));
    SB_LUT4 encoder0_position_31__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n41132), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_12 (.CI(n41132), .I0(n1924), 
            .I1(VCC_net), .CO(n41133));
    SB_CARRY add_224_23 (.CI(n40432), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n40433));
    SB_LUT4 encoder0_position_31__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n41131), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_11 (.CI(n41131), .I0(n1925), 
            .I1(VCC_net), .CO(n41132));
    SB_CARRY add_145_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n40381));
    SB_LUT4 encoder0_position_31__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n41130), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_10 (.CI(n41130), .I0(n1926), 
            .I1(VCC_net), .CO(n41131));
    SB_LUT4 encoder0_position_31__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n41129), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_CARRY encoder0_position_31__I_0_add_1302_9 (.CI(n41129), .I0(n1927), 
            .I1(VCC_net), .CO(n41130));
    SB_LUT4 encoder0_position_31__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n41128), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_8 (.CI(n41128), .I0(n1928), 
            .I1(VCC_net), .CO(n41129));
    SB_LUT4 encoder0_position_31__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n41127), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_7 (.CI(n41127), .I0(n1929), 
            .I1(GND_net), .CO(n41128));
    SB_LUT4 encoder0_position_31__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n41126), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_12_lut (.I0(n52520), .I1(n1224), 
            .I2(VCC_net), .I3(n40897), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_1302_6 (.CI(n41126), .I0(n1930), 
            .I1(GND_net), .CO(n41127));
    SB_LUT4 encoder0_position_31__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n41125), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_5 (.CI(n41125), .I0(n1931), 
            .I1(VCC_net), .CO(n41126));
    SB_LUT4 encoder0_position_31__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n41124), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_4 (.CI(n41124), .I0(n1932), 
            .I1(GND_net), .CO(n41125));
    SB_LUT4 encoder0_position_31__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n41123), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_3 (.CI(n41123), .I0(n1933), 
            .I1(VCC_net), .CO(n41124));
    SB_LUT4 encoder0_position_31__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n41123));
    SB_LUT4 encoder0_position_31__I_0_add_1235_18_lut (.I0(n52641), .I1(n1818), 
            .I2(VCC_net), .I3(n41122), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_10_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36274_3_lut_4_lut (.I0(n2346), .I1(n2247), .I2(n2228), .I3(n50223), 
            .O(n2426));
    defparam i36274_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16017_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n44527), .I3(GND_net), .O(n29539));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16017_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16018_3_lut (.I0(h3), .I1(reg_B[0]), .I2(n48513), .I3(GND_net), 
            .O(n29540));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i16018_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16019_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n48426), .I3(GND_net), .O(n29541));   // verilog/coms.v(127[12] 300[6])
    defparam i16019_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16020_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29542));   // verilog/coms.v(127[12] 300[6])
    defparam i16020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5132));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5133));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1821 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5193));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_4_lut_adj_1821.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_2_lut_adj_1822 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5149));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i2_2_lut_adj_1822.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1823 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5142));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i6_4_lut_adj_1823.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1824 (.I0(dti_counter[0]), .I1(n14_adj_5142), .I2(n10_adj_5149), 
            .I3(dti_counter[3]), .O(n25316));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i7_4_lut_adj_1824.LUT_INIT = 16'hfffe;
    SB_LUT4 i36997_2_lut (.I0(n25316), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_416));
    defparam i36997_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i16149_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n48426), .I3(GND_net), .O(n29671));   // verilog/coms.v(127[12] 300[6])
    defparam i16149_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16084_3_lut (.I0(h1), .I1(reg_B[2]), .I2(n48513), .I3(GND_net), 
            .O(n29606));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i16084_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16085_4_lut (.I0(state_7__N_4103[3]), .I1(data[3]), .I2(n4_adj_5120), 
            .I3(n27954), .O(n29607));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16085_4_lut.LUT_INIT = 16'hccca;
    motorControl control (.GND_net(GND_net), .setpoint({setpoint}), .motor_state({motor_state}), 
            .\Ki[11] (Ki[11]), .\Ki[14] (Ki[14]), .\Ki[12] (Ki[12]), .\Ki[3] (Ki[3]), 
            .\Ki[4] (Ki[4]), .\Ki[15] (Ki[15]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), 
            .\Kp[2] (Kp[2]), .\Ki[5] (Ki[5]), .\Ki[13] (Ki[13]), .\Ki[0] (Ki[0]), 
            .\Ki[1] (Ki[1]), .\Ki[6] (Ki[6]), .\Ki[2] (Ki[2]), .\Kp[3] (Kp[3]), 
            .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .IntegralLimit({IntegralLimit}), 
            .\Kp[7] (Kp[7]), .duty({duty}), .clk32MHz(clk32MHz), .\Ki[7] (Ki[7]), 
            .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .VCC_net(VCC_net), 
            .PWMLimit({PWMLimit}), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), 
            .\Kp[15] (Kp[15])) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(271[16] 283[4])
    SB_LUT4 i16086_3_lut (.I0(h2), .I1(reg_B[1]), .I2(n48513), .I3(GND_net), 
            .O(n29608));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i16086_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16087_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n44527), .I3(GND_net), .O(n29609));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16087_3_lut.LUT_INIT = 16'hacac;
    \quadrature_decoder(1,500000)_U0  quad_counter0 (.\a_new[1] (a_new[1]), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .n1653(CLK_c), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .b_prev(b_prev), .direction_N_3907(direction_N_3907), .encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .n29600(n29600), .n1617(n1617), .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(285[57] 292[6])
    SB_LUT4 i16088_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n44527), .I3(GND_net), .O(n29610));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16088_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16089_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n44527), .I3(GND_net), .O(n29611));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16089_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16090_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n44527), .I3(GND_net), .O(n29612));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16090_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16091_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n44527), .I3(GND_net), .O(n29613));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16091_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16092_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n44527), .I3(GND_net), .O(n29614));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16092_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16093_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n44527), .I3(GND_net), .O(n29615));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16093_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16094_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n44527), .I3(GND_net), .O(n29616));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16094_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16095_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n44527), .I3(GND_net), .O(n29617));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16095_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16096_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n44527), .I3(GND_net), .O(n29618));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16096_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16097_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n44527), .I3(GND_net), .O(n29619));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16097_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5134));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36019_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5193), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[0]), .O(n51311));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i36019_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i35971_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5193), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[1]), .O(n51320));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i35971_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i36027_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5193), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[2]), .O(n51321));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i36027_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i36026_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5193), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[3]), .O(n51322));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i36026_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i36025_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5193), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[4]), .O(n51323));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i36025_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i36024_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5193), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[5]), .O(n51324));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i36024_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i36023_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5193), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[6]), .O(n51325));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i36023_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i36022_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5193), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[7]), .O(n51326));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i36022_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i1_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5193), 
            .I2(commutation_state_prev[0]), .I3(dti_N_416), .O(n29044));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 unary_minus_10_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5135));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5305[1]), .I1(r_SM_Main_adj_5305[0]), 
            .I2(r_SM_Main_adj_5305[2]), .I3(r_SM_Main_2__N_3613[1]), .O(n53403));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5136));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5137));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31089_4_lut_4_lut_4_lut (.I0(h1), .I1(h3), .I2(h2), .I3(commutation_state[2]), 
            .O(n46452));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i31089_4_lut_4_lut_4_lut.LUT_INIT = 16'hc544;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5138));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_3_lut (.I0(h1), .I1(h3), .I2(h2), .I3(GND_net), 
            .O(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n29137), 
            .I3(rx_data_ready), .O(n45179));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3542[2]), .O(n45591));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5139));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5140));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5102));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5141));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13_3_lut_4_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3542[2]), .O(n29137));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13_3_lut_4_lut_4_lut.LUT_INIT = 16'h4303;
    SB_LUT4 unary_minus_10_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21762_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(84[16:31])
    defparam i21762_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21761_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(82[16:31])
    defparam i21761_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22131_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(80[16:31])
    defparam i22131_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16022_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(n29252), 
            .I3(state_3__N_528[1]), .O(n29544));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16022_4_lut_4_lut.LUT_INIT = 16'hfc7c;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5143));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5144));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i701_3_lut (.I0(n1026), .I1(n1093_adj_5173), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5145));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i706_3_lut (.I0(n1031), .I1(n1098_adj_5178), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5146));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15847_2_lut (.I0(n29048), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n29375));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i15847_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36845_4_lut (.I0(commutation_state[1]), .I1(n25316), .I2(dti), 
            .I3(commutation_state[2]), .O(n29048));
    defparam i36845_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 encoder0_position_31__I_0_i705_3_lut (.I0(n1030), .I1(n1097_adj_5177), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i704_3_lut (.I0(n1029), .I1(n1096_adj_5176), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i703_3_lut (.I0(n1028), .I1(n1095_adj_5175), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16098_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n44527), .I3(GND_net), .O(n29620));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16098_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1825 (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_5122), .I3(control_mode[2]), .O(n27765));   // verilog/TinyFPGA_B.v(268[5:22])
    defparam i1_2_lut_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 i31034_3_lut (.I0(n4_adj_5165), .I1(n7284), .I2(n46394), .I3(GND_net), 
            .O(n46395));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31035_3_lut (.I0(encoder0_position[29]), .I1(n46395), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6635_3_lut_4_lut_4_lut (.I0(commutation_state[1]), .I1(commutation_state[2]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_367));
    defparam i6635_3_lut_4_lut_4_lut.LUT_INIT = 16'h1a14;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i27_3_lut (.I0(encoder0_position[26]), 
            .I1(n7_adj_5162), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1826 (.I0(n4_adj_5165), .I1(n5_adj_5164), .I2(n731), 
            .I3(n6_adj_5163), .O(n5_adj_5123));
    defparam i1_4_lut_adj_1826.LUT_INIT = 16'heeea;
    SB_LUT4 i16033_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_5101), 
            .I3(n27898), .O(n29555));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16033_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i6637_3_lut_4_lut_4_lut (.I0(commutation_state[1]), .I1(commutation_state[2]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_384));
    defparam i6637_3_lut_4_lut_4_lut.LUT_INIT = 16'ha141;
    SB_LUT4 i16034_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_5096), 
            .I3(n27903), .O(n29556));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16034_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16035_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_5096), 
            .I3(n27898), .O(n29557));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16035_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16036_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_5156), 
            .I3(n27903), .O(n29558));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16036_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16037_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_5156), 
            .I3(n27898), .O(n29559));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16037_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16038_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n35507), 
            .I3(n27903), .O(n29560));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16038_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16039_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n35507), 
            .I3(n27898), .O(n29561));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16039_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16041_4_lut (.I0(state_7__N_4103[3]), .I1(data[0]), .I2(n10_adj_5233), 
            .I3(n27911), .O(n29563));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16041_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16042_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n48426), 
            .I3(GND_net), .O(n29564));   // verilog/coms.v(127[12] 300[6])
    defparam i16042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16043_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n48426), 
            .I3(GND_net), .O(n29565));   // verilog/coms.v(127[12] 300[6])
    defparam i16043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5147));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16044_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n29106), .I3(GND_net), .O(n29566));   // verilog/coms.v(127[12] 300[6])
    defparam i16044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16045_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n48489), .I3(GND_net), 
            .O(n29567));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16047_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n48426), .I3(GND_net), .O(n29569));   // verilog/coms.v(127[12] 300[6])
    defparam i16047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_scaled_23__I_4_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_279));   // verilog/TinyFPGA_B.v(321[33:52])
    defparam encoder1_position_scaled_23__I_4_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i16048_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n48426), .I3(GND_net), .O(n29570));   // verilog/coms.v(127[12] 300[6])
    defparam i16048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31052_2_lut (.I0(n114), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n46413));
    defparam i31052_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1827 (.I0(n3_adj_5166), .I1(n2_adj_5167), .I2(n5_adj_5123), 
            .I3(GND_net), .O(n46394));
    defparam i1_3_lut_adj_1827.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_1828 (.I0(n113), .I1(n45520), .I2(n3303), .I3(n46413), 
            .O(n48537));
    defparam i2_4_lut_adj_1828.LUT_INIT = 16'hcdff;
    SB_LUT4 i1_4_lut_adj_1829 (.I0(n63), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n48537), .I3(n25059), .O(n44955));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1829.LUT_INIT = 16'hd5f5;
    SB_LUT4 i3_4_lut_adj_1830 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n48551));
    defparam i3_4_lut_adj_1830.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_1831 (.I0(enable_slow_N_4190), .I1(data_ready), 
            .I2(state_adj_5296[1]), .I3(state_adj_5296[0]), .O(n45289));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1831.LUT_INIT = 16'hccd0;
    SB_LUT4 i16053_4_lut (.I0(rw), .I1(state_adj_5296[0]), .I2(state_adj_5296[1]), 
            .I3(n5741), .O(n29575));   // verilog/eeprom.v(26[8] 58[4])
    defparam i16053_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i16057_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5305[1]), .I2(n20247), 
            .I3(n4), .O(n29579));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i16057_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i16061_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_4087[0]), 
            .I3(enable_slow_N_4190), .O(n29583));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16061_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i21914_1_lut_2_lut (.I0(n25316), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n1910));
    defparam i21914_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i16078_3_lut_4_lut (.I0(n1617), .I1(b_prev), .I2(a_new[1]), 
            .I3(direction_N_3907), .O(n29600));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16078_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i21771_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27761), .I3(n1195), .O(n35272));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i21771_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfbb;
    SB_LUT4 i1_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27761), .I3(GND_net), .O(n27762));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1832 (.I0(\ID_READOUT_FSM.state [0]), 
            .I1(\ID_READOUT_FSM.state [1]), .I2(n27761), .I3(n1195), .O(n6970));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_2_lut_3_lut_4_lut_adj_1832.LUT_INIT = 16'h0400;
    SB_LUT4 i1_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27761), .I3(GND_net), .O(n6662));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 mux_236_i19_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i20_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i21_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i22_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i23_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i24_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5148));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16069_3_lut_4_lut (.I0(n1658), .I1(b_prev_adj_5153), .I2(a_new_adj_5272[1]), 
            .I3(direction_N_3907_adj_5157), .O(n29591));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16069_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 mux_236_i1_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), .I2(motor_state_23__N_123[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_236_i2_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), .I2(motor_state_23__N_123[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i3_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), .I2(motor_state_23__N_123[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i4_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), .I2(motor_state_23__N_123[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i5_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), .I2(motor_state_23__N_123[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    \grp_debouncer(3,1000)  debounce (.reg_B({reg_B}), .CLK_c(CLK_c), .GND_net(GND_net), 
            .VCC_net(VCC_net), .n29608(n29608), .data_o({h1, h2, h3}), 
            .n29606(n29606), .data_i({hall1, hall2, hall3}), .n48513(n48513), 
            .n29540(n29540));   // verilog/TinyFPGA_B.v(98[26] 102[3])
    SB_LUT4 mux_236_i6_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), .I2(motor_state_23__N_123[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i31040_3_lut (.I0(n3_adj_5166), .I1(n7283), .I2(n46394), .I3(GND_net), 
            .O(n46401));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i7_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), .I2(motor_state_23__N_123[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i31041_3_lut (.I0(encoder0_position[30]), .I1(n46401), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i31041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i8_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), .I2(motor_state_23__N_123[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i9_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), .I2(motor_state_23__N_123[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i10_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i11_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i12_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i13_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_5316[0]), .I1(n51345), .I2(n6387), 
            .I3(n10), .O(n8_adj_5184));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_LUT4 i22958_4_lut (.I0(n834), .I1(n831), .I2(n832), .I3(n833), 
            .O(n36490));
    defparam i22958_4_lut.LUT_INIT = 16'hfcec;
    coms neopxl_color_23__I_0 (.CLK_c(CLK_c), .n122(n122), .GND_net(GND_net), 
         .n63(n63_adj_5188), .n3684(n3684), .n8(n8_adj_5192), .n3303(n3303), 
         .\FRAME_MATCHER.state_31__N_2788[2] (\FRAME_MATCHER.state_31__N_2788 [2]), 
         .\FRAME_MATCHER.i_31__N_2626 (\FRAME_MATCHER.i_31__N_2626 ), .n4452(n4452), 
         .n7(n7_adj_5191), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .\data_in[1] ({\data_in[1] }), 
         .\data_in[0] ({\data_in[0] }), .\data_in[3] ({\data_in[3] }), .\data_in[2] ({\data_in[2] }), 
         .n771(n771), .n29106(n29106), .n29671(n29671), .control_mode({control_mode}), 
         .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), .n63_adj_10(n63), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .n48070(n48070), 
         .n29670(n29670), .n29669(n29669), .n29668(n29668), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .n29667(n29667), 
         .n25095(n25095), .n29666(n29666), .n29665(n29665), .n29664(n29664), 
         .PWMLimit({PWMLimit}), .n29663(n29663), .rx_data_ready(rx_data_ready), 
         .setpoint({setpoint}), .n29662(n29662), .n29661(n29661), .n29660(n29660), 
         .n29659(n29659), .n29658(n29658), .n29657(n29657), .n29656(n29656), 
         .n29655(n29655), .\data_out_frame[8] ({\data_out_frame[8] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .n29654(n29654), .n29653(n29653), .n29652(n29652), .n29651(n29651), 
         .n29650(n29650), .n29649(n29649), .n29648(n29648), .n29647(n29647), 
         .n29646(n29646), .n29645(n29645), .n29644(n29644), .n29643(n29643), 
         .n29642(n29642), .n53344(n53344), .n53345(n53345), .DE_c(DE_c), 
         .LED_c(LED_c), .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .rx_data({rx_data}), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .\data_in_frame[3] ({\data_in_frame[3] }), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .tx_active(tx_active), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .\state[2] (state_adj_5316[2]), 
         .\state[3] (state_adj_5316[3]), .n10(n10_adj_5100), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .n30122(n30122), .IntegralLimit({IntegralLimit}), 
         .n30121(n30121), .n30120(n30120), .n30119(n30119), .n30118(n30118), 
         .n30117(n30117), .n30116(n30116), .n30115(n30115), .n30114(n30114), 
         .n30113(n30113), .n30112(n30112), .n30111(n30111), .n30110(n30110), 
         .n30109(n30109), .n30108(n30108), .n30107(n30107), .n30106(n30106), 
         .n30105(n30105), .n30104(n30104), .n30103(n30103), .n30102(n30102), 
         .n30101(n30101), .n30100(n30100), .n30099(n30099), .n30098(n30098), 
         .n30097(n30097), .n30096(n30096), .n30095(n30095), .n30094(n30094), 
         .n30093(n30093), .n30092(n30092), .n30091(n30091), .n30090(n30090), 
         .n30089(n30089), .n30088(n30088), .n30087(n30087), .n30086(n30086), 
         .n30085(n30085), .n30084(n30084), .n30083(n30083), .n30082(n30082), 
         .n30081(n30081), .n30080(n30080), .n30079(n30079), .n30078(n30078), 
         .n30077(n30077), .n30076(n30076), .n30075(n30075), .n30074(n30074), 
         .n30073(n30073), .n30072(n30072), .n30071(n30071), .n30070(n30070), 
         .n30069(n30069), .n30068(n30068), .\Kp[1] (Kp[1]), .n30067(n30067), 
         .\Kp[2] (Kp[2]), .n30066(n30066), .\Kp[3] (Kp[3]), .n30065(n30065), 
         .\Kp[4] (Kp[4]), .n30064(n30064), .\Kp[5] (Kp[5]), .n30063(n30063), 
         .\Kp[6] (Kp[6]), .n30062(n30062), .\Kp[7] (Kp[7]), .n30061(n30061), 
         .\Kp[8] (Kp[8]), .n30060(n30060), .\Kp[9] (Kp[9]), .n30059(n30059), 
         .\Kp[10] (Kp[10]), .n30058(n30058), .\Kp[11] (Kp[11]), .n30057(n30057), 
         .\Kp[12] (Kp[12]), .n30056(n30056), .\Kp[13] (Kp[13]), .n30055(n30055), 
         .\Kp[14] (Kp[14]), .n30054(n30054), .\Kp[15] (Kp[15]), .n30053(n30053), 
         .\Ki[1] (Ki[1]), .n30052(n30052), .\Ki[2] (Ki[2]), .n30051(n30051), 
         .\Ki[3] (Ki[3]), .n30050(n30050), .\Ki[4] (Ki[4]), .n30049(n30049), 
         .\Ki[5] (Ki[5]), .n30048(n30048), .\Ki[6] (Ki[6]), .n30047(n30047), 
         .\Ki[7] (Ki[7]), .n30046(n30046), .\Ki[8] (Ki[8]), .n30045(n30045), 
         .\Ki[9] (Ki[9]), .n30044(n30044), .\Ki[10] (Ki[10]), .n30043(n30043), 
         .\Ki[11] (Ki[11]), .n30042(n30042), .\Ki[12] (Ki[12]), .n30041(n30041), 
         .\Ki[13] (Ki[13]), .n30040(n30040), .\Ki[14] (Ki[14]), .n30039(n30039), 
         .\Ki[15] (Ki[15]), .n30038(n30038), .n30037(n30037), .n30036(n30036), 
         .n30035(n30035), .n30034(n30034), .n30033(n30033), .n30032(n30032), 
         .n30031(n30031), .n30030(n30030), .n30029(n30029), .n30028(n30028), 
         .n30027(n30027), .n30026(n30026), .n30025(n30025), .n30024(n30024), 
         .n30023(n30023), .n30022(n30022), .n30021(n30021), .n30020(n30020), 
         .n30019(n30019), .n30018(n30018), .n30017(n30017), .n30016(n30016), 
         .n30015(n30015), .n30014(n30014), .n30013(n30013), .n30012(n30012), 
         .n30011(n30011), .n30010(n30010), .n30009(n30009), .n30008(n30008), 
         .n30007(n30007), .n30006(n30006), .n30005(n30005), .n30004(n30004), 
         .n30003(n30003), .n30002(n30002), .n30001(n30001), .n30000(n30000), 
         .n29999(n29999), .n29998(n29998), .n29997(n29997), .n29996(n29996), 
         .n29995(n29995), .n29994(n29994), .n29993(n29993), .n29991(n29991), 
         .n29990(n29990), .n29989(n29989), .n29988(n29988), .n29987(n29987), 
         .n29986(n29986), .n29985(n29985), .n29984(n29984), .n29983(n29983), 
         .n29982(n29982), .n29981(n29981), .n29980(n29980), .n29979(n29979), 
         .n29978(n29978), .n29977(n29977), .n29976(n29976), .n29975(n29975), 
         .n29974(n29974), .n29973(n29973), .n29972(n29972), .n29971(n29971), 
         .n29970(n29970), .n29969(n29969), .n29968(n29968), .n29967(n29967), 
         .n29966(n29966), .n29965(n29965), .n29964(n29964), .n29963(n29963), 
         .n29962(n29962), .n29961(n29961), .n29960(n29960), .n29959(n29959), 
         .n29958(n29958), .n29957(n29957), .n29956(n29956), .n29955(n29955), 
         .n29954(n29954), .n29953(n29953), .n29952(n29952), .n29951(n29951), 
         .n29950(n29950), .n29949(n29949), .n29948(n29948), .n29947(n29947), 
         .n29946(n29946), .n29945(n29945), .n29944(n29944), .n29943(n29943), 
         .n29942(n29942), .n29941(n29941), .n29940(n29940), .n29939(n29939), 
         .n29938(n29938), .n29937(n29937), .n29936(n29936), .n29935(n29935), 
         .n29934(n29934), .n29933(n29933), .n29932(n29932), .n29931(n29931), 
         .n29930(n29930), .n29929(n29929), .n29928(n29928), .n29927(n29927), 
         .n29926(n29926), .n29925(n29925), .n29924(n29924), .n29923(n29923), 
         .n29922(n29922), .n29921(n29921), .n29920(n29920), .n29919(n29919), 
         .n29918(n29918), .n29917(n29917), .n29916(n29916), .n29915(n29915), 
         .n29914(n29914), .n29913(n29913), .n29912(n29912), .n29911(n29911), 
         .n29910(n29910), .n29909(n29909), .n29908(n29908), .n29907(n29907), 
         .n29906(n29906), .n29905(n29905), .n29904(n29904), .n29903(n29903), 
         .n29902(n29902), .n29901(n29901), .n29900(n29900), .n29899(n29899), 
         .n29898(n29898), .n29897(n29897), .n29896(n29896), .n29895(n29895), 
         .n29894(n29894), .n29893(n29893), .n29892(n29892), .n29891(n29891), 
         .n29890(n29890), .n29889(n29889), .n29888(n29888), .n29887(n29887), 
         .n29886(n29886), .n29885(n29885), .n29884(n29884), .n29883(n29883), 
         .n29882(n29882), .n29881(n29881), .n29880(n29880), .n29879(n29879), 
         .n29878(n29878), .n29877(n29877), .neopxl_color({neopxl_color}), 
         .n29876(n29876), .n29875(n29875), .n29874(n29874), .n29873(n29873), 
         .n29872(n29872), .n29871(n29871), .n29870(n29870), .n29869(n29869), 
         .n29868(n29868), .n29867(n29867), .n29866(n29866), .n29865(n29865), 
         .n29864(n29864), .n29863(n29863), .n29862(n29862), .n29861(n29861), 
         .n29860(n29860), .n29859(n29859), .n29858(n29858), .n29857(n29857), 
         .n29856(n29856), .n29855(n29855), .n44955(n44955), .n29570(n29570), 
         .n29569(n29569), .n29566(n29566), .n29565(n29565), .\Ki[0] (Ki[0]), 
         .n29564(n29564), .\Kp[0] (Kp[0]), .n29542(n29542), .n29541(n29541), 
         .n25059(n25059), .n123(n123), .ID({ID}), .n48426(n48426), .n45588(n45588), 
         .n113(n113), .n114(n114), .\state[0] (state_adj_5316[0]), .n6935(n6935), 
         .n29165(n29165), .tx_o(tx_o), .r_SM_Main({r_SM_Main_adj_5305}), 
         .\r_SM_Main_2__N_3613[1] (r_SM_Main_2__N_3613[1]), .\r_Bit_Index[0] (r_Bit_Index_adj_5307[0]), 
         .n45528(n45528), .n29578(n29578), .n29579(n29579), .n53403(n53403), 
         .VCC_net(VCC_net), .n20247(n20247), .n4(n4), .tx_enable(tx_enable), 
         .n29175(n29175), .r_SM_Main_adj_18({r_SM_Main}), .r_Rx_Data(r_Rx_Data), 
         .RX_N_10(RX_N_10), .\r_SM_Main_2__N_3542[2] (r_SM_Main_2__N_3542[2]), 
         .\r_Bit_Index[0]_adj_14 (r_Bit_Index[0]), .n27903(n27903), .n4_adj_15(n4_adj_5101), 
         .n45526(n45526), .n29587(n29587), .n29582(n29582), .n45179(n45179), 
         .n29561(n29561), .n29560(n29560), .n29559(n29559), .n29558(n29558), 
         .n29557(n29557), .n29556(n29556), .n29555(n29555), .n45591(n45591), 
         .n4_adj_16(n4_adj_5096), .n4_adj_17(n4_adj_5156), .n27898(n27898), 
         .n35507(n35507)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(238[8] 261[4])
    SB_LUT4 mux_238_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[0]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_236_i14_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i15_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i16_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i17_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[16]), .I3(encoder0_position_scaled[16]), 
            .O(motor_state[16]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i23085_4_lut (.I0(n829), .I1(n828), .I2(n36490), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i23085_4_lut.LUT_INIT = 16'heccc;
    EEPROM eeprom (.CLK_c(CLK_c), .enable_slow_N_4190(enable_slow_N_4190), 
           .\state[1] (state_adj_5296[1]), .n5740({n5741}), .\state[0] (state_adj_5296[0]), 
           .GND_net(GND_net), .\state[3] (state_adj_5316[3]), .\state[0]_adj_4 (state_adj_5316[0]), 
           .read(read), .\state[2] (state_adj_5316[2]), .n29575(n29575), 
           .rw(rw), .n45289(n45289), .data_ready(data_ready), .n6387(n6387), 
           .sda_enable(sda_enable), .\state_7__N_4087[0] (state_7__N_4087[0]), 
           .n51345(n51345), .n10(n10), .n27911(n27911), .n27954(n27954), 
           .scl_enable(scl_enable), .n29607(n29607), .data({data}), .n35513(n35513), 
           .n4(n4_adj_5097), .n29598(n29598), .n29597(n29597), .n29596(n29596), 
           .n29595(n29595), .VCC_net(VCC_net), .\state_7__N_4103[3] (state_7__N_4103[3]), 
           .n6935(n6935), .\saved_addr[0] (saved_addr[0]), .n10_adj_5(n10_adj_5100), 
           .n10_adj_6(n10_adj_5233), .n8(n8_adj_5184), .scl(scl), .n30125(n30125), 
           .sda_out(sda_out), .n29583(n29583), .n29563(n29563), .n29538(n29538), 
           .n4_adj_7(n4_adj_5120)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(387[10] 398[6])
    SB_LUT4 mux_238_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5124), .I3(n15_adj_5150), .O(motor_state_23__N_123[1]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i2_4_lut.LUT_INIT = 16'h0aca;
    \quadrature_decoder(1,500000)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .\a_new[1] (a_new_adj_5272[1]), .ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1653(CLK_c), .ENCODER1_A_N_keep(ENCODER1_A_N), .VCC_net(VCC_net), 
            .b_prev(b_prev_adj_5153), .direction_N_3907(direction_N_3907_adj_5157), 
            .n29591(n29591), .n1658(n1658)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(294[57] 301[6])
    SB_LUT4 mux_236_i18_3_lut_4_lut (.I0(n27765), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16099_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n44527), .I3(GND_net), .O(n29621));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16099_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16100_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n44527), .I3(GND_net), .O(n29622));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16100_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16101_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n44527), .I3(GND_net), .O(n29623));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16102_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n44527), .I3(GND_net), .O(n29624));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16102_3_lut.LUT_INIT = 16'hacac;
    pwm PWM (.pwm_setpoint({pwm_setpoint}), .GND_net(GND_net), .pwm_out(pwm_out), 
        .clk32MHz(clk32MHz), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    SB_LUT4 i16103_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n44527), .I3(GND_net), .O(n29625));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16104_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n44527), .I3(GND_net), .O(n29626));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16105_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n44527), .I3(GND_net), .O(n29627));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16106_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n44527), .I3(GND_net), .O(n29628));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16106_3_lut.LUT_INIT = 16'hacac;
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (\state[0] , \state[1] , n44527, 
            GND_net, CLK_c, VCC_net, timer, n29252, neopxl_color, 
            n29639, \neo_pixel_transmitter.t0 , n29638, n29637, n29636, 
            n29635, n29634, n29633, n29632, n29631, n29630, n29629, 
            n29628, n29627, n29626, n29625, n29624, n29623, n29622, 
            n29621, n29620, n29619, n29618, n29617, n29616, n29615, 
            n29614, n29613, n29612, n29611, n29610, n29609, \state_3__N_528[1] , 
            LED_c, n29544, n29539, NEOPXL_c) /* synthesis syn_module_defined=1 */ ;
    output \state[0] ;
    output \state[1] ;
    output n44527;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output [31:0]timer;
    output n29252;
    input [23:0]neopxl_color;
    input n29639;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input n29638;
    input n29637;
    input n29636;
    input n29635;
    input n29634;
    input n29633;
    input n29632;
    input n29631;
    input n29630;
    input n29629;
    input n29628;
    input n29627;
    input n29626;
    input n29625;
    input n29624;
    input n29623;
    input n29622;
    input n29621;
    input n29620;
    input n29619;
    input n29618;
    input n29617;
    input n29616;
    input n29615;
    input n29614;
    input n29613;
    input n29612;
    input n29611;
    input n29610;
    input n29609;
    output \state_3__N_528[1] ;
    input LED_c;
    input n29544;
    input n29539;
    output NEOPXL_c;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n27768, n4, n42258, n46573, \neo_pixel_transmitter.done , 
        start, n7, n8, n46580;
    wire [31:0]n133;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n41761, n41762, n41760, n41759, \neo_pixel_transmitter.done_N_736 , 
        n53316, n41758, start_N_727, n7_adj_4944, n41757, n41756;
    wire [31:0]n133_adj_5095;
    
    wire n41755, n41754, n2589;
    wire [31:0]n2654;
    
    wire n2621, n2688, n2604, n2703, n2600, n2699, n41753, n2605, 
        n2704, n2602, n2701, n2607, n2706, n2606, n2705, n2598, 
        n2697, n2601, n2700, n2609, n2708, n2603, n2702, n2608, 
        n2707, n2597, n2696, n2595, n2694, n2596, n2695, n2594, 
        n2693, n2593, n2692, n2591, n2690, n2592, n2691, n2590, 
        n2689, n2709, n2599, n2698, n30, n41752, n41751, n41750, 
        n41749, n41748, n37, n36, n42, n41747, n41746, n41745, 
        n41744, n41743, n41742, n40, n2687, n41, n41741, n41740, 
        n41739, n41738, n39, n2720, n41737, n6801, n6, n29377, 
        n29446, n41736, n2499;
    wire [31:0]n2555;
    
    wire n2522, n2509, n2502, n2507, n2498, n2508, n2505, n2496, 
        n2504, n2500, n2501, n2503, n2506, n2494, n2495, n2493, 
        n2492, n2491, n2490, n2497, n28, n35, n2588, n34, n40_adj_4960, 
        n38, n39_adj_4961, n37_adj_4962, n41735, n41734, n2407;
    wire [31:0]n2456;
    
    wire n2423, n2409, n2406, n41733, n2404, n2400, n2399, n2397, 
        n2398, n2396, n2395, n2393, n2394, n2392, n2405, n2403, 
        n2401, n2408, n41732, n2402, n2391, n2489, n22, n36_adj_4963, 
        n27, n34_adj_4964, n33, n37_adj_4965, n39_adj_4966, n41731, 
        n41730, n41729, n41728, n41727, n41726, n41725, n1400, 
        n1301, n41717, n1334;
    wire [31:0]n1367;
    
    wire n1302, n41716, n1303, n41715, n1304, n41714;
    wire [31:0]one_wire_N_679;
    
    wire n27952, n36444, n1305, n41713, n1306, n41712, n1307, 
        n41711, n1308, n41710, n4_adj_4976, n1309, n41709, n50005, 
        n50011, n51335, n46581, n2307;
    wire [31:0]n2357;
    
    wire n2324, n2298, n2302, n2303, n2308, n2300, n2294, n2293, 
        n2292, n2297, n2296, n2301, n2295, n2299, n2306, n2309, 
        n46472, n45634, n103, n2305, n2304, n34_adj_4981, n25, 
        n32, n2390, n31, n35_adj_4982, n37_adj_4983, n16, n2201;
    wire [31:0]n2258;
    
    wire n2225, n6_adj_4984, n2199, n2200, n2198, n2204, n2207, 
        n2203, n2208, n2205, n2209, n2206, n2193, n2202, n2197, 
        n2195, n2196, n2194, n30_adj_4985, n36282, n2291, n34_adj_4986, 
        n32_adj_4987, n33_adj_4988, n31_adj_4989, n2109;
    wire [31:0]n2159;
    
    wire n2126, n2098, n2099, n2097, n2102, n2108, n2107, n2104, 
        n2101, n2105, n2103, n2100, n2106, n2096, n2095, n2094, 
        n2192, n28_adj_4990, n24, n32_adj_4991, n30_adj_4992, n31_adj_4993, 
        n29, n50448, n50449, n50446, n50445, n1999;
    wire [31:0]n2060;
    
    wire n2027, n1997, n1998, n1996, n2003, n2007, n2001, n2002, 
        n2000, n2006, n2004, n2008, n2009, n2005, n1995, n2093, 
        n18, n24_adj_4997, n30_adj_4998, n28_adj_4999, n29_adj_5000, 
        n27_adj_5001;
    wire [31:0]n1;
    
    wire n40603, n50003, n40602, n50001, n40601, n49999, n50391, 
        n50392, n50395, n50394, n1898;
    wire [31:0]n1961;
    
    wire n1928, n1897, n40600, n49997, n1896, n1901, n1909, n1907, 
        n1903, n1900, n1904, n1899, n1905, n1908, n1906, n1902, 
        n36276, n28_adj_5004, n26, n27_adj_5005, n1994, n25_adj_5006;
    wire [3:0]state_3__N_528;
    
    wire n2984, n2885, n41597, n2918;
    wire [31:0]n2951;
    
    wire n2886, n41596, n2887, n41595, n2888, n41594, n2889, n41593, 
        n2890, n41592, n1809;
    wire [31:0]n1862;
    
    wire n1829, n1803, n1802, n2891, n41591, n1801, n41786, n2892, 
        n41590, n1799, n1800, n1798, n1797, n1805, n1804, n1807, 
        n1806, n1808, n2893, n41589, n40599, n49995, n20, n26_adj_5008, 
        n2894, n41588, n1895, n16_adj_5009, n24_adj_5010, n28_adj_5011, 
        n1706;
    wire [31:0]n1763;
    
    wire n1730, n1703, n1707, n1701, n1700, n1699, n1499, n41091, 
        n1433, n1698, n1705, n41785, n1709, n2895, n41587, n1702, 
        n2896, n41586, n2897, n41585, n1704, n1708, n24_adj_5012, 
        n17, n1796, n22_adj_5013, n26_adj_5014, n2898, n41584;
    wire [31:0]n1466;
    
    wire n1401, n41090, n2899, n41583, n40598, n49993, n2900, 
        n41582, n16_adj_5016, n22_adj_5017, n2901, n41581, n1697, 
        n20_adj_5018, n24_adj_5019, n2902, n41580, n2903, n41579, 
        n1631, n53097, n1402, n41089, n2904, n41578, n2905, n41577, 
        n2906, n41576, n2907, n41575, n2908, n41574, n2909, n41573, 
        n40597, n49991, n41784, n1403, n41088, n41783, n41782, 
        n40596, n49989, n41781, n41780, n41779, n1502;
    wire [31:0]n1565;
    
    wire n1532, n1601, n1501, n1600, n1504, n1603, n1500, n1599, 
        n1508, n1607, n1505, n1604, n1406, n41778, n1407, n1506, 
        n1409, n1408, n1507, n1405, n1404, n1503, n41777, n18_adj_5021, 
        n20_adj_5022, n1509, n15, n40595, n49987, n1608, n41087, 
        n1605, n1606, n1609, n1602, n15_adj_5023, n1598, n19, 
        n18_adj_5024, n41776, n22_adj_5025, n41775, n41774, n41773, 
        n40594, n49985, n41772, n41771, n41770, n1235, n53096, 
        n41769, n41763, n40593, n49983, n41086, n41085, n40592, 
        n49981, n41084, n41083, n41082, n1207, n1209, n12_adj_5026, 
        n1205, n1204, n1206, n1208, n13_adj_5027, n1203, n1202, 
        n1136, n53095, n40591, n49979, n1109, n36266, n1106, n1103, 
        n1108, n12_adj_5028, n1107, n1105, n1104, n40590, n49977, 
        n40589, n49975, n41768, n40588, n49973, n40587, n49971, 
        n41767, n41766, n41765, n41764, n40586, n49969, n40585, 
        n49967, n40584, n40583, n40582, n40581, n40580, n40579, 
        n40578, n40577, n40576, n40575, n40574, n40573, n50397, 
        n50398, n50401, n14_adj_5046, n12_adj_5047, n16_adj_5048, 
        n50400, n42233, n42232, n42231, n42230, n42229, n42228, 
        n42227, n42226, n42225, n42224, n42223, n42222, n42221, 
        n42220, n42219, n42218, n42217, n42216, n42215, n42214, 
        n42213, n42212, n40741, n42211, n51824, n42210, n51330, 
        n46577, n51825, n46623, n42209, n42208, \neo_pixel_transmitter.done_N_742 , 
        n42207, n40740, n42206, n42205, n42204, n42203, n42202, 
        n42201, n42200, n42199, n42198, n42197, n42196, n42195, 
        n42194, n42193, n40739, n42192, n42191, n42190, n42189, 
        n42188, n42187, n42186, n42185, n42184, n40738, n42183, 
        n42182, n42181, n42180, n42179, n42178, n42177, n42176, 
        n42175, n42174, n42173, n42172, n42171, n42170, n42169, 
        n42168, n42167, n42166, n42165, n42164, n40737, n42163, 
        n42162, n42161, n42160, n42159, n40736, n42158, n42157, 
        n42156, n42155, n40735, n53209, n53212, n42154, n42153, 
        n42152, n42151;
    wire [31:0]n971;
    
    wire n40557, n1037, n53099, n42150, n42149, n42148, n42147, 
        n42146, n42145, n42144, n40556, n42143, n42142, n36179, 
        n48, n53167, n53170, n42141, n42140, n42139, n2_adj_5049, 
        n52397, n46, n47, n45, n44, n43, n54, n49, n1923, 
        n42138, n40734, n42137, n42136, n42135, n42134, n42133, 
        n29362, n40555, n51314, n42132, n42131, n42130, n42129, 
        n42128, n42127, n40733, n29316, n40554, n42126, n42125, 
        n26353, n40553, n42124, n42123, n42122, n42121, n42120, 
        n42119, n42118, n42117, n42116, n51333, n42115, n42114, 
        n42113, n42112, n40732, n42111, n42110, n42109, n42108, 
        n42107, n42106, n42105, n42104, n42103, n42102, n42101, 
        n42100, n42099, n42098, n42097, n42096, n42095, n42094, 
        n42093, n42092, n42091, n52396, n52398, n1006, n1009, 
        n1008, n42090, n42089, n1007, n52405, n7_adj_5050, n42088, 
        n42087, n40731, n8_adj_5051, n42086, n42085, n42084, n42083, 
        n42082, n42081, n42080, n42079, n42078, n42077, n42076, 
        n42075, n42074, n42073, n42072, n42071, n42070, n42069, 
        n42068, n42067, n42066, n42065, n42064, n42063, n42062, 
        n42061, n42060, n42059, n42058, n42057, n42056, n42055, 
        n42054, n42053, n42052, n42051, n42050, n42049, n42048, 
        n42047, n42046, n42045, n42044, n42043, n42042, n42041, 
        n42040, n42039, n42038, n42037, n42036, n42035, n42034, 
        n42033, n42032, n2786, n42031;
    wire [31:0]n2753;
    
    wire n42030, n42029, n42028, n42027, n42026, n42025, n42024, 
        n42023, n42022, n42021, n42020, n42019, n42018, n42017, 
        n42016, n42015, n42014, n42013, n42012, n42011, n42010, 
        n42009, n2819, n42008, n2787, n42007, n2788, n42006, n2789, 
        n42005, n2790, n42004, n2791, n42003, n2792, n42002, n2793, 
        n42001, n2794, n42000, n2795, n41999, n2796, n41998, n53098, 
        n2797, n41997, n2798, n41996, n2799, n41995, n2800, n41994, 
        n2801, n41993, n2802, n41992, n2803, n41991, n2804, n41990, 
        n2805, n41989, n2806, n41988, n2807, n41987, n2808, n41986, 
        n2809, n41985, n3083, n41984, n3017;
    wire [31:0]n3050;
    
    wire n2985, n41983, n2986, n41982, n2987, n41981, n2988, n41980, 
        n2989, n41979, n2990, n41978, n2991, n41977, n2992, n41976, 
        n2993, n41975, n2994, n41974, n2995, n41973, n2996, n41972, 
        n2997, n41971, n2998, n41970, n2999, n41969, n3000, n41968, 
        n3001, n41967, n3002, n41966, n3003, n41965, n3004, n41964, 
        n3005, n41963, n3006, n41962, n3007, n41961, n3008, n41960, 
        n32309, n41959, n50124, n41958, n3116;
    wire [31:0]n3149;
    
    wire n3084, n41957, n3085, n41956, n3086, n41955, n3087, n41954, 
        n3088, n41953, n3089, n41952, n3090, n41951, n3091, n41950, 
        n3092, n41949, n40547, n3093, n41948, n3094, n41947, n3095, 
        n41946, n40546, n3096, n41945, n3097, n41944, n3098, n41943, 
        n3099, n41942, n3100, n41941, n3101, n41940, n3102, n41939, 
        n3103, n41938, n3104, n41937, n3105, n41936, n3106, n41935, 
        n3107, n41934, n3108, n41933, n40545, n3109, n41932, n40544, 
        n40543, n40542, n48491, n26355, n29324, n12_adj_5052, n16_adj_5053, 
        n17_adj_5054, n32_adj_5055, n42_adj_5056, n38_adj_5057, n43_adj_5058, 
        n40_adj_5059, n46_adj_5060, n39_adj_5061, n47_adj_5062, n44_adj_5063, 
        n33_adj_5064, n40_adj_5065, n45_adj_5066, n42_adj_5067, n48_adj_5068, 
        n41_adj_5069, n49_adj_5070, n36_adj_5071, n46_adj_5072, n42_adj_5073, 
        n34_adj_5074, n43_adj_5075, n50, n48_adj_5076, n49_adj_5077, 
        n47_adj_5078, n29_adj_5079, n11_adj_5080, n19_adj_5081, n27_adj_5082, 
        n23_adj_5083, n15_adj_5084, n49547, n49549, n49543, n49541, 
        n31_adj_5085, n49539, n49551, n49545, n39_adj_5086, n49563, 
        n49561, n3209, n49567, n49569, n49571, n49573, n49575, 
        n49577, n49579, n49581, n49583, n49585, n59, n61, n42492, 
        n48405;
    wire [4:0]color_bit_N_722;
    
    wire n51343, n53110, n52269, n31_adj_5087, n39_adj_5088, n26_adj_5089, 
        n38_adj_5090, n44_adj_5091, n42_adj_5092, n43_adj_5093, n41_adj_5094, 
        n53107;
    
    SB_LUT4 i31206_4_lut (.I0(n27768), .I1(n4), .I2(n42258), .I3(\state[0] ), 
            .O(n46573));
    defparam i31206_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i20_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[1] ), 
            .I2(start), .I3(n46573), .O(n7));
    defparam i20_4_lut.LUT_INIT = 16'hcecf;
    SB_LUT4 i1_4_lut (.I0(n8), .I1(n7), .I2(n46580), .I3(\state[1] ), 
            .O(n44527));
    defparam i1_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 bit_ctr_2058_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[6]), 
            .I3(n41761), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_8 (.CI(n41761), .I0(GND_net), .I1(bit_ctr[6]), 
            .CO(n41762));
    SB_LUT4 bit_ctr_2058_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[5]), 
            .I3(n41760), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_7 (.CI(n41760), .I0(GND_net), .I1(bit_ctr[5]), 
            .CO(n41761));
    SB_LUT4 bit_ctr_2058_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[4]), 
            .I3(n41759), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(CLK_c), .E(n53316), .D(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY bit_ctr_2058_add_4_6 (.CI(n41759), .I0(GND_net), .I1(bit_ctr[4]), 
            .CO(n41760));
    SB_LUT4 bit_ctr_2058_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[3]), 
            .I3(n41758), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFE start_103 (.Q(start), .C(CLK_c), .E(n7_adj_4944), .D(start_N_727));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY bit_ctr_2058_add_4_5 (.CI(n41758), .I0(GND_net), .I1(bit_ctr[3]), 
            .CO(n41759));
    SB_LUT4 bit_ctr_2058_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[2]), 
            .I3(n41757), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_4 (.CI(n41757), .I0(GND_net), .I1(bit_ctr[2]), 
            .CO(n41758));
    SB_LUT4 bit_ctr_2058_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[1]), 
            .I3(n41756), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_3 (.CI(n41756), .I0(GND_net), .I1(bit_ctr[1]), 
            .CO(n41757));
    SB_LUT4 bit_ctr_2058_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_ctr[0]), 
            .CO(n41756));
    SB_LUT4 timer_2057_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n41755), .O(n133_adj_5095[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2057_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n41754), .O(n133_adj_5095[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_32 (.CI(n41754), .I0(GND_net), .I1(timer[30]), 
            .CO(n41755));
    SB_LUT4 mod_5_i1811_3_lut (.I0(n2589), .I1(n2654[30]), .I2(n2621), 
            .I3(GND_net), .O(n2688));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1826_3_lut (.I0(n2604), .I1(n2654[15]), .I2(n2621), 
            .I3(GND_net), .O(n2703));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1822_3_lut (.I0(n2600), .I1(n2654[19]), .I2(n2621), 
            .I3(GND_net), .O(n2699));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2057_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n41753), .O(n133_adj_5095[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1827_3_lut (.I0(n2605), .I1(n2654[14]), .I2(n2621), 
            .I3(GND_net), .O(n2704));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1824_3_lut (.I0(n2602), .I1(n2654[17]), .I2(n2621), 
            .I3(GND_net), .O(n2701));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1829_3_lut (.I0(n2607), .I1(n2654[12]), .I2(n2621), 
            .I3(GND_net), .O(n2706));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1828_3_lut (.I0(n2606), .I1(n2654[13]), .I2(n2621), 
            .I3(GND_net), .O(n2705));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1820_3_lut (.I0(n2598), .I1(n2654[21]), .I2(n2621), 
            .I3(GND_net), .O(n2697));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1823_3_lut (.I0(n2601), .I1(n2654[18]), .I2(n2621), 
            .I3(GND_net), .O(n2700));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1831_3_lut (.I0(n2609), .I1(n2654[10]), .I2(n2621), 
            .I3(GND_net), .O(n2708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1825_3_lut (.I0(n2603), .I1(n2654[16]), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1830_3_lut (.I0(n2608), .I1(n2654[11]), .I2(n2621), 
            .I3(GND_net), .O(n2707));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1819_3_lut (.I0(n2597), .I1(n2654[22]), .I2(n2621), 
            .I3(GND_net), .O(n2696));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1817_3_lut (.I0(n2595), .I1(n2654[24]), .I2(n2621), 
            .I3(GND_net), .O(n2694));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1818_3_lut (.I0(n2596), .I1(n2654[23]), .I2(n2621), 
            .I3(GND_net), .O(n2695));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1816_3_lut (.I0(n2594), .I1(n2654[25]), .I2(n2621), 
            .I3(GND_net), .O(n2693));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1815_3_lut (.I0(n2593), .I1(n2654[26]), .I2(n2621), 
            .I3(GND_net), .O(n2692));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1813_3_lut (.I0(n2591), .I1(n2654[28]), .I2(n2621), 
            .I3(GND_net), .O(n2690));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1814_3_lut (.I0(n2592), .I1(n2654[27]), .I2(n2621), 
            .I3(GND_net), .O(n2691));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1812_3_lut (.I0(n2590), .I1(n2654[29]), .I2(n2621), 
            .I3(GND_net), .O(n2689));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1832_3_lut (.I0(bit_ctr[9]), .I1(n2654[9]), .I2(n2621), 
            .I3(GND_net), .O(n2709));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1821_3_lut (.I0(n2599), .I1(n2654[20]), .I2(n2621), 
            .I3(GND_net), .O(n2698));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_3_lut (.I0(bit_ctr[8]), .I1(n2698), .I2(n2709), .I3(GND_net), 
            .O(n30));
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY timer_2057_add_4_31 (.CI(n41753), .I0(GND_net), .I1(timer[29]), 
            .CO(n41754));
    SB_LUT4 timer_2057_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n41752), .O(n133_adj_5095[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_30 (.CI(n41752), .I0(GND_net), .I1(timer[28]), 
            .CO(n41753));
    SB_LUT4 timer_2057_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n41751), .O(n133_adj_5095[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_29 (.CI(n41751), .I0(GND_net), .I1(timer[27]), 
            .CO(n41752));
    SB_LUT4 timer_2057_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n41750), .O(n133_adj_5095[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_28 (.CI(n41750), .I0(GND_net), .I1(timer[26]), 
            .CO(n41751));
    SB_LUT4 timer_2057_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n41749), .O(n133_adj_5095[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_27 (.CI(n41749), .I0(GND_net), .I1(timer[25]), 
            .CO(n41750));
    SB_LUT4 timer_2057_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n41748), .O(n133_adj_5095[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut (.I0(n2693), .I1(n2695), .I2(n2694), .I3(n2696), 
            .O(n37));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2689), .I1(n2691), .I2(n2690), .I3(n2692), 
            .O(n36));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n2697), .I2(n30), .I3(n2705), .O(n42));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_2057_add_4_26 (.CI(n41748), .I0(GND_net), .I1(timer[24]), 
            .CO(n41749));
    SB_LUT4 timer_2057_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n41747), .O(n133_adj_5095[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_25 (.CI(n41747), .I0(GND_net), .I1(timer[23]), 
            .CO(n41748));
    SB_LUT4 timer_2057_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n41746), .O(n133_adj_5095[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_24 (.CI(n41746), .I0(GND_net), .I1(timer[22]), 
            .CO(n41747));
    SB_LUT4 timer_2057_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n41745), .O(n133_adj_5095[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_23 (.CI(n41745), .I0(GND_net), .I1(timer[21]), 
            .CO(n41746));
    SB_LUT4 timer_2057_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n41744), .O(n133_adj_5095[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_22 (.CI(n41744), .I0(GND_net), .I1(timer[20]), 
            .CO(n41745));
    SB_LUT4 timer_2057_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n41743), .O(n133_adj_5095[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_21 (.CI(n41743), .I0(GND_net), .I1(timer[19]), 
            .CO(n41744));
    SB_LUT4 timer_2057_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n41742), .O(n133_adj_5095[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut (.I0(n2707), .I1(n2702), .I2(n2708), .I3(n2700), 
            .O(n40));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n2703), .I1(n36), .I2(n2688), .I3(n2687), 
            .O(n41));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_2057_add_4_20 (.CI(n41742), .I0(GND_net), .I1(timer[18]), 
            .CO(n41743));
    SB_LUT4 timer_2057_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n41741), .O(n133_adj_5095[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_19 (.CI(n41741), .I0(GND_net), .I1(timer[17]), 
            .CO(n41742));
    SB_LUT4 timer_2057_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n41740), .O(n133_adj_5095[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_18 (.CI(n41740), .I0(GND_net), .I1(timer[16]), 
            .CO(n41741));
    SB_LUT4 timer_2057_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n41739), .O(n133_adj_5095[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_17 (.CI(n41739), .I0(GND_net), .I1(timer[15]), 
            .CO(n41740));
    SB_LUT4 timer_2057_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n41738), .O(n133_adj_5095[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_16 (.CI(n41738), .I0(GND_net), .I1(timer[14]), 
            .CO(n41739));
    SB_LUT4 i16_4_lut (.I0(n2706), .I1(n2701), .I2(n2704), .I3(n2699), 
            .O(n39));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_2057_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n41737), .O(n133_adj_5095[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n6801), 
            .I3(GND_net), .O(n6));   // verilog/neopixel.v(36[4] 116[11])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i15855_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n29252), 
            .I3(GND_net), .O(n29377));   // verilog/neopixel.v(36[4] 116[11])
    defparam i15855_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_DFFESR bit_ctr_2058__i31 (.Q(bit_ctr[31]), .C(CLK_c), .E(n6801), 
            .D(n133[31]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i30 (.Q(bit_ctr[30]), .C(CLK_c), .E(n6801), 
            .D(n133[30]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i29 (.Q(bit_ctr[29]), .C(CLK_c), .E(n6801), 
            .D(n133[29]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i28 (.Q(bit_ctr[28]), .C(CLK_c), .E(n6801), 
            .D(n133[28]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i27 (.Q(bit_ctr[27]), .C(CLK_c), .E(n6801), 
            .D(n133[27]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i26 (.Q(bit_ctr[26]), .C(CLK_c), .E(n6801), 
            .D(n133[26]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i25 (.Q(bit_ctr[25]), .C(CLK_c), .E(n6801), 
            .D(n133[25]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i24 (.Q(bit_ctr[24]), .C(CLK_c), .E(n6801), 
            .D(n133[24]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i23 (.Q(bit_ctr[23]), .C(CLK_c), .E(n6801), 
            .D(n133[23]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i22 (.Q(bit_ctr[22]), .C(CLK_c), .E(n6801), 
            .D(n133[22]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i0 (.Q(bit_ctr[0]), .C(CLK_c), .E(n6801), 
            .D(n133[0]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i21 (.Q(bit_ctr[21]), .C(CLK_c), .E(n6801), 
            .D(n133[21]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_CARRY timer_2057_add_4_15 (.CI(n41737), .I0(GND_net), .I1(timer[13]), 
            .CO(n41738));
    SB_DFFESR bit_ctr_2058__i20 (.Q(bit_ctr[20]), .C(CLK_c), .E(n6801), 
            .D(n133[20]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i19 (.Q(bit_ctr[19]), .C(CLK_c), .E(n6801), 
            .D(n133[19]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i18 (.Q(bit_ctr[18]), .C(CLK_c), .E(n6801), 
            .D(n133[18]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i17 (.Q(bit_ctr[17]), .C(CLK_c), .E(n6801), 
            .D(n133[17]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 timer_2057_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n41736), .O(n133_adj_5095[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_14 (.CI(n41736), .I0(GND_net), .I1(timer[12]), 
            .CO(n41737));
    SB_LUT4 mod_5_i1753_3_lut (.I0(n2499), .I1(n2555[21]), .I2(n2522), 
            .I3(GND_net), .O(n2598));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1763_3_lut (.I0(n2509), .I1(n2555[11]), .I2(n2522), 
            .I3(GND_net), .O(n2608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1756_3_lut (.I0(n2502), .I1(n2555[18]), .I2(n2522), 
            .I3(GND_net), .O(n2601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1761_3_lut (.I0(n2507), .I1(n2555[13]), .I2(n2522), 
            .I3(GND_net), .O(n2606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1752_3_lut (.I0(n2498), .I1(n2555[22]), .I2(n2522), 
            .I3(GND_net), .O(n2597));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1762_3_lut (.I0(n2508), .I1(n2555[12]), .I2(n2522), 
            .I3(GND_net), .O(n2607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1759_3_lut (.I0(n2505), .I1(n2555[15]), .I2(n2522), 
            .I3(GND_net), .O(n2604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1750_3_lut (.I0(n2496), .I1(n2555[24]), .I2(n2522), 
            .I3(GND_net), .O(n2595));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1758_3_lut (.I0(n2504), .I1(n2555[16]), .I2(n2522), 
            .I3(GND_net), .O(n2603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1754_3_lut (.I0(n2500), .I1(n2555[20]), .I2(n2522), 
            .I3(GND_net), .O(n2599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1755_3_lut (.I0(n2501), .I1(n2555[19]), .I2(n2522), 
            .I3(GND_net), .O(n2600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1757_3_lut (.I0(n2503), .I1(n2555[17]), .I2(n2522), 
            .I3(GND_net), .O(n2602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1760_3_lut (.I0(n2506), .I1(n2555[14]), .I2(n2522), 
            .I3(GND_net), .O(n2605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1748_3_lut (.I0(n2494), .I1(n2555[26]), .I2(n2522), 
            .I3(GND_net), .O(n2593));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1749_3_lut (.I0(n2495), .I1(n2555[25]), .I2(n2522), 
            .I3(GND_net), .O(n2594));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1747_3_lut (.I0(n2493), .I1(n2555[27]), .I2(n2522), 
            .I3(GND_net), .O(n2592));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1746_3_lut (.I0(n2492), .I1(n2555[28]), .I2(n2522), 
            .I3(GND_net), .O(n2591));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1745_3_lut (.I0(n2491), .I1(n2555[29]), .I2(n2522), 
            .I3(GND_net), .O(n2590));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1744_3_lut (.I0(n2490), .I1(n2555[30]), .I2(n2522), 
            .I3(GND_net), .O(n2589));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1764_3_lut (.I0(bit_ctr[10]), .I1(n2555[10]), .I2(n2522), 
            .I3(GND_net), .O(n2609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1751_3_lut (.I0(n2497), .I1(n2555[23]), .I2(n2522), 
            .I3(GND_net), .O(n2596));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut (.I0(bit_ctr[9]), .I1(n2596), .I2(n2609), .I3(GND_net), 
            .O(n28));
    defparam i6_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1526 (.I0(n2592), .I1(n2594), .I2(n2593), .I3(n2605), 
            .O(n35));
    defparam i13_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2589), .I1(n2590), .I2(n2588), .I3(n2591), 
            .O(n34));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1527 (.I0(n35), .I1(n2595), .I2(n28), .I3(n2604), 
            .O(n40_adj_4960));
    defparam i18_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1528 (.I0(n2602), .I1(n2600), .I2(n2599), .I3(n2603), 
            .O(n38));
    defparam i16_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2608), .I1(n34), .I2(n2598), .I3(GND_net), 
            .O(n39_adj_4961));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut (.I0(n2607), .I1(n2597), .I2(n2606), .I3(n2601), 
            .O(n37_adj_4962));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n37_adj_4962), .I1(n39_adj_4961), .I2(n38), 
            .I3(n40_adj_4960), .O(n2621));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_2057_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n41735), .O(n133_adj_5095[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_13 (.CI(n41735), .I0(GND_net), .I1(timer[11]), 
            .CO(n41736));
    SB_LUT4 timer_2057_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n41734), .O(n133_adj_5095[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1693_3_lut (.I0(n2407), .I1(n2456[14]), .I2(n2423), 
            .I3(GND_net), .O(n2506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1693_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2057_add_4_12 (.CI(n41734), .I0(GND_net), .I1(timer[10]), 
            .CO(n41735));
    SB_LUT4 mod_5_i1695_3_lut (.I0(n2409), .I1(n2456[12]), .I2(n2423), 
            .I3(GND_net), .O(n2508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1692_3_lut (.I0(n2406), .I1(n2456[15]), .I2(n2423), 
            .I3(GND_net), .O(n2505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2057_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n41733), .O(n133_adj_5095[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1690_3_lut (.I0(n2404), .I1(n2456[17]), .I2(n2423), 
            .I3(GND_net), .O(n2503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1686_3_lut (.I0(n2400), .I1(n2456[21]), .I2(n2423), 
            .I3(GND_net), .O(n2499));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1685_3_lut (.I0(n2399), .I1(n2456[22]), .I2(n2423), 
            .I3(GND_net), .O(n2498));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1683_3_lut (.I0(n2397), .I1(n2456[24]), .I2(n2423), 
            .I3(GND_net), .O(n2496));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1684_3_lut (.I0(n2398), .I1(n2456[23]), .I2(n2423), 
            .I3(GND_net), .O(n2497));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1682_3_lut (.I0(n2396), .I1(n2456[25]), .I2(n2423), 
            .I3(GND_net), .O(n2495));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1681_3_lut (.I0(n2395), .I1(n2456[26]), .I2(n2423), 
            .I3(GND_net), .O(n2494));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1679_3_lut (.I0(n2393), .I1(n2456[28]), .I2(n2423), 
            .I3(GND_net), .O(n2492));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1680_3_lut (.I0(n2394), .I1(n2456[27]), .I2(n2423), 
            .I3(GND_net), .O(n2493));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1678_3_lut (.I0(n2392), .I1(n2456[29]), .I2(n2423), 
            .I3(GND_net), .O(n2491));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1691_3_lut (.I0(n2405), .I1(n2456[16]), .I2(n2423), 
            .I3(GND_net), .O(n2504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1689_3_lut (.I0(n2403), .I1(n2456[18]), .I2(n2423), 
            .I3(GND_net), .O(n2502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1687_3_lut (.I0(n2401), .I1(n2456[20]), .I2(n2423), 
            .I3(GND_net), .O(n2500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1694_3_lut (.I0(n2408), .I1(n2456[13]), .I2(n2423), 
            .I3(GND_net), .O(n2507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1694_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2057_add_4_11 (.CI(n41733), .I0(GND_net), .I1(timer[9]), 
            .CO(n41734));
    SB_LUT4 timer_2057_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n41732), .O(n133_adj_5095[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1696_3_lut (.I0(bit_ctr[11]), .I1(n2456[11]), .I2(n2423), 
            .I3(GND_net), .O(n2509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1696_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2057_add_4_10 (.CI(n41732), .I0(GND_net), .I1(timer[8]), 
            .CO(n41733));
    SB_LUT4 mod_5_i1688_3_lut (.I0(n2402), .I1(n2456[19]), .I2(n2423), 
            .I3(GND_net), .O(n2501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1677_3_lut (.I0(n2391), .I1(n2456[30]), .I2(n2423), 
            .I3(GND_net), .O(n2490));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n2490), .I1(n2489), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1529 (.I0(n2507), .I1(n2500), .I2(n2502), .I3(n2504), 
            .O(n36_adj_4963));
    defparam i15_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_3_lut_adj_1530 (.I0(n2501), .I1(bit_ctr[10]), .I2(n2509), 
            .I3(GND_net), .O(n27));
    defparam i6_3_lut_adj_1530.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1531 (.I0(n2495), .I1(n2497), .I2(n2496), .I3(n2498), 
            .O(n34_adj_4964));
    defparam i13_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1532 (.I0(n2491), .I1(n2493), .I2(n2492), .I3(n2494), 
            .O(n33));
    defparam i12_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1533 (.I0(n2505), .I1(n2508), .I2(n2506), .I3(n22), 
            .O(n37_adj_4965));
    defparam i16_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1534 (.I0(n27), .I1(n36_adj_4963), .I2(n2499), 
            .I3(n2503), .O(n39_adj_4966));
    defparam i18_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1535 (.I0(n39_adj_4966), .I1(n37_adj_4965), .I2(n33), 
            .I3(n34_adj_4964), .O(n2522));
    defparam i20_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_2057_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n41731), .O(n133_adj_5095[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_9 (.CI(n41731), .I0(GND_net), .I1(timer[7]), 
            .CO(n41732));
    SB_LUT4 timer_2057_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n41730), .O(n133_adj_5095[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_8 (.CI(n41730), .I0(GND_net), .I1(timer[6]), 
            .CO(n41731));
    SB_LUT4 timer_2057_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n41729), .O(n133_adj_5095[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_7 (.CI(n41729), .I0(GND_net), .I1(timer[5]), 
            .CO(n41730));
    SB_LUT4 timer_2057_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n41728), .O(n133_adj_5095[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_6 (.CI(n41728), .I0(GND_net), .I1(timer[4]), 
            .CO(n41729));
    SB_LUT4 timer_2057_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n41727), .O(n133_adj_5095[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_5 (.CI(n41727), .I0(GND_net), .I1(timer[3]), 
            .CO(n41728));
    SB_LUT4 timer_2057_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n41726), .O(n133_adj_5095[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_4 (.CI(n41726), .I0(GND_net), .I1(timer[2]), 
            .CO(n41727));
    SB_LUT4 timer_2057_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n41725), .O(n133_adj_5095[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_3 (.CI(n41725), .I0(GND_net), .I1(timer[1]), 
            .CO(n41726));
    SB_LUT4 timer_2057_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133_adj_5095[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n41725));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1334), .I1(n1301), .I2(VCC_net), 
            .I3(n41717), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'h8228;
    SB_DFFESR bit_ctr_2058__i16 (.Q(bit_ctr[16]), .C(CLK_c), .E(n6801), 
            .D(n133[16]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_add_937_10_lut (.I0(GND_net), .I1(n1302), .I2(VCC_net), 
            .I3(n41716), .O(n1367[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_10 (.CI(n41716), .I0(n1302), .I1(VCC_net), 
            .CO(n41717));
    SB_LUT4 mod_5_add_937_9_lut (.I0(GND_net), .I1(n1303), .I2(VCC_net), 
            .I3(n41715), .O(n1367[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_9 (.CI(n41715), .I0(n1303), .I1(VCC_net), .CO(n41716));
    SB_DFFESR bit_ctr_2058__i15 (.Q(bit_ctr[15]), .C(CLK_c), .E(n6801), 
            .D(n133[15]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_add_937_8_lut (.I0(GND_net), .I1(n1304), .I2(VCC_net), 
            .I3(n41714), .O(n1367[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_8 (.CI(n41714), .I0(n1304), .I1(VCC_net), .CO(n41715));
    SB_LUT4 i22912_4_lut (.I0(one_wire_N_679[8]), .I1(n27952), .I2(one_wire_N_679[10]), 
            .I3(one_wire_N_679[9]), .O(n36444));
    defparam i22912_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1536 (.I0(one_wire_N_679[2]), .I1(one_wire_N_679[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4));
    defparam i1_2_lut_adj_1536.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_937_7_lut (.I0(GND_net), .I1(n1305), .I2(VCC_net), 
            .I3(n41713), .O(n1367[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_7 (.CI(n41713), .I0(n1305), .I1(VCC_net), .CO(n41714));
    SB_LUT4 mod_5_add_937_6_lut (.I0(GND_net), .I1(n1306), .I2(VCC_net), 
            .I3(n41712), .O(n1367[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_6 (.CI(n41712), .I0(n1306), .I1(VCC_net), .CO(n41713));
    SB_LUT4 mod_5_add_937_5_lut (.I0(GND_net), .I1(n1307), .I2(VCC_net), 
            .I3(n41711), .O(n1367[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_5 (.CI(n41711), .I0(n1307), .I1(VCC_net), .CO(n41712));
    SB_LUT4 mod_5_add_937_4_lut (.I0(GND_net), .I1(n1308), .I2(VCC_net), 
            .I3(n41710), .O(n1367[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_4 (.CI(n41710), .I0(n1308), .I1(VCC_net), .CO(n41711));
    SB_LUT4 i2_2_lut (.I0(one_wire_N_679[2]), .I1(n4_adj_4976), .I2(GND_net), 
            .I3(GND_net), .O(n42258));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_937_3_lut (.I0(GND_net), .I1(n1309), .I2(GND_net), 
            .I3(n41709), .O(n1367[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_2058__i14 (.Q(bit_ctr[14]), .C(CLK_c), .E(n6801), 
            .D(n133[14]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_CARRY mod_5_add_937_3 (.CI(n41709), .I0(n1309), .I1(GND_net), .CO(n41710));
    SB_LUT4 i1_2_lut_adj_1537 (.I0(one_wire_N_679[5]), .I1(one_wire_N_679[4]), 
            .I2(GND_net), .I3(GND_net), .O(n50005));   // verilog/neopixel.v(104[14:39])
    defparam i1_2_lut_adj_1537.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1538 (.I0(one_wire_N_679[8]), .I1(one_wire_N_679[7]), 
            .I2(one_wire_N_679[6]), .I3(n50005), .O(n50011));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_2_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(VCC_net), .O(n1367[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(GND_net), 
            .CO(n41709));
    SB_LUT4 i1_4_lut_adj_1539 (.I0(one_wire_N_679[10]), .I1(n27952), .I2(one_wire_N_679[9]), 
            .I3(n50011), .O(n27768));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i31210_4_lut (.I0(n27768), .I1(n42258), .I2(n4), .I3(\state[0] ), 
            .O(n46580));
    defparam i31210_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i35979_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n51335));
    defparam i35979_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR bit_ctr_2058__i13 (.Q(bit_ctr[13]), .C(CLK_c), .E(n6801), 
            .D(n133[13]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i12 (.Q(bit_ctr[12]), .C(CLK_c), .E(n6801), 
            .D(n133[12]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i11 (.Q(bit_ctr[11]), .C(CLK_c), .E(n6801), 
            .D(n133[11]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 i31211_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n46580), .I3(GND_net), .O(n46581));
    defparam i31211_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_i1625_3_lut (.I0(n2307), .I1(n2357[15]), .I2(n2324), 
            .I3(GND_net), .O(n2406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1616_3_lut (.I0(n2298), .I1(n2357[24]), .I2(n2324), 
            .I3(GND_net), .O(n2397));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1620_3_lut (.I0(n2302), .I1(n2357[20]), .I2(n2324), 
            .I3(GND_net), .O(n2401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1621_3_lut (.I0(n2303), .I1(n2357[19]), .I2(n2324), 
            .I3(GND_net), .O(n2402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1626_3_lut (.I0(n2308), .I1(n2357[14]), .I2(n2324), 
            .I3(GND_net), .O(n2407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1618_3_lut (.I0(n2300), .I1(n2357[22]), .I2(n2324), 
            .I3(GND_net), .O(n2399));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1612_3_lut (.I0(n2294), .I1(n2357[28]), .I2(n2324), 
            .I3(GND_net), .O(n2393));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1611_3_lut (.I0(n2293), .I1(n2357[29]), .I2(n2324), 
            .I3(GND_net), .O(n2392));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1610_3_lut (.I0(n2292), .I1(n2357[30]), .I2(n2324), 
            .I3(GND_net), .O(n2391));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1615_3_lut (.I0(n2297), .I1(n2357[25]), .I2(n2324), 
            .I3(GND_net), .O(n2396));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15_4_lut_adj_1540 (.I0(n46581), .I1(n51335), .I2(\state[1] ), 
            .I3(n36444), .O(n7_adj_4944));
    defparam i15_4_lut_adj_1540.LUT_INIT = 16'h3a0a;
    SB_LUT4 mod_5_i1614_3_lut (.I0(n2296), .I1(n2357[26]), .I2(n2324), 
            .I3(GND_net), .O(n2395));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36905_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(start_N_727));   // verilog/neopixel.v(36[4] 116[11])
    defparam i36905_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 mod_5_i1619_3_lut (.I0(n2301), .I1(n2357[21]), .I2(n2324), 
            .I3(GND_net), .O(n2400));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1613_3_lut (.I0(n2295), .I1(n2357[27]), .I2(n2324), 
            .I3(GND_net), .O(n2394));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1628_3_lut (.I0(bit_ctr[12]), .I1(n2357[12]), .I2(n2324), 
            .I3(GND_net), .O(n2409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1617_3_lut (.I0(n2299), .I1(n2357[23]), .I2(n2324), 
            .I3(GND_net), .O(n2398));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1624_3_lut (.I0(n2306), .I1(n2357[16]), .I2(n2324), 
            .I3(GND_net), .O(n2405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1627_3_lut (.I0(n2309), .I1(n2357[13]), .I2(n2324), 
            .I3(GND_net), .O(n2408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31108_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n46472));
    defparam i31108_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i36846_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n45634));
    defparam i36846_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1541 (.I0(one_wire_N_679[2]), .I1(n45634), .I2(one_wire_N_679[3]), 
            .I3(n4_adj_4976), .O(n103));
    defparam i1_4_lut_adj_1541.LUT_INIT = 16'h45cd;
    SB_LUT4 mod_5_i1623_3_lut (.I0(n2305), .I1(n2357[17]), .I2(n2324), 
            .I3(GND_net), .O(n2404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1622_3_lut (.I0(n2304), .I1(n2357[18]), .I2(n2324), 
            .I3(GND_net), .O(n2403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut_adj_1542 (.I0(n2403), .I1(n2404), .I2(n2408), .I3(n2405), 
            .O(n34_adj_4981));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(n2398), .I1(bit_ctr[11]), .I2(n2409), .I3(GND_net), 
            .O(n25));   // verilog/neopixel.v(22[26:36])
    defparam i5_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1543 (.I0(n2394), .I1(n2400), .I2(n2395), .I3(n2396), 
            .O(n32));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2391), .I1(n2392), .I2(n2390), .I3(n2393), 
            .O(n31));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1544 (.I0(n2399), .I1(n2407), .I2(n2402), .I3(n2401), 
            .O(n35_adj_4982));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1545 (.I0(n25), .I1(n34_adj_4981), .I2(n2397), 
            .I3(n2406), .O(n37_adj_4983));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_679[7]), .I1(one_wire_N_679[9]), .I2(n46472), 
            .I3(n103), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i19_4_lut_adj_1546 (.I0(n37_adj_4983), .I1(n35_adj_4982), .I2(n31), 
            .I3(n32), .O(n2423));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1551_3_lut (.I0(n2201), .I1(n2258[22]), .I2(n2225), 
            .I3(GND_net), .O(n2300));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1547 (.I0(one_wire_N_679[8]), .I1(one_wire_N_679[4]), 
            .I2(n16), .I3(n27952), .O(n6_adj_4984));
    defparam i1_4_lut_adj_1547.LUT_INIT = 16'hffef;
    SB_LUT4 mod_5_i1549_3_lut (.I0(n2199), .I1(n2258[24]), .I2(n2225), 
            .I3(GND_net), .O(n2298));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1550_3_lut (.I0(n2200), .I1(n2258[23]), .I2(n2225), 
            .I3(GND_net), .O(n2299));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1548_3_lut (.I0(n2198), .I1(n2258[25]), .I2(n2225), 
            .I3(GND_net), .O(n2297));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut (.I0(one_wire_N_679[10]), .I1(one_wire_N_679[6]), .I2(one_wire_N_679[5]), 
            .I3(n6_adj_4984), .O(n53316));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1554_3_lut (.I0(n2204), .I1(n2258[19]), .I2(n2225), 
            .I3(GND_net), .O(n2303));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1557_3_lut (.I0(n2207), .I1(n2258[16]), .I2(n2225), 
            .I3(GND_net), .O(n2306));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1553_3_lut (.I0(n2203), .I1(n2258[20]), .I2(n2225), 
            .I3(GND_net), .O(n2302));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1558_3_lut (.I0(n2208), .I1(n2258[15]), .I2(n2225), 
            .I3(GND_net), .O(n2307));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1555_3_lut (.I0(n2205), .I1(n2258[18]), .I2(n2225), 
            .I3(GND_net), .O(n2304));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1559_3_lut (.I0(n2209), .I1(n2258[14]), .I2(n2225), 
            .I3(GND_net), .O(n2308));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1556_3_lut (.I0(n2206), .I1(n2258[17]), .I2(n2225), 
            .I3(GND_net), .O(n2305));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1543_3_lut (.I0(n2193), .I1(n2258[30]), .I2(n2225), 
            .I3(GND_net), .O(n2292));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1552_3_lut (.I0(n2202), .I1(n2258[21]), .I2(n2225), 
            .I3(GND_net), .O(n2301));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1547_3_lut (.I0(n2197), .I1(n2258[26]), .I2(n2225), 
            .I3(GND_net), .O(n2296));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1239_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_1239_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 mod_5_i1545_3_lut (.I0(n2195), .I1(n2258[28]), .I2(n2225), 
            .I3(GND_net), .O(n2294));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1546_3_lut (.I0(n2196), .I1(n2258[27]), .I2(n2225), 
            .I3(GND_net), .O(n2295));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1544_3_lut (.I0(n2194), .I1(n2258[29]), .I2(n2225), 
            .I3(GND_net), .O(n2293));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1560_3_lut (.I0(bit_ctr[13]), .I1(n2258[13]), .I2(n2225), 
            .I3(GND_net), .O(n2309));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1548 (.I0(n2293), .I1(n2295), .I2(n2294), .I3(n2296), 
            .O(n30_adj_4985));
    defparam i11_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i22754_2_lut (.I0(bit_ctr[12]), .I1(n2309), .I2(GND_net), 
            .I3(GND_net), .O(n36282));
    defparam i22754_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15_4_lut_adj_1549 (.I0(n2301), .I1(n30_adj_4985), .I2(n2292), 
            .I3(n2291), .O(n34_adj_4986));
    defparam i15_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1550 (.I0(n2305), .I1(n2308), .I2(n36282), .I3(n2304), 
            .O(n32_adj_4987));
    defparam i13_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1551 (.I0(n2307), .I1(n2302), .I2(n2306), .I3(n2303), 
            .O(n33_adj_4988));
    defparam i14_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1552 (.I0(n2297), .I1(n2299), .I2(n2298), .I3(n2300), 
            .O(n31_adj_4989));
    defparam i12_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1553 (.I0(n31_adj_4989), .I1(n33_adj_4988), .I2(n32_adj_4987), 
            .I3(n34_adj_4986), .O(n2324));
    defparam i18_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1491_3_lut (.I0(n2109), .I1(n2159[15]), .I2(n2126), 
            .I3(GND_net), .O(n2208));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1480_3_lut (.I0(n2098), .I1(n2159[26]), .I2(n2126), 
            .I3(GND_net), .O(n2197));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1481_3_lut (.I0(n2099), .I1(n2159[25]), .I2(n2126), 
            .I3(GND_net), .O(n2198));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1479_3_lut (.I0(n2097), .I1(n2159[27]), .I2(n2126), 
            .I3(GND_net), .O(n2196));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1484_3_lut (.I0(n2102), .I1(n2159[22]), .I2(n2126), 
            .I3(GND_net), .O(n2201));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1490_3_lut (.I0(n2108), .I1(n2159[16]), .I2(n2126), 
            .I3(GND_net), .O(n2207));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1489_3_lut (.I0(n2107), .I1(n2159[17]), .I2(n2126), 
            .I3(GND_net), .O(n2206));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1486_3_lut (.I0(n2104), .I1(n2159[20]), .I2(n2126), 
            .I3(GND_net), .O(n2203));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1492_3_lut (.I0(bit_ctr[14]), .I1(n2159[14]), .I2(n2126), 
            .I3(GND_net), .O(n2209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1483_3_lut (.I0(n2101), .I1(n2159[23]), .I2(n2126), 
            .I3(GND_net), .O(n2200));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1487_3_lut (.I0(n2105), .I1(n2159[19]), .I2(n2126), 
            .I3(GND_net), .O(n2204));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1485_3_lut (.I0(n2103), .I1(n2159[21]), .I2(n2126), 
            .I3(GND_net), .O(n2202));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1482_3_lut (.I0(n2100), .I1(n2159[24]), .I2(n2126), 
            .I3(GND_net), .O(n2199));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1488_3_lut (.I0(n2106), .I1(n2159[18]), .I2(n2126), 
            .I3(GND_net), .O(n2205));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1478_3_lut (.I0(n2096), .I1(n2159[28]), .I2(n2126), 
            .I3(GND_net), .O(n2195));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1477_3_lut (.I0(n2095), .I1(n2159[29]), .I2(n2126), 
            .I3(GND_net), .O(n2194));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1476_3_lut (.I0(n2094), .I1(n2159[30]), .I2(n2126), 
            .I3(GND_net), .O(n2193));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut (.I0(n2193), .I1(n2194), .I2(n2192), .I3(n2195), 
            .O(n28_adj_4990));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n2205), .I1(n2199), .I2(GND_net), .I3(GND_net), 
            .O(n24));   // verilog/neopixel.v(22[26:36])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14_3_lut (.I0(n2202), .I1(n28_adj_4990), .I2(n2204), .I3(GND_net), 
            .O(n32_adj_4991));   // verilog/neopixel.v(22[26:36])
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut_adj_1554 (.I0(bit_ctr[13]), .I1(n24), .I2(n2200), 
            .I3(n2209), .O(n30_adj_4992));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1554.LUT_INIT = 16'hfefc;
    SB_LUT4 i13_4_lut_adj_1555 (.I0(n2203), .I1(n2206), .I2(n2207), .I3(n2201), 
            .O(n31_adj_4993));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1556 (.I0(n2196), .I1(n2198), .I2(n2197), .I3(n2208), 
            .O(n29));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1557 (.I0(n29), .I1(n31_adj_4993), .I2(n30_adj_4992), 
            .I3(n32_adj_4991), .O(n2225));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i34966_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50448));
    defparam i34966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34967_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50449));
    defparam i34967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34964_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50446));
    defparam i34964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34963_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50445));
    defparam i34963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1413_3_lut (.I0(n1999), .I1(n2060[26]), .I2(n2027), 
            .I3(GND_net), .O(n2098));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1411_3_lut (.I0(n1997), .I1(n2060[28]), .I2(n2027), 
            .I3(GND_net), .O(n2096));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1412_3_lut (.I0(n1998), .I1(n2060[27]), .I2(n2027), 
            .I3(GND_net), .O(n2097));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1410_3_lut (.I0(n1996), .I1(n2060[29]), .I2(n2027), 
            .I3(GND_net), .O(n2095));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1424_3_lut (.I0(bit_ctr[15]), .I1(n2060[15]), .I2(n2027), 
            .I3(GND_net), .O(n2109));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1417_3_lut (.I0(n2003), .I1(n2060[22]), .I2(n2027), 
            .I3(GND_net), .O(n2102));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1421_3_lut (.I0(n2007), .I1(n2060[18]), .I2(n2027), 
            .I3(GND_net), .O(n2106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1415_3_lut (.I0(n2001), .I1(n2060[24]), .I2(n2027), 
            .I3(GND_net), .O(n2100));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1416_3_lut (.I0(n2002), .I1(n2060[23]), .I2(n2027), 
            .I3(GND_net), .O(n2101));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR bit_ctr_2058__i10 (.Q(bit_ctr[10]), .C(CLK_c), .E(n6801), 
            .D(n133[10]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_i1414_3_lut (.I0(n2000), .I1(n2060[25]), .I2(n2027), 
            .I3(GND_net), .O(n2099));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR bit_ctr_2058__i9 (.Q(bit_ctr[9]), .C(CLK_c), .E(n6801), 
            .D(n133[9]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i8 (.Q(bit_ctr[8]), .C(CLK_c), .E(n6801), 
            .D(n133[8]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_i1420_3_lut (.I0(n2006), .I1(n2060[19]), .I2(n2027), 
            .I3(GND_net), .O(n2105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1418_3_lut (.I0(n2004), .I1(n2060[21]), .I2(n2027), 
            .I3(GND_net), .O(n2103));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1422_3_lut (.I0(n2008), .I1(n2060[17]), .I2(n2027), 
            .I3(GND_net), .O(n2107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1423_3_lut (.I0(n2009), .I1(n2060[16]), .I2(n2027), 
            .I3(GND_net), .O(n2108));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1419_3_lut (.I0(n2005), .I1(n2060[20]), .I2(n2027), 
            .I3(GND_net), .O(n2104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1409_3_lut (.I0(n1995), .I1(n2060[30]), .I2(n2027), 
            .I3(GND_net), .O(n2094));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1558 (.I0(n2094), .I1(n2093), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i1_2_lut_adj_1558.LUT_INIT = 16'heeee;
    SB_LUT4 i7_2_lut (.I0(n2104), .I1(n2108), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4997));
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(CLK_c), .D(n29639));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i13_4_lut_adj_1559 (.I0(n2107), .I1(n2103), .I2(n2105), .I3(n18), 
            .O(n30_adj_4998));
    defparam i13_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(CLK_c), .D(n29638));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i11_4_lut_adj_1560 (.I0(n2099), .I1(n2101), .I2(n2100), .I3(n2106), 
            .O(n28_adj_4999));
    defparam i11_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1561 (.I0(bit_ctr[14]), .I1(n24_adj_4997), .I2(n2102), 
            .I3(n2109), .O(n29_adj_5000));
    defparam i12_4_lut_adj_1561.LUT_INIT = 16'hfefc;
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(CLK_c), .D(n29637));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(CLK_c), .D(n29636));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(CLK_c), .D(n29635));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(CLK_c), .D(n29634));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i10_4_lut_adj_1562 (.I0(n2095), .I1(n2097), .I2(n2096), .I3(n2098), 
            .O(n27_adj_5001));
    defparam i10_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1563 (.I0(n27_adj_5001), .I1(n29_adj_5000), .I2(n28_adj_4999), 
            .I3(n30_adj_4998), .O(n2126));
    defparam i16_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(CLK_c), .D(n29633));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(CLK_c), .D(n29632));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(CLK_c), .D(n29631));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(CLK_c), .D(n29630));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(CLK_c), .D(n29629));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(CLK_c), .D(n29628));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(CLK_c), .D(n29627));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(CLK_c), .D(n29626));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(CLK_c), .D(n29625));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(CLK_c), .D(n29624));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(CLK_c), .D(n29623));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(CLK_c), .D(n29622));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(CLK_c), .D(n29621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_33_lut (.I0(n50003), .I1(timer[31]), .I2(n1[31]), 
            .I3(n40603), .O(n27952)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n50001), .I1(timer[30]), .I2(n1[30]), 
            .I3(n40602), .O(n50003)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n40602), .I0(timer[30]), .I1(n1[30]), 
            .CO(n40603));
    SB_LUT4 sub_14_add_2_31_lut (.I0(n49999), .I1(timer[29]), .I2(n1[29]), 
            .I3(n40601), .O(n50001)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i34909_3_lut (.I0(neopxl_color[8]), .I1(neopxl_color[9]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n50391));
    defparam i34909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34910_3_lut (.I0(neopxl_color[10]), .I1(neopxl_color[11]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50392));
    defparam i34910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34913_3_lut (.I0(neopxl_color[14]), .I1(neopxl_color[15]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50395));
    defparam i34913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34912_3_lut (.I0(neopxl_color[12]), .I1(neopxl_color[13]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50394));
    defparam i34912_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR bit_ctr_2058__i7 (.Q(bit_ctr[7]), .C(CLK_c), .E(n6801), 
            .D(n133[7]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_CARRY sub_14_add_2_31 (.CI(n40601), .I0(timer[29]), .I1(n1[29]), 
            .CO(n40602));
    SB_LUT4 mod_5_i1344_3_lut (.I0(n1898), .I1(n1961[28]), .I2(n1928), 
            .I3(GND_net), .O(n1997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1343_3_lut (.I0(n1897), .I1(n1961[29]), .I2(n1928), 
            .I3(GND_net), .O(n1996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_add_2_30_lut (.I0(n49997), .I1(timer[28]), .I2(n1[28]), 
            .I3(n40600), .O(n49999)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_DFFESR bit_ctr_2058__i6 (.Q(bit_ctr[6]), .C(CLK_c), .E(n6801), 
            .D(n133[6]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_i1342_3_lut (.I0(n1896), .I1(n1961[30]), .I2(n1928), 
            .I3(GND_net), .O(n1995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1347_3_lut (.I0(n1901), .I1(n1961[25]), .I2(n1928), 
            .I3(GND_net), .O(n2000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1355_3_lut (.I0(n1909), .I1(n1961[17]), .I2(n1928), 
            .I3(GND_net), .O(n2008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1355_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR bit_ctr_2058__i5 (.Q(bit_ctr[5]), .C(CLK_c), .E(n6801), 
            .D(n133[5]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_i1353_3_lut (.I0(n1907), .I1(n1961[19]), .I2(n1928), 
            .I3(GND_net), .O(n2006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1349_3_lut (.I0(n1903), .I1(n1961[23]), .I2(n1928), 
            .I3(GND_net), .O(n2002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1346_3_lut (.I0(n1900), .I1(n1961[26]), .I2(n1928), 
            .I3(GND_net), .O(n1999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1350_3_lut (.I0(n1904), .I1(n1961[22]), .I2(n1928), 
            .I3(GND_net), .O(n2003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1345_3_lut (.I0(n1899), .I1(n1961[27]), .I2(n1928), 
            .I3(GND_net), .O(n1998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1351_3_lut (.I0(n1905), .I1(n1961[21]), .I2(n1928), 
            .I3(GND_net), .O(n2004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1354_3_lut (.I0(n1908), .I1(n1961[18]), .I2(n1928), 
            .I3(GND_net), .O(n2007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1352_3_lut (.I0(n1906), .I1(n1961[20]), .I2(n1928), 
            .I3(GND_net), .O(n2005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1348_3_lut (.I0(n1902), .I1(n1961[24]), .I2(n1928), 
            .I3(GND_net), .O(n2001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1356_3_lut (.I0(bit_ctr[16]), .I1(n1961[16]), .I2(n1928), 
            .I3(GND_net), .O(n2009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22748_2_lut (.I0(bit_ctr[15]), .I1(n2009), .I2(GND_net), 
            .I3(GND_net), .O(n36276));
    defparam i22748_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1564 (.I0(n2001), .I1(n2005), .I2(n2007), .I3(n2004), 
            .O(n28_adj_5004));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1565 (.I0(n1998), .I1(n2003), .I2(n1999), .I3(n36276), 
            .O(n26));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1566 (.I0(n2002), .I1(n2006), .I2(n2008), .I3(n2000), 
            .O(n27_adj_5005));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1995), .I1(n1996), .I2(n1994), .I3(n1997), 
            .O(n25_adj_5006));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1567 (.I0(n25_adj_5006), .I1(n27_adj_5005), .I2(n26), 
            .I3(n28_adj_5004), .O(n2027));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_30 (.CI(n40600), .I0(timer[28]), .I1(n1[28]), 
            .CO(n40601));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(CLK_c), .E(n29252), .D(state_3__N_528[0]), 
            .S(n29377));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2918), .I1(n2885), .I2(VCC_net), 
            .I3(n41597), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(GND_net), .I1(n2886), .I2(VCC_net), 
            .I3(n41596), .O(n2951[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_26 (.CI(n41596), .I0(n2886), .I1(VCC_net), 
            .CO(n41597));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(GND_net), .I1(n2887), .I2(VCC_net), 
            .I3(n41595), .O(n2951[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_25 (.CI(n41595), .I0(n2887), .I1(VCC_net), 
            .CO(n41596));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(GND_net), .I1(n2888), .I2(VCC_net), 
            .I3(n41594), .O(n2951[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_24 (.CI(n41594), .I0(n2888), .I1(VCC_net), 
            .CO(n41595));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(GND_net), .I1(n2889), .I2(VCC_net), 
            .I3(n41593), .O(n2951[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_23 (.CI(n41593), .I0(n2889), .I1(VCC_net), 
            .CO(n41594));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(GND_net), .I1(n2890), .I2(VCC_net), 
            .I3(n41592), .O(n2951[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_22 (.CI(n41592), .I0(n2890), .I1(VCC_net), 
            .CO(n41593));
    SB_LUT4 mod_5_i1287_3_lut (.I0(n1809), .I1(n1862[18]), .I2(n1829), 
            .I3(GND_net), .O(n1908));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1281_3_lut (.I0(n1803), .I1(n1862[24]), .I2(n1829), 
            .I3(GND_net), .O(n1902));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1280_3_lut (.I0(n1802), .I1(n1862[25]), .I2(n1829), 
            .I3(GND_net), .O(n1901));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2009_21_lut (.I0(GND_net), .I1(n2891), .I2(VCC_net), 
            .I3(n41591), .O(n2951[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1279_3_lut (.I0(n1801), .I1(n1862[26]), .I2(n1829), 
            .I3(GND_net), .O(n1900));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1279_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_2009_21 (.CI(n41591), .I0(n2891), .I1(VCC_net), 
            .CO(n41592));
    SB_LUT4 bit_ctr_2058_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[31]), 
            .I3(n41786), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_20_lut (.I0(GND_net), .I1(n2892), .I2(VCC_net), 
            .I3(n41590), .O(n2951[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1277_3_lut (.I0(n1799), .I1(n1862[28]), .I2(n1829), 
            .I3(GND_net), .O(n1898));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1278_3_lut (.I0(n1800), .I1(n1862[27]), .I2(n1829), 
            .I3(GND_net), .O(n1899));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1276_3_lut (.I0(n1798), .I1(n1862[29]), .I2(n1829), 
            .I3(GND_net), .O(n1897));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1276_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_2009_20 (.CI(n41590), .I0(n2892), .I1(VCC_net), 
            .CO(n41591));
    SB_LUT4 mod_5_i1275_3_lut (.I0(n1797), .I1(n1862[30]), .I2(n1829), 
            .I3(GND_net), .O(n1896));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1283_3_lut (.I0(n1805), .I1(n1862[22]), .I2(n1829), 
            .I3(GND_net), .O(n1904));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1282_3_lut (.I0(n1804), .I1(n1862[23]), .I2(n1829), 
            .I3(GND_net), .O(n1903));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1285_3_lut (.I0(n1807), .I1(n1862[20]), .I2(n1829), 
            .I3(GND_net), .O(n1906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1284_3_lut (.I0(n1806), .I1(n1862[21]), .I2(n1829), 
            .I3(GND_net), .O(n1905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1288_3_lut (.I0(bit_ctr[17]), .I1(n1862[17]), .I2(n1829), 
            .I3(GND_net), .O(n1909));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1286_3_lut (.I0(n1808), .I1(n1862[19]), .I2(n1829), 
            .I3(GND_net), .O(n1907));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2009_19_lut (.I0(GND_net), .I1(n2893), .I2(VCC_net), 
            .I3(n41589), .O(n2951[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(CLK_c), .D(n29620));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_29_lut (.I0(n49995), .I1(timer[27]), .I2(n1[27]), 
            .I3(n40599), .O(n49997)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2009_19 (.CI(n41589), .I0(n2893), .I1(VCC_net), 
            .CO(n41590));
    SB_LUT4 i5_3_lut_adj_1568 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), 
            .I3(GND_net), .O(n20));
    defparam i5_3_lut_adj_1568.LUT_INIT = 16'heaea;
    SB_LUT4 i11_4_lut_adj_1569 (.I0(n1905), .I1(n1906), .I2(n1903), .I3(n1904), 
            .O(n26_adj_5008));
    defparam i11_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_18_lut (.I0(GND_net), .I1(n2894), .I2(VCC_net), 
            .I3(n41588), .O(n2951[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1570 (.I0(n1896), .I1(n1895), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_5009));
    defparam i1_2_lut_adj_1570.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1571 (.I0(n1897), .I1(n1899), .I2(n1898), .I3(n1900), 
            .O(n24_adj_5010));
    defparam i9_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1572 (.I0(n1901), .I1(n26_adj_5008), .I2(n20), 
            .I3(n1902), .O(n28_adj_5011));
    defparam i13_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1573 (.I0(n1908), .I1(n28_adj_5011), .I2(n24_adj_5010), 
            .I3(n16_adj_5009), .O(n1928));
    defparam i14_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_18 (.CI(n41588), .I0(n2894), .I1(VCC_net), 
            .CO(n41589));
    SB_CARRY sub_14_add_2_29 (.CI(n40599), .I0(timer[27]), .I1(n1[27]), 
            .CO(n40600));
    SB_LUT4 mod_5_i1216_3_lut (.I0(n1706), .I1(n1763[22]), .I2(n1730), 
            .I3(GND_net), .O(n1805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1213_3_lut (.I0(n1703), .I1(n1763[25]), .I2(n1730), 
            .I3(GND_net), .O(n1802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1217_3_lut (.I0(n1707), .I1(n1763[21]), .I2(n1730), 
            .I3(GND_net), .O(n1806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1211_3_lut (.I0(n1701), .I1(n1763[27]), .I2(n1730), 
            .I3(GND_net), .O(n1800));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1210_3_lut (.I0(n1700), .I1(n1763[28]), .I2(n1730), 
            .I3(GND_net), .O(n1799));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1209_3_lut (.I0(n1699), .I1(n1763[29]), .I2(n1730), 
            .I3(GND_net), .O(n1798));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1433), .I1(n1400), .I2(VCC_net), 
            .I3(n41091), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_i1208_3_lut (.I0(n1698), .I1(n1763[30]), .I2(n1730), 
            .I3(GND_net), .O(n1797));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1220_3_lut (.I0(bit_ctr[18]), .I1(n1763[18]), .I2(n1730), 
            .I3(GND_net), .O(n1809));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1215_3_lut (.I0(n1705), .I1(n1763[23]), .I2(n1730), 
            .I3(GND_net), .O(n1804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_ctr_2058_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[30]), 
            .I3(n41785), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1219_3_lut (.I0(n1709), .I1(n1763[19]), .I2(n1730), 
            .I3(GND_net), .O(n1808));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2009_17_lut (.I0(GND_net), .I1(n2895), .I2(VCC_net), 
            .I3(n41587), .O(n2951[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_32 (.CI(n41785), .I0(GND_net), .I1(bit_ctr[30]), 
            .CO(n41786));
    SB_LUT4 mod_5_i1212_3_lut (.I0(n1702), .I1(n1763[26]), .I2(n1730), 
            .I3(GND_net), .O(n1801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1212_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_2009_17 (.CI(n41587), .I0(n2895), .I1(VCC_net), 
            .CO(n41588));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(GND_net), .I1(n2896), .I2(VCC_net), 
            .I3(n41586), .O(n2951[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_16 (.CI(n41586), .I0(n2896), .I1(VCC_net), 
            .CO(n41587));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(GND_net), .I1(n2897), .I2(VCC_net), 
            .I3(n41585), .O(n2951[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1214_3_lut (.I0(n1704), .I1(n1763[24]), .I2(n1730), 
            .I3(GND_net), .O(n1803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1218_3_lut (.I0(n1708), .I1(n1763[20]), .I2(n1730), 
            .I3(GND_net), .O(n1807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1574 (.I0(n1807), .I1(n1803), .I2(n1801), .I3(n1808), 
            .O(n24_adj_5012));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[17]), .I1(n1804), .I2(n1809), .I3(GND_net), 
            .O(n17));   // verilog/neopixel.v(22[26:36])
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut (.I0(n1797), .I1(n1798), .I2(n1796), .I3(n1799), 
            .O(n22_adj_5013));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1575 (.I0(n17), .I1(n24_adj_5012), .I2(n1800), 
            .I3(n1806), .O(n26_adj_5014));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1576 (.I0(n1802), .I1(n26_adj_5014), .I2(n22_adj_5013), 
            .I3(n1805), .O(n1829));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_15 (.CI(n41585), .I0(n2897), .I1(VCC_net), 
            .CO(n41586));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(GND_net), .I1(n2898), .I2(VCC_net), 
            .I3(n41584), .O(n2951[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_14 (.CI(n41584), .I0(n2898), .I1(VCC_net), 
            .CO(n41585));
    SB_LUT4 mod_5_add_1004_11_lut (.I0(GND_net), .I1(n1401), .I2(VCC_net), 
            .I3(n41090), .O(n1466[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_13_lut (.I0(GND_net), .I1(n2899), .I2(VCC_net), 
            .I3(n41583), .O(n2951[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_28_lut (.I0(n49993), .I1(timer[26]), .I2(n1[26]), 
            .I3(n40598), .O(n49995)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2009_13 (.CI(n41583), .I0(n2899), .I1(VCC_net), 
            .CO(n41584));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(GND_net), .I1(n2900), .I2(VCC_net), 
            .I3(n41582), .O(n2951[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_12 (.CI(n41582), .I0(n2900), .I1(VCC_net), 
            .CO(n41583));
    SB_LUT4 i3_3_lut_adj_1577 (.I0(n1699), .I1(bit_ctr[18]), .I2(n1709), 
            .I3(GND_net), .O(n16_adj_5016));
    defparam i3_3_lut_adj_1577.LUT_INIT = 16'heaea;
    SB_LUT4 i9_4_lut_adj_1578 (.I0(n1702), .I1(n1704), .I2(n1703), .I3(n1705), 
            .O(n22_adj_5017));
    defparam i9_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_11_lut (.I0(GND_net), .I1(n2901), .I2(VCC_net), 
            .I3(n41581), .O(n2951[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_3_lut_adj_1579 (.I0(n1707), .I1(n1698), .I2(n1697), .I3(GND_net), 
            .O(n20_adj_5018));
    defparam i7_3_lut_adj_1579.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1580 (.I0(n1701), .I1(n22_adj_5017), .I2(n16_adj_5016), 
            .I3(n1700), .O(n24_adj_5019));
    defparam i11_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_11 (.CI(n41581), .I0(n2901), .I1(VCC_net), 
            .CO(n41582));
    SB_LUT4 i12_4_lut_adj_1581 (.I0(n1706), .I1(n24_adj_5019), .I2(n20_adj_5018), 
            .I3(n1708), .O(n1730));
    defparam i12_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_10_lut (.I0(GND_net), .I1(n2902), .I2(VCC_net), 
            .I3(n41580), .O(n2951[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_10 (.CI(n41580), .I0(n2902), .I1(VCC_net), 
            .CO(n41581));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(GND_net), .I1(n2903), .I2(VCC_net), 
            .I3(n41579), .O(n2951[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_11 (.CI(n41090), .I0(n1401), .I1(VCC_net), 
            .CO(n41091));
    SB_CARRY mod_5_add_2009_9 (.CI(n41579), .I0(n2903), .I1(VCC_net), 
            .CO(n41580));
    SB_CARRY sub_14_add_2_28 (.CI(n40598), .I0(timer[26]), .I1(n1[26]), 
            .CO(n40599));
    SB_LUT4 i37614_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53097));
    defparam i37614_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1004_10_lut (.I0(GND_net), .I1(n1402), .I2(VCC_net), 
            .I3(n41089), .O(n1466[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_8_lut (.I0(GND_net), .I1(n2904), .I2(VCC_net), 
            .I3(n41578), .O(n2951[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_8 (.CI(n41578), .I0(n2904), .I1(VCC_net), 
            .CO(n41579));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(GND_net), .I1(n2905), .I2(VCC_net), 
            .I3(n41577), .O(n2951[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_7 (.CI(n41577), .I0(n2905), .I1(VCC_net), 
            .CO(n41578));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(GND_net), .I1(n2906), .I2(VCC_net), 
            .I3(n41576), .O(n2951[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_6 (.CI(n41576), .I0(n2906), .I1(VCC_net), 
            .CO(n41577));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(GND_net), .I1(n2907), .I2(VCC_net), 
            .I3(n41575), .O(n2951[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_5 (.CI(n41575), .I0(n2907), .I1(VCC_net), 
            .CO(n41576));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(GND_net), .I1(n2908), .I2(VCC_net), 
            .I3(n41574), .O(n2951[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_4 (.CI(n41574), .I0(n2908), .I1(VCC_net), 
            .CO(n41575));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(GND_net), .I1(n2909), .I2(GND_net), 
            .I3(n41573), .O(n2951[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_3 (.CI(n41573), .I0(n2909), .I1(GND_net), 
            .CO(n41574));
    SB_LUT4 sub_14_add_2_27_lut (.I0(n49991), .I1(timer[25]), .I2(n1[25]), 
            .I3(n40597), .O(n49993)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2009_2_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(VCC_net), .O(n2951[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(GND_net), 
            .CO(n41573));
    SB_CARRY mod_5_add_1004_10 (.CI(n41089), .I0(n1402), .I1(VCC_net), 
            .CO(n41090));
    SB_LUT4 bit_ctr_2058_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[29]), 
            .I3(n41784), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_9_lut (.I0(GND_net), .I1(n1403), .I2(VCC_net), 
            .I3(n41088), .O(n1466[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_31 (.CI(n41784), .I0(GND_net), .I1(bit_ctr[29]), 
            .CO(n41785));
    SB_LUT4 bit_ctr_2058_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[28]), 
            .I3(n41783), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_9 (.CI(n41088), .I0(n1403), .I1(VCC_net), 
            .CO(n41089));
    SB_CARRY bit_ctr_2058_add_4_30 (.CI(n41783), .I0(GND_net), .I1(bit_ctr[28]), 
            .CO(n41784));
    SB_LUT4 bit_ctr_2058_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[27]), 
            .I3(n41782), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_27 (.CI(n40597), .I0(timer[25]), .I1(n1[25]), 
            .CO(n40598));
    SB_LUT4 sub_14_add_2_26_lut (.I0(n49989), .I1(timer[24]), .I2(n1[24]), 
            .I3(n40596), .O(n49991)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_CARRY bit_ctr_2058_add_4_29 (.CI(n41782), .I0(GND_net), .I1(bit_ctr[27]), 
            .CO(n41783));
    SB_LUT4 bit_ctr_2058_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[26]), 
            .I3(n41781), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_28 (.CI(n41781), .I0(GND_net), .I1(bit_ctr[26]), 
            .CO(n41782));
    SB_LUT4 bit_ctr_2058_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[25]), 
            .I3(n41780), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_27 (.CI(n41780), .I0(GND_net), .I1(bit_ctr[25]), 
            .CO(n41781));
    SB_LUT4 bit_ctr_2058_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[24]), 
            .I3(n41779), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_26 (.CI(n41779), .I0(GND_net), .I1(bit_ctr[24]), 
            .CO(n41780));
    SB_LUT4 mod_5_i1076_3_lut (.I0(n1502), .I1(n1565[28]), .I2(n1532), 
            .I3(GND_net), .O(n1601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1075_3_lut (.I0(n1501), .I1(n1565[29]), .I2(n1532), 
            .I3(GND_net), .O(n1600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1078_3_lut (.I0(n1504), .I1(n1565[26]), .I2(n1532), 
            .I3(GND_net), .O(n1603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1074_3_lut (.I0(n1500), .I1(n1565[30]), .I2(n1532), 
            .I3(GND_net), .O(n1599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1082_3_lut (.I0(n1508), .I1(n1565[22]), .I2(n1532), 
            .I3(GND_net), .O(n1607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1079_3_lut (.I0(n1505), .I1(n1565[25]), .I2(n1532), 
            .I3(GND_net), .O(n1604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1012_3_lut (.I0(n1406), .I1(n1466[25]), .I2(n1433), 
            .I3(GND_net), .O(n1505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_ctr_2058_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[23]), 
            .I3(n41778), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_25 (.CI(n41778), .I0(GND_net), .I1(bit_ctr[23]), 
            .CO(n41779));
    SB_LUT4 mod_5_i1007_3_lut (.I0(n1401), .I1(n1466[30]), .I2(n1433), 
            .I3(GND_net), .O(n1500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1013_3_lut (.I0(n1407), .I1(n1466[24]), .I2(n1433), 
            .I3(GND_net), .O(n1506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1015_3_lut (.I0(n1409), .I1(n1466[22]), .I2(n1433), 
            .I3(GND_net), .O(n1508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1014_3_lut (.I0(n1408), .I1(n1466[23]), .I2(n1433), 
            .I3(GND_net), .O(n1507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1011_3_lut (.I0(n1405), .I1(n1466[26]), .I2(n1433), 
            .I3(GND_net), .O(n1504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1009_3_lut (.I0(n1403), .I1(n1466[28]), .I2(n1433), 
            .I3(GND_net), .O(n1502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1010_3_lut (.I0(n1404), .I1(n1466[27]), .I2(n1433), 
            .I3(GND_net), .O(n1503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1008_3_lut (.I0(n1402), .I1(n1466[29]), .I2(n1433), 
            .I3(GND_net), .O(n1501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_ctr_2058_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[22]), 
            .I3(n41777), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut (.I0(n1501), .I1(n1503), .I2(n1502), .I3(n1504), 
            .O(n18_adj_5021));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1582 (.I0(n1506), .I1(n18_adj_5021), .I2(n1500), 
            .I3(n1499), .O(n20_adj_5022));
    defparam i9_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(n1505), .I1(bit_ctr[20]), .I2(n1509), .I3(GND_net), 
            .O(n15));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_CARRY sub_14_add_2_26 (.CI(n40596), .I0(timer[24]), .I1(n1[24]), 
            .CO(n40597));
    SB_LUT4 i10_4_lut_adj_1583 (.I0(n15), .I1(n20_adj_5022), .I2(n1507), 
            .I3(n1508), .O(n1532));
    defparam i10_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_25_lut (.I0(n49987), .I1(timer[23]), .I2(n1[23]), 
            .I3(n40595), .O(n49989)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_i1016_3_lut (.I0(bit_ctr[21]), .I1(n1466[21]), .I2(n1433), 
            .I3(GND_net), .O(n1509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1083_3_lut (.I0(n1509), .I1(n1565[21]), .I2(n1532), 
            .I3(GND_net), .O(n1608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(GND_net), .I1(n1404), .I2(VCC_net), 
            .I3(n41087), .O(n1466[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_24 (.CI(n41777), .I0(GND_net), .I1(bit_ctr[22]), 
            .CO(n41778));
    SB_LUT4 mod_5_i1080_3_lut (.I0(n1506), .I1(n1565[24]), .I2(n1532), 
            .I3(GND_net), .O(n1605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1081_3_lut (.I0(n1507), .I1(n1565[23]), .I2(n1532), 
            .I3(GND_net), .O(n1606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1084_3_lut (.I0(bit_ctr[20]), .I1(n1565[20]), .I2(n1532), 
            .I3(GND_net), .O(n1609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1077_3_lut (.I0(n1503), .I1(n1565[27]), .I2(n1532), 
            .I3(GND_net), .O(n1602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut_adj_1584 (.I0(n1602), .I1(bit_ctr[19]), .I2(n1609), 
            .I3(GND_net), .O(n15_adj_5023));
    defparam i3_3_lut_adj_1584.LUT_INIT = 16'heaea;
    SB_LUT4 i7_4_lut_adj_1585 (.I0(n1606), .I1(n1605), .I2(n1608), .I3(n1598), 
            .O(n19));
    defparam i7_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut_adj_1586 (.I0(n1604), .I1(n1607), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5024));
    defparam i6_2_lut_adj_1586.LUT_INIT = 16'heeee;
    SB_LUT4 bit_ctr_2058_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[21]), 
            .I3(n41776), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_1587 (.I0(n19), .I1(n15_adj_5023), .I2(n1599), 
            .I3(n1603), .O(n22_adj_5025));
    defparam i10_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_CARRY bit_ctr_2058_add_4_23 (.CI(n41776), .I0(GND_net), .I1(bit_ctr[21]), 
            .CO(n41777));
    SB_LUT4 i11_4_lut_adj_1588 (.I0(n1600), .I1(n22_adj_5025), .I2(n18_adj_5024), 
            .I3(n1601), .O(n1631));
    defparam i11_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_2058_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[20]), 
            .I3(n41775), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_22 (.CI(n41775), .I0(GND_net), .I1(bit_ctr[20]), 
            .CO(n41776));
    SB_LUT4 bit_ctr_2058_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[19]), 
            .I3(n41774), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_25 (.CI(n40595), .I0(timer[23]), .I1(n1[23]), 
            .CO(n40596));
    SB_CARRY bit_ctr_2058_add_4_21 (.CI(n41774), .I0(GND_net), .I1(bit_ctr[19]), 
            .CO(n41775));
    SB_LUT4 bit_ctr_2058_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[18]), 
            .I3(n41773), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_8 (.CI(n41087), .I0(n1404), .I1(VCC_net), 
            .CO(n41088));
    SB_LUT4 sub_14_add_2_24_lut (.I0(n49985), .I1(timer[22]), .I2(n1[22]), 
            .I3(n40594), .O(n49987)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n40594), .I0(timer[22]), .I1(n1[22]), 
            .CO(n40595));
    SB_CARRY bit_ctr_2058_add_4_20 (.CI(n41773), .I0(GND_net), .I1(bit_ctr[18]), 
            .CO(n41774));
    SB_LUT4 bit_ctr_2058_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[17]), 
            .I3(n41772), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_19 (.CI(n41772), .I0(GND_net), .I1(bit_ctr[17]), 
            .CO(n41773));
    SB_LUT4 bit_ctr_2058_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[16]), 
            .I3(n41771), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_18 (.CI(n41771), .I0(GND_net), .I1(bit_ctr[16]), 
            .CO(n41772));
    SB_LUT4 bit_ctr_2058_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[15]), 
            .I3(n41770), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_17 (.CI(n41770), .I0(GND_net), .I1(bit_ctr[15]), 
            .CO(n41771));
    SB_LUT4 i37613_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53096));
    defparam i37613_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2058_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[14]), 
            .I3(n41769), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_16 (.CI(n41769), .I0(GND_net), .I1(bit_ctr[14]), 
            .CO(n41770));
    SB_CARRY bit_ctr_2058_add_4_9 (.CI(n41762), .I0(GND_net), .I1(bit_ctr[7]), 
            .CO(n41763));
    SB_LUT4 sub_14_add_2_23_lut (.I0(n49983), .I1(timer[21]), .I2(n1[21]), 
            .I3(n40593), .O(n49985)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_23 (.CI(n40593), .I0(timer[21]), .I1(n1[21]), 
            .CO(n40594));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(GND_net), .I1(n1405), .I2(VCC_net), 
            .I3(n41086), .O(n1466[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_7 (.CI(n41086), .I0(n1405), .I1(VCC_net), 
            .CO(n41087));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(GND_net), .I1(n1406), .I2(VCC_net), 
            .I3(n41085), .O(n1466[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_6 (.CI(n41085), .I0(n1406), .I1(VCC_net), 
            .CO(n41086));
    SB_LUT4 sub_14_add_2_22_lut (.I0(n49981), .I1(timer[20]), .I2(n1[20]), 
            .I3(n40592), .O(n49983)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1004_5_lut (.I0(GND_net), .I1(n1407), .I2(VCC_net), 
            .I3(n41084), .O(n1466[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_5 (.CI(n41084), .I0(n1407), .I1(VCC_net), 
            .CO(n41085));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(GND_net), .I1(n1408), .I2(VCC_net), 
            .I3(n41083), .O(n1466[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_4 (.CI(n41083), .I0(n1408), .I1(VCC_net), 
            .CO(n41084));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(GND_net), .I1(n1409), .I2(GND_net), 
            .I3(n41082), .O(n1466[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_22 (.CI(n40592), .I0(timer[20]), .I1(n1[20]), 
            .CO(n40593));
    SB_LUT4 i4_3_lut_adj_1589 (.I0(bit_ctr[23]), .I1(n1207), .I2(n1209), 
            .I3(GND_net), .O(n12_adj_5026));
    defparam i4_3_lut_adj_1589.LUT_INIT = 16'hecec;
    SB_LUT4 i5_4_lut (.I0(n1205), .I1(n1204), .I2(n1206), .I3(n1208), 
            .O(n13_adj_5027));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1590 (.I0(n13_adj_5027), .I1(n1203), .I2(n12_adj_5026), 
            .I3(n1202), .O(n1235));
    defparam i7_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 i37612_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53095));
    defparam i37612_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1004_3 (.CI(n41082), .I0(n1409), .I1(GND_net), 
            .CO(n41083));
    SB_LUT4 sub_14_add_2_21_lut (.I0(n49979), .I1(timer[19]), .I2(n1[19]), 
            .I3(n40591), .O(n49981)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1004_2_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(VCC_net), .O(n1466[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22738_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n36266));
    defparam i22738_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1591 (.I0(n1106), .I1(n1103), .I2(n1108), .I3(n36266), 
            .O(n12_adj_5028));
    defparam i5_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1592 (.I0(n1107), .I1(n12_adj_5028), .I2(n1105), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(GND_net), 
            .CO(n41082));
    SB_CARRY sub_14_add_2_21 (.CI(n40591), .I0(timer[19]), .I1(n1[19]), 
            .CO(n40592));
    SB_LUT4 sub_14_add_2_20_lut (.I0(n49977), .I1(timer[18]), .I2(n1[18]), 
            .I3(n40590), .O(n49979)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_20 (.CI(n40590), .I0(timer[18]), .I1(n1[18]), 
            .CO(n40591));
    SB_LUT4 sub_14_add_2_19_lut (.I0(n49975), .I1(timer[17]), .I2(n1[17]), 
            .I3(n40589), .O(n49977)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_2058_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[13]), 
            .I3(n41768), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_19 (.CI(n40589), .I0(timer[17]), .I1(n1[17]), 
            .CO(n40590));
    SB_LUT4 sub_14_add_2_18_lut (.I0(n49973), .I1(timer[16]), .I2(n1[16]), 
            .I3(n40588), .O(n49975)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(CLK_c), .D(n29619));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(CLK_c), .D(n29618));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(CLK_c), .D(n29617));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(CLK_c), .D(n29616));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(CLK_c), .D(n29615));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(CLK_c), .D(n29614));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(CLK_c), .D(n29613));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(CLK_c), .D(n29612));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(CLK_c), .D(n29611));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(CLK_c), .D(n29610));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(CLK_c), .D(n29609));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_2058__i4 (.Q(bit_ctr[4]), .C(CLK_c), .E(n6801), 
            .D(n133[4]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_CARRY sub_14_add_2_18 (.CI(n40588), .I0(timer[16]), .I1(n1[16]), 
            .CO(n40589));
    SB_LUT4 sub_14_add_2_17_lut (.I0(n49971), .I1(timer[15]), .I2(n1[15]), 
            .I3(n40587), .O(n49973)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_DFF timer_2057__i0 (.Q(timer[0]), .C(CLK_c), .D(n133_adj_5095[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY sub_14_add_2_17 (.CI(n40587), .I0(timer[15]), .I1(n1[15]), 
            .CO(n40588));
    SB_CARRY bit_ctr_2058_add_4_15 (.CI(n41768), .I0(GND_net), .I1(bit_ctr[13]), 
            .CO(n41769));
    SB_LUT4 bit_ctr_2058_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[12]), 
            .I3(n41767), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_14 (.CI(n41767), .I0(GND_net), .I1(bit_ctr[12]), 
            .CO(n41768));
    SB_LUT4 bit_ctr_2058_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[11]), 
            .I3(n41766), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_13 (.CI(n41766), .I0(GND_net), .I1(bit_ctr[11]), 
            .CO(n41767));
    SB_LUT4 bit_ctr_2058_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[10]), 
            .I3(n41765), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_12 (.CI(n41765), .I0(GND_net), .I1(bit_ctr[10]), 
            .CO(n41766));
    SB_LUT4 bit_ctr_2058_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[9]), 
            .I3(n41764), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_11 (.CI(n41764), .I0(GND_net), .I1(bit_ctr[9]), 
            .CO(n41765));
    SB_LUT4 bit_ctr_2058_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[8]), 
            .I3(n41763), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_10 (.CI(n41763), .I0(GND_net), .I1(bit_ctr[8]), 
            .CO(n41764));
    SB_LUT4 bit_ctr_2058_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[7]), 
            .I3(n41762), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_16_lut (.I0(n49969), .I1(timer[14]), .I2(n1[14]), 
            .I3(n40586), .O(n49971)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_16 (.CI(n40586), .I0(timer[14]), .I1(n1[14]), 
            .CO(n40587));
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_15_lut (.I0(n49967), .I1(timer[13]), .I2(n1[13]), 
            .I3(n40585), .O(n49969)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_15 (.CI(n40585), .I0(timer[13]), .I1(n1[13]), 
            .CO(n40586));
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_679[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n40584), .O(n49967)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_14 (.CI(n40584), .I0(timer[12]), .I1(n1[12]), 
            .CO(n40585));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n40583), .O(one_wire_N_679[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n40583), .I0(timer[11]), .I1(n1[11]), 
            .CO(n40584));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n40582), .O(one_wire_N_679[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n40582), .I0(timer[10]), .I1(n1[10]), 
            .CO(n40583));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n40581), .O(one_wire_N_679[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n40581), .I0(timer[9]), .I1(n1[9]), 
            .CO(n40582));
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n40580), .O(one_wire_N_679[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n40580), .I0(timer[8]), .I1(n1[8]), 
            .CO(n40581));
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_2058__i3 (.Q(bit_ctr[3]), .C(CLK_c), .E(n6801), 
            .D(n133[3]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i2 (.Q(bit_ctr[2]), .C(CLK_c), .E(n6801), 
            .D(n133[2]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n40579), .O(one_wire_N_679[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n40579), .I0(timer[7]), .I1(n1[7]), .CO(n40580));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n40578), .O(one_wire_N_679[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n40578), .I0(timer[6]), .I1(n1[6]), .CO(n40579));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n40577), .O(one_wire_N_679[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n40577), .I0(timer[5]), .I1(n1[5]), .CO(n40578));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n40576), .O(one_wire_N_679[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_6 (.CI(n40576), .I0(timer[4]), .I1(n1[4]), .CO(n40577));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n40575), .O(one_wire_N_679[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n40575), .I0(timer[3]), .I1(n1[3]), .CO(n40576));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n40574), .O(one_wire_N_679[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n40574), .I0(timer[2]), .I1(n1[2]), .CO(n40575));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_679[3]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n40573), .O(n4_adj_4976)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_3 (.CI(n40573), .I0(timer[1]), .I1(n1[1]), .CO(n40574));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n40573));
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34915_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n50397));
    defparam i34915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34916_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n50398));
    defparam i34916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34919_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n50401));
    defparam i34919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1593 (.I0(n1307), .I1(n1302), .I2(n1301), .I3(GND_net), 
            .O(n14_adj_5046));   // verilog/neopixel.v(22[26:36])
    defparam i5_3_lut_adj_1593.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_2_lut (.I0(n1305), .I1(n1306), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_5047));   // verilog/neopixel.v(22[26:36])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1594 (.I0(bit_ctr[22]), .I1(n14_adj_5046), .I2(n1308), 
            .I3(n1309), .O(n16_adj_5048));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1594.LUT_INIT = 16'hfefc;
    SB_LUT4 i8_4_lut_adj_1595 (.I0(n1303), .I1(n16_adj_5048), .I2(n12_adj_5047), 
            .I3(n1304), .O(n1334));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i34918_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n50400));
    defparam i34918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n42233), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n42232), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n42232), .I0(n1104), .I1(n1136), .CO(n42233));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n42231), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n42231), .I0(n1105), .I1(n1136), .CO(n42232));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n42230), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n42230), .I0(n1106), .I1(n1136), .CO(n42231));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n42229), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n42229), .I0(n1107), .I1(n1136), .CO(n42230));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n42228), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n42228), .I0(n1108), .I1(n1136), .CO(n42229));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n53095), 
            .I3(n42227), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n42227), .I0(n1109), .I1(n53095), .CO(n42228));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n53095), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n53095), 
            .CO(n42227));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n42226), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n42225), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n42225), .I0(n1203), .I1(n1235), .CO(n42226));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n42224), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_870_8 (.CI(n42224), .I0(n1204), .I1(n1235), .CO(n42225));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n42223), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n42223), .I0(n1205), .I1(n1235), .CO(n42224));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n42222), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n42222), .I0(n1206), .I1(n1235), .CO(n42223));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n42221), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n42221), .I0(n1207), .I1(n1235), .CO(n42222));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n42220), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n42220), .I0(n1208), .I1(n1235), .CO(n42221));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n53096), 
            .I3(n42219), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n42219), .I0(n1209), .I1(n53096), .CO(n42220));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n53096), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n53096), 
            .CO(n42219));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n42218), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n42217), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_13 (.CI(n42217), .I0(n1599), .I1(n1631), .CO(n42218));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n42216), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n42216), .I0(n1600), .I1(n1631), .CO(n42217));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n42215), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n42215), .I0(n1601), .I1(n1631), .CO(n42216));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n42214), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n42214), .I0(n1602), .I1(n1631), .CO(n42215));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n42213), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n42213), .I0(n1603), .I1(n1631), .CO(n42214));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n42212), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1532), .I1(n1499), .I2(VCC_net), 
            .I3(n40741), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1138_8 (.CI(n42212), .I0(n1604), .I1(n1631), .CO(n42213));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n42211), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n42211), .I0(n1605), .I1(n1631), .CO(n42212));
    SB_LUT4 i36517_4_lut (.I0(n42258), .I1(n4), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n51824));
    defparam i36517_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n42210), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i53_4_lut (.I0(n51330), .I1(n36444), .I2(\state[1] ), .I3(n27768), 
            .O(n46577));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_CARRY mod_5_add_1138_6 (.CI(n42210), .I0(n1606), .I1(n1631), .CO(n42211));
    SB_LUT4 i52_4_lut (.I0(n46577), .I1(n51825), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n46623));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n42209), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n42209), .I0(n1607), .I1(n1631), .CO(n42210));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n42208), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i42_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_742 ));
    defparam i42_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1138_4 (.CI(n42208), .I0(n1608), .I1(n1631), .CO(n42209));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n53097), 
            .I3(n42207), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n42207), .I0(n1609), .I1(n53097), .CO(n42208));
    SB_LUT4 mod_5_add_1071_12_lut (.I0(GND_net), .I1(n1500), .I2(VCC_net), 
            .I3(n40740), .O(n1565[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n53097), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n53097), 
            .CO(n42207));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1730), .I1(n1697), .I2(VCC_net), 
            .I3(n42206), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(GND_net), .I1(n1698), .I2(VCC_net), 
            .I3(n42205), .O(n1763[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_14 (.CI(n42205), .I0(n1698), .I1(VCC_net), 
            .CO(n42206));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(GND_net), .I1(n1699), .I2(VCC_net), 
            .I3(n42204), .O(n1763[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_13 (.CI(n42204), .I0(n1699), .I1(VCC_net), 
            .CO(n42205));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(GND_net), .I1(n1700), .I2(VCC_net), 
            .I3(n42203), .O(n1763[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_12 (.CI(n42203), .I0(n1700), .I1(VCC_net), 
            .CO(n42204));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(GND_net), .I1(n1701), .I2(VCC_net), 
            .I3(n42202), .O(n1763[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_11 (.CI(n42202), .I0(n1701), .I1(VCC_net), 
            .CO(n42203));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(GND_net), .I1(n1702), .I2(VCC_net), 
            .I3(n42201), .O(n1763[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_10 (.CI(n42201), .I0(n1702), .I1(VCC_net), 
            .CO(n42202));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(GND_net), .I1(n1703), .I2(VCC_net), 
            .I3(n42200), .O(n1763[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_9 (.CI(n42200), .I0(n1703), .I1(VCC_net), 
            .CO(n42201));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(GND_net), .I1(n1704), .I2(VCC_net), 
            .I3(n42199), .O(n1763[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_12 (.CI(n40740), .I0(n1500), .I1(VCC_net), 
            .CO(n40741));
    SB_CARRY mod_5_add_1205_8 (.CI(n42199), .I0(n1704), .I1(VCC_net), 
            .CO(n42200));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(GND_net), .I1(n1705), .I2(VCC_net), 
            .I3(n42198), .O(n1763[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_7 (.CI(n42198), .I0(n1705), .I1(VCC_net), 
            .CO(n42199));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(GND_net), .I1(n1706), .I2(VCC_net), 
            .I3(n42197), .O(n1763[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_6 (.CI(n42197), .I0(n1706), .I1(VCC_net), 
            .CO(n42198));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(GND_net), .I1(n1707), .I2(VCC_net), 
            .I3(n42196), .O(n1763[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_5 (.CI(n42196), .I0(n1707), .I1(VCC_net), 
            .CO(n42197));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(GND_net), .I1(n1708), .I2(VCC_net), 
            .I3(n42195), .O(n1763[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_4 (.CI(n42195), .I0(n1708), .I1(VCC_net), 
            .CO(n42196));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(GND_net), .I1(n1709), .I2(GND_net), 
            .I3(n42194), .O(n1763[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_3 (.CI(n42194), .I0(n1709), .I1(GND_net), 
            .CO(n42195));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(VCC_net), .O(n1763[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(GND_net), 
            .CO(n42194));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1829), .I1(n1796), .I2(VCC_net), 
            .I3(n42193), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1071_11_lut (.I0(GND_net), .I1(n1501), .I2(VCC_net), 
            .I3(n40739), .O(n1565[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(GND_net), .I1(n1797), .I2(VCC_net), 
            .I3(n42192), .O(n1862[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_15 (.CI(n42192), .I0(n1797), .I1(VCC_net), 
            .CO(n42193));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(GND_net), .I1(n1798), .I2(VCC_net), 
            .I3(n42191), .O(n1862[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_14 (.CI(n42191), .I0(n1798), .I1(VCC_net), 
            .CO(n42192));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(GND_net), .I1(n1799), .I2(VCC_net), 
            .I3(n42190), .O(n1862[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_13 (.CI(n42190), .I0(n1799), .I1(VCC_net), 
            .CO(n42191));
    SB_CARRY mod_5_add_1071_11 (.CI(n40739), .I0(n1501), .I1(VCC_net), 
            .CO(n40740));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(GND_net), .I1(n1800), .I2(VCC_net), 
            .I3(n42189), .O(n1862[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_12 (.CI(n42189), .I0(n1800), .I1(VCC_net), 
            .CO(n42190));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(GND_net), .I1(n1801), .I2(VCC_net), 
            .I3(n42188), .O(n1862[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_11 (.CI(n42188), .I0(n1801), .I1(VCC_net), 
            .CO(n42189));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(GND_net), .I1(n1802), .I2(VCC_net), 
            .I3(n42187), .O(n1862[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_10 (.CI(n42187), .I0(n1802), .I1(VCC_net), 
            .CO(n42188));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(GND_net), .I1(n1803), .I2(VCC_net), 
            .I3(n42186), .O(n1862[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_9 (.CI(n42186), .I0(n1803), .I1(VCC_net), 
            .CO(n42187));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(GND_net), .I1(n1804), .I2(VCC_net), 
            .I3(n42185), .O(n1862[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_8 (.CI(n42185), .I0(n1804), .I1(VCC_net), 
            .CO(n42186));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(GND_net), .I1(n1805), .I2(VCC_net), 
            .I3(n42184), .O(n1862[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_10_lut (.I0(GND_net), .I1(n1502), .I2(VCC_net), 
            .I3(n40738), .O(n1565[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_7 (.CI(n42184), .I0(n1805), .I1(VCC_net), 
            .CO(n42185));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(GND_net), .I1(n1806), .I2(VCC_net), 
            .I3(n42183), .O(n1862[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_6 (.CI(n42183), .I0(n1806), .I1(VCC_net), 
            .CO(n42184));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(GND_net), .I1(n1807), .I2(VCC_net), 
            .I3(n42182), .O(n1862[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_5 (.CI(n42182), .I0(n1807), .I1(VCC_net), 
            .CO(n42183));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(GND_net), .I1(n1808), .I2(VCC_net), 
            .I3(n42181), .O(n1862[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_4 (.CI(n42181), .I0(n1808), .I1(VCC_net), 
            .CO(n42182));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(GND_net), .I1(n1809), .I2(GND_net), 
            .I3(n42180), .O(n1862[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_3 (.CI(n42180), .I0(n1809), .I1(GND_net), 
            .CO(n42181));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(VCC_net), .O(n1862[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(GND_net), 
            .CO(n42180));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1928), .I1(n1895), .I2(VCC_net), 
            .I3(n42179), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(GND_net), .I1(n1896), .I2(VCC_net), 
            .I3(n42178), .O(n1961[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_16 (.CI(n42178), .I0(n1896), .I1(VCC_net), 
            .CO(n42179));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(GND_net), .I1(n1897), .I2(VCC_net), 
            .I3(n42177), .O(n1961[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_15 (.CI(n42177), .I0(n1897), .I1(VCC_net), 
            .CO(n42178));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(GND_net), .I1(n1898), .I2(VCC_net), 
            .I3(n42176), .O(n1961[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_14 (.CI(n42176), .I0(n1898), .I1(VCC_net), 
            .CO(n42177));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(GND_net), .I1(n1899), .I2(VCC_net), 
            .I3(n42175), .O(n1961[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_13 (.CI(n42175), .I0(n1899), .I1(VCC_net), 
            .CO(n42176));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(GND_net), .I1(n1900), .I2(VCC_net), 
            .I3(n42174), .O(n1961[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_12 (.CI(n42174), .I0(n1900), .I1(VCC_net), 
            .CO(n42175));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(GND_net), .I1(n1901), .I2(VCC_net), 
            .I3(n42173), .O(n1961[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_11 (.CI(n42173), .I0(n1901), .I1(VCC_net), 
            .CO(n42174));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(GND_net), .I1(n1902), .I2(VCC_net), 
            .I3(n42172), .O(n1961[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_10 (.CI(n42172), .I0(n1902), .I1(VCC_net), 
            .CO(n42173));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(GND_net), .I1(n1903), .I2(VCC_net), 
            .I3(n42171), .O(n1961[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_9 (.CI(n42171), .I0(n1903), .I1(VCC_net), 
            .CO(n42172));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(GND_net), .I1(n1904), .I2(VCC_net), 
            .I3(n42170), .O(n1961[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_8 (.CI(n42170), .I0(n1904), .I1(VCC_net), 
            .CO(n42171));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(GND_net), .I1(n1905), .I2(VCC_net), 
            .I3(n42169), .O(n1961[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_7 (.CI(n42169), .I0(n1905), .I1(VCC_net), 
            .CO(n42170));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(GND_net), .I1(n1906), .I2(VCC_net), 
            .I3(n42168), .O(n1961[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_6 (.CI(n42168), .I0(n1906), .I1(VCC_net), 
            .CO(n42169));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(GND_net), .I1(n1907), .I2(VCC_net), 
            .I3(n42167), .O(n1961[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_5 (.CI(n42167), .I0(n1907), .I1(VCC_net), 
            .CO(n42168));
    SB_CARRY mod_5_add_1071_10 (.CI(n40738), .I0(n1502), .I1(VCC_net), 
            .CO(n40739));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(GND_net), .I1(n1908), .I2(VCC_net), 
            .I3(n42166), .O(n1961[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_4 (.CI(n42166), .I0(n1908), .I1(VCC_net), 
            .CO(n42167));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(GND_net), .I1(n1909), .I2(GND_net), 
            .I3(n42165), .O(n1961[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_3 (.CI(n42165), .I0(n1909), .I1(GND_net), 
            .CO(n42166));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(VCC_net), .O(n1961[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(GND_net), 
            .CO(n42165));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n2027), .I1(n1994), .I2(VCC_net), 
            .I3(n42164), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1071_9_lut (.I0(GND_net), .I1(n1503), .I2(VCC_net), 
            .I3(n40737), .O(n1565[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(GND_net), .I1(n1995), .I2(VCC_net), 
            .I3(n42163), .O(n2060[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_17 (.CI(n42163), .I0(n1995), .I1(VCC_net), 
            .CO(n42164));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(GND_net), .I1(n1996), .I2(VCC_net), 
            .I3(n42162), .O(n2060[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_16 (.CI(n42162), .I0(n1996), .I1(VCC_net), 
            .CO(n42163));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(GND_net), .I1(n1997), .I2(VCC_net), 
            .I3(n42161), .O(n2060[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_15 (.CI(n42161), .I0(n1997), .I1(VCC_net), 
            .CO(n42162));
    SB_CARRY mod_5_add_1071_9 (.CI(n40737), .I0(n1503), .I1(VCC_net), 
            .CO(n40738));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(GND_net), .I1(n1998), .I2(VCC_net), 
            .I3(n42160), .O(n2060[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_14 (.CI(n42160), .I0(n1998), .I1(VCC_net), 
            .CO(n42161));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(GND_net), .I1(n1999), .I2(VCC_net), 
            .I3(n42159), .O(n2060[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_13 (.CI(n42159), .I0(n1999), .I1(VCC_net), 
            .CO(n42160));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(GND_net), .I1(n1504), .I2(VCC_net), 
            .I3(n40736), .O(n1565[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_8 (.CI(n40736), .I0(n1504), .I1(VCC_net), 
            .CO(n40737));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(GND_net), .I1(n2000), .I2(VCC_net), 
            .I3(n42158), .O(n2060[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_12 (.CI(n42158), .I0(n2000), .I1(VCC_net), 
            .CO(n42159));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(GND_net), .I1(n2001), .I2(VCC_net), 
            .I3(n42157), .O(n2060[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_11 (.CI(n42157), .I0(n2001), .I1(VCC_net), 
            .CO(n42158));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(GND_net), .I1(n2002), .I2(VCC_net), 
            .I3(n42156), .O(n2060[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_10 (.CI(n42156), .I0(n2002), .I1(VCC_net), 
            .CO(n42157));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(GND_net), .I1(n2003), .I2(VCC_net), 
            .I3(n42155), .O(n2060[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_9 (.CI(n42155), .I0(n2003), .I1(VCC_net), 
            .CO(n42156));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(GND_net), .I1(n1505), .I2(VCC_net), 
            .I3(n40735), .O(n1565[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_1__bdd_4_lut (.I0(bit_ctr[1]), .I1(n50394), .I2(n50395), 
            .I3(bit_ctr[2]), .O(n53209));
    defparam bit_ctr_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n53209_bdd_4_lut (.I0(n53209), .I1(n50392), .I2(n50391), .I3(bit_ctr[2]), 
            .O(n53212));
    defparam n53209_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1406_8_lut (.I0(GND_net), .I1(n2004), .I2(VCC_net), 
            .I3(n42154), .O(n2060[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_8 (.CI(n42154), .I0(n2004), .I1(VCC_net), 
            .CO(n42155));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(GND_net), .I1(n2005), .I2(VCC_net), 
            .I3(n42153), .O(n2060[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_7 (.CI(n42153), .I0(n2005), .I1(VCC_net), 
            .CO(n42154));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(GND_net), .I1(n2006), .I2(VCC_net), 
            .I3(n42152), .O(n2060[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_6 (.CI(n42152), .I0(n2006), .I1(VCC_net), 
            .CO(n42153));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(GND_net), .I1(n2007), .I2(VCC_net), 
            .I3(n42151), .O(n2060[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_5 (.CI(n42151), .I0(n2007), .I1(VCC_net), 
            .CO(n42152));
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n40557), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37616_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53099));
    defparam i37616_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1406_4_lut (.I0(GND_net), .I1(n2008), .I2(VCC_net), 
            .I3(n42150), .O(n2060[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_4 (.CI(n42150), .I0(n2008), .I1(VCC_net), 
            .CO(n42151));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(GND_net), .I1(n2009), .I2(GND_net), 
            .I3(n42149), .O(n2060[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_3 (.CI(n42149), .I0(n2009), .I1(GND_net), 
            .CO(n42150));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(VCC_net), .O(n2060[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(GND_net), 
            .CO(n42149));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2126), .I1(n2093), .I2(VCC_net), 
            .I3(n42148), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(GND_net), .I1(n2094), .I2(VCC_net), 
            .I3(n42147), .O(n2159[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_18 (.CI(n42147), .I0(n2094), .I1(VCC_net), 
            .CO(n42148));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(GND_net), .I1(n2095), .I2(VCC_net), 
            .I3(n42146), .O(n2159[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_17 (.CI(n42146), .I0(n2095), .I1(VCC_net), 
            .CO(n42147));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(GND_net), .I1(n2096), .I2(VCC_net), 
            .I3(n42145), .O(n2159[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_16 (.CI(n42145), .I0(n2096), .I1(VCC_net), 
            .CO(n42146));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(GND_net), .I1(n2097), .I2(VCC_net), 
            .I3(n42144), .O(n2159[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_15 (.CI(n42144), .I0(n2097), .I1(VCC_net), 
            .CO(n42145));
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n40556), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_14_lut (.I0(GND_net), .I1(n2098), .I2(VCC_net), 
            .I3(n42143), .O(n2159[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_14 (.CI(n42143), .I0(n2098), .I1(VCC_net), 
            .CO(n42144));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(GND_net), .I1(n2099), .I2(VCC_net), 
            .I3(n42142), .O(n2159[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n40556), .I0(GND_net), .I1(VCC_net), 
            .CO(n40557));
    SB_CARRY mod_5_add_1473_13 (.CI(n42142), .I0(n2099), .I1(VCC_net), 
            .CO(n42143));
    SB_LUT4 i22654_2_lut (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(GND_net), .O(n36179));
    defparam i22654_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1596 (.I0(bit_ctr[8]), .I1(bit_ctr[18]), .I2(bit_ctr[24]), 
            .I3(bit_ctr[9]), .O(n48));
    defparam i20_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1071_7 (.CI(n40735), .I0(n1505), .I1(VCC_net), 
            .CO(n40736));
    SB_LUT4 bit_ctr_1__bdd_4_lut_37707 (.I0(bit_ctr[1]), .I1(n50445), .I2(n50446), 
            .I3(bit_ctr[2]), .O(n53167));
    defparam bit_ctr_1__bdd_4_lut_37707.LUT_INIT = 16'he4aa;
    SB_LUT4 n53167_bdd_4_lut (.I0(n53167), .I1(n50449), .I2(n50448), .I3(bit_ctr[2]), 
            .O(n53170));
    defparam n53167_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1473_12_lut (.I0(GND_net), .I1(n2100), .I2(VCC_net), 
            .I3(n42141), .O(n2159[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_12 (.CI(n42141), .I0(n2100), .I1(VCC_net), 
            .CO(n42142));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(GND_net), .I1(n2101), .I2(VCC_net), 
            .I3(n42140), .O(n2159[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_11 (.CI(n42140), .I0(n2101), .I1(VCC_net), 
            .CO(n42141));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(GND_net), .I1(n2102), .I2(VCC_net), 
            .I3(n42139), .O(n2159[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_10 (.CI(n42139), .I0(n2102), .I1(VCC_net), 
            .CO(n42140));
    SB_LUT4 i36914_2_lut (.I0(n971[28]), .I1(n2_adj_5049), .I2(GND_net), 
            .I3(GND_net), .O(n52397));   // verilog/neopixel.v(22[26:36])
    defparam i36914_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i18_4_lut_adj_1597 (.I0(bit_ctr[26]), .I1(bit_ctr[28]), .I2(bit_ctr[6]), 
            .I3(bit_ctr[19]), .O(n46));
    defparam i18_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1598 (.I0(bit_ctr[13]), .I1(bit_ctr[20]), .I2(bit_ctr[23]), 
            .I3(bit_ctr[16]), .O(n47));
    defparam i19_4_lut_adj_1598.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1599 (.I0(bit_ctr[15]), .I1(bit_ctr[14]), .I2(bit_ctr[21]), 
            .I3(bit_ctr[22]), .O(n45));
    defparam i17_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1600 (.I0(bit_ctr[11]), .I1(bit_ctr[7]), .I2(bit_ctr[17]), 
            .I3(bit_ctr[29]), .O(n44));
    defparam i16_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1601 (.I0(bit_ctr[12]), .I1(bit_ctr[30]), .I2(n36179), 
            .I3(bit_ctr[25]), .O(n43));
    defparam i15_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1602 (.I0(bit_ctr[27]), .I1(bit_ctr[31]), .I2(bit_ctr[10]), 
            .I3(bit_ctr[5]), .O(n49));
    defparam i21_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44), .O(\state_3__N_528[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i467_2_lut (.I0(LED_c), .I1(\state_3__N_528[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n1923));   // verilog/neopixel.v(40[18] 45[12])
    defparam i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_612_i8_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n8));
    defparam equal_612_i8_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 mod_5_add_1473_9_lut (.I0(GND_net), .I1(n2103), .I2(VCC_net), 
            .I3(n42138), .O(n2159[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_9 (.CI(n42138), .I0(n2103), .I1(VCC_net), 
            .CO(n42139));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(GND_net), .I1(n1506), .I2(VCC_net), 
            .I3(n40734), .O(n1565[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_8_lut (.I0(GND_net), .I1(n2104), .I2(VCC_net), 
            .I3(n42137), .O(n2159[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_6 (.CI(n40734), .I0(n1506), .I1(VCC_net), 
            .CO(n40735));
    SB_CARRY mod_5_add_1473_8 (.CI(n42137), .I0(n2104), .I1(VCC_net), 
            .CO(n42138));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(GND_net), .I1(n2105), .I2(VCC_net), 
            .I3(n42136), .O(n2159[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_7 (.CI(n42136), .I0(n2105), .I1(VCC_net), 
            .CO(n42137));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(GND_net), .I1(n2106), .I2(VCC_net), 
            .I3(n42135), .O(n2159[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_6 (.CI(n42135), .I0(n2106), .I1(VCC_net), 
            .CO(n42136));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(GND_net), .I1(n2107), .I2(VCC_net), 
            .I3(n42134), .O(n2159[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_5 (.CI(n42134), .I0(n2107), .I1(VCC_net), 
            .CO(n42135));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(GND_net), .I1(n2108), .I2(VCC_net), 
            .I3(n42133), .O(n2159[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_4 (.CI(n42133), .I0(n2108), .I1(VCC_net), 
            .CO(n42134));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n29362), .I2(VCC_net), 
            .I3(n40555), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(n51314), .I1(n6), .I2(n1923), .I3(\state[1] ), 
            .O(n29446));
    defparam i3_4_lut.LUT_INIT = 16'hc040;
    SB_LUT4 mod_5_add_1473_3_lut (.I0(GND_net), .I1(n2109), .I2(GND_net), 
            .I3(n42132), .O(n2159[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_3 (.CI(n42132), .I0(n2109), .I1(GND_net), 
            .CO(n42133));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(VCC_net), .O(n2159[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(GND_net), 
            .CO(n42132));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2225), .I1(n2192), .I2(VCC_net), 
            .I3(n42131), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(GND_net), .I1(n2193), .I2(VCC_net), 
            .I3(n42130), .O(n2258[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_19 (.CI(n42130), .I0(n2193), .I1(VCC_net), 
            .CO(n42131));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(GND_net), .I1(n2194), .I2(VCC_net), 
            .I3(n42129), .O(n2258[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_18 (.CI(n42129), .I0(n2194), .I1(VCC_net), 
            .CO(n42130));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(GND_net), .I1(n2195), .I2(VCC_net), 
            .I3(n42128), .O(n2258[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_17 (.CI(n42128), .I0(n2195), .I1(VCC_net), 
            .CO(n42129));
    SB_CARRY mod_5_add_669_5 (.CI(n40555), .I0(n29362), .I1(VCC_net), 
            .CO(n40556));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(GND_net), .I1(n2196), .I2(VCC_net), 
            .I3(n42127), .O(n2258[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_5_lut (.I0(GND_net), .I1(n1507), .I2(VCC_net), 
            .I3(n40733), .O(n1565[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_16 (.CI(n42127), .I0(n2196), .I1(VCC_net), 
            .CO(n42128));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n29316), .I2(VCC_net), 
            .I3(n40554), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_15_lut (.I0(GND_net), .I1(n2197), .I2(VCC_net), 
            .I3(n42126), .O(n2258[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n40554), .I0(n29316), .I1(VCC_net), 
            .CO(n40555));
    SB_CARRY mod_5_add_1540_15 (.CI(n42126), .I0(n2197), .I1(VCC_net), 
            .CO(n42127));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(GND_net), .I1(n2198), .I2(VCC_net), 
            .I3(n42125), .O(n2258[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n26353), .I2(GND_net), 
            .I3(n40553), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_14 (.CI(n42125), .I0(n2198), .I1(VCC_net), 
            .CO(n42126));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(GND_net), .I1(n2199), .I2(VCC_net), 
            .I3(n42124), .O(n2258[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_5 (.CI(n40733), .I0(n1507), .I1(VCC_net), 
            .CO(n40734));
    SB_CARRY mod_5_add_1540_13 (.CI(n42124), .I0(n2199), .I1(VCC_net), 
            .CO(n42125));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(GND_net), .I1(n2200), .I2(VCC_net), 
            .I3(n42123), .O(n2258[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_12 (.CI(n42123), .I0(n2200), .I1(VCC_net), 
            .CO(n42124));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(GND_net), .I1(n2201), .I2(VCC_net), 
            .I3(n42122), .O(n2258[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_11 (.CI(n42122), .I0(n2201), .I1(VCC_net), 
            .CO(n42123));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(GND_net), .I1(n2202), .I2(VCC_net), 
            .I3(n42121), .O(n2258[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_10 (.CI(n42121), .I0(n2202), .I1(VCC_net), 
            .CO(n42122));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(GND_net), .I1(n2203), .I2(VCC_net), 
            .I3(n42120), .O(n2258[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_9 (.CI(n42120), .I0(n2203), .I1(VCC_net), 
            .CO(n42121));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(GND_net), .I1(n2204), .I2(VCC_net), 
            .I3(n42119), .O(n2258[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_8 (.CI(n42119), .I0(n2204), .I1(VCC_net), 
            .CO(n42120));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(GND_net), .I1(n2205), .I2(VCC_net), 
            .I3(n42118), .O(n2258[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_7 (.CI(n42118), .I0(n2205), .I1(VCC_net), 
            .CO(n42119));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(GND_net), .I1(n2206), .I2(VCC_net), 
            .I3(n42117), .O(n2258[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_6 (.CI(n42117), .I0(n2206), .I1(VCC_net), 
            .CO(n42118));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(GND_net), .I1(n2207), .I2(VCC_net), 
            .I3(n42116), .O(n2258[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26_4_lut_adj_1603 (.I0(n8), .I1(n51333), .I2(\state[1] ), 
            .I3(n46580), .O(n6801));
    defparam i26_4_lut_adj_1603.LUT_INIT = 16'hc5c0;
    SB_CARRY mod_5_add_1540_5 (.CI(n42116), .I0(n2207), .I1(VCC_net), 
            .CO(n42117));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(GND_net), .I1(n2208), .I2(VCC_net), 
            .I3(n42115), .O(n2258[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_4 (.CI(n42115), .I0(n2208), .I1(VCC_net), 
            .CO(n42116));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(GND_net), .I1(n2209), .I2(GND_net), 
            .I3(n42114), .O(n2258[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_3 (.CI(n42114), .I0(n2209), .I1(GND_net), 
            .CO(n42115));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(VCC_net), .O(n2258[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(GND_net), 
            .CO(n42114));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2324), .I1(n2291), .I2(VCC_net), 
            .I3(n42113), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(GND_net), .I1(n2292), .I2(VCC_net), 
            .I3(n42112), .O(n2357[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_4_lut (.I0(GND_net), .I1(n1508), .I2(VCC_net), 
            .I3(n40732), .O(n1565[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_20 (.CI(n42112), .I0(n2292), .I1(VCC_net), 
            .CO(n42113));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(GND_net), .I1(n2293), .I2(VCC_net), 
            .I3(n42111), .O(n2357[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_19 (.CI(n42111), .I0(n2293), .I1(VCC_net), 
            .CO(n42112));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(GND_net), .I1(n2294), .I2(VCC_net), 
            .I3(n42110), .O(n2357[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_18 (.CI(n42110), .I0(n2294), .I1(VCC_net), 
            .CO(n42111));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(GND_net), .I1(n2295), .I2(VCC_net), 
            .I3(n42109), .O(n2357[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_17 (.CI(n42109), .I0(n2295), .I1(VCC_net), 
            .CO(n42110));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(GND_net), .I1(n2296), .I2(VCC_net), 
            .I3(n42108), .O(n2357[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_16 (.CI(n42108), .I0(n2296), .I1(VCC_net), 
            .CO(n42109));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(GND_net), .I1(n2297), .I2(VCC_net), 
            .I3(n42107), .O(n2357[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_15 (.CI(n42107), .I0(n2297), .I1(VCC_net), 
            .CO(n42108));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(GND_net), .I1(n2298), .I2(VCC_net), 
            .I3(n42106), .O(n2357[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_14 (.CI(n42106), .I0(n2298), .I1(VCC_net), 
            .CO(n42107));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(GND_net), .I1(n2299), .I2(VCC_net), 
            .I3(n42105), .O(n2357[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n40553), .I0(n26353), .I1(GND_net), 
            .CO(n40554));
    SB_CARRY mod_5_add_1607_13 (.CI(n42105), .I0(n2299), .I1(VCC_net), 
            .CO(n42106));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(GND_net), .I1(n2300), .I2(VCC_net), 
            .I3(n42104), .O(n2357[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_12 (.CI(n42104), .I0(n2300), .I1(VCC_net), 
            .CO(n42105));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(GND_net), .I1(n2301), .I2(VCC_net), 
            .I3(n42103), .O(n2357[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_11 (.CI(n42103), .I0(n2301), .I1(VCC_net), 
            .CO(n42104));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(GND_net), .I1(n2302), .I2(VCC_net), 
            .I3(n42102), .O(n2357[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_10 (.CI(n42102), .I0(n2302), .I1(VCC_net), 
            .CO(n42103));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(GND_net), .I1(n2303), .I2(VCC_net), 
            .I3(n42101), .O(n2357[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_9 (.CI(n42101), .I0(n2303), .I1(VCC_net), 
            .CO(n42102));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(GND_net), .I1(n2304), .I2(VCC_net), 
            .I3(n42100), .O(n2357[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_8 (.CI(n42100), .I0(n2304), .I1(VCC_net), 
            .CO(n42101));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(GND_net), .I1(n2305), .I2(VCC_net), 
            .I3(n42099), .O(n2357[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_7 (.CI(n42099), .I0(n2305), .I1(VCC_net), 
            .CO(n42100));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(GND_net), .I1(n2306), .I2(VCC_net), 
            .I3(n42098), .O(n2357[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_6 (.CI(n42098), .I0(n2306), .I1(VCC_net), 
            .CO(n42099));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(GND_net), .I1(n2307), .I2(VCC_net), 
            .I3(n42097), .O(n2357[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_5 (.CI(n42097), .I0(n2307), .I1(VCC_net), 
            .CO(n42098));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(GND_net), .I1(n2308), .I2(VCC_net), 
            .I3(n42096), .O(n2357[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_4 (.CI(n42096), .I0(n2308), .I1(VCC_net), 
            .CO(n42097));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(GND_net), .I1(n2309), .I2(GND_net), 
            .I3(n42095), .O(n2357[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_3 (.CI(n42095), .I0(n2309), .I1(GND_net), 
            .CO(n42096));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(VCC_net), .O(n2357[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(GND_net), 
            .CO(n42095));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2423), .I1(n2390), .I2(VCC_net), 
            .I3(n42094), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(GND_net), .I1(n2391), .I2(VCC_net), 
            .I3(n42093), .O(n2456[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_21 (.CI(n42093), .I0(n2391), .I1(VCC_net), 
            .CO(n42094));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(GND_net), .I1(n2392), .I2(VCC_net), 
            .I3(n42092), .O(n2456[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_20 (.CI(n42092), .I0(n2392), .I1(VCC_net), 
            .CO(n42093));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(GND_net), .I1(n2393), .I2(VCC_net), 
            .I3(n42091), .O(n2456[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_19 (.CI(n42091), .I0(n2393), .I1(VCC_net), 
            .CO(n42092));
    SB_LUT4 i36913_2_lut (.I0(n971[29]), .I1(n2_adj_5049), .I2(GND_net), 
            .I3(GND_net), .O(n52396));   // verilog/neopixel.v(22[26:36])
    defparam i36913_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i36915_2_lut (.I0(n971[30]), .I1(n2_adj_5049), .I2(GND_net), 
            .I3(GND_net), .O(n52398));   // verilog/neopixel.v(22[26:36])
    defparam i36915_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mod_5_i673_3_lut (.I0(n29362), .I1(n971[29]), .I2(n2_adj_5049), 
            .I3(GND_net), .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i673_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2_adj_5049), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n26353), .I1(n971[27]), .I2(n2_adj_5049), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_add_1674_18_lut (.I0(GND_net), .I1(n2394), .I2(VCC_net), 
            .I3(n42090), .O(n2456[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_18 (.CI(n42090), .I0(n2394), .I1(VCC_net), 
            .CO(n42091));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(GND_net), .I1(n2395), .I2(VCC_net), 
            .I3(n42089), .O(n2456[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i674_3_lut (.I0(n29316), .I1(n971[28]), .I2(n2_adj_5049), 
            .I3(GND_net), .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36922_2_lut (.I0(n971[31]), .I1(n2_adj_5049), .I2(GND_net), 
            .I3(GND_net), .O(n52405));   // verilog/neopixel.v(22[26:36])
    defparam i36922_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n7_adj_5050));
    defparam i1_3_lut.LUT_INIT = 16'heaea;
    SB_CARRY mod_5_add_1674_17 (.CI(n42089), .I0(n2395), .I1(VCC_net), 
            .CO(n42090));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(GND_net), .I1(n2396), .I2(VCC_net), 
            .I3(n42088), .O(n2456[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_16 (.CI(n42088), .I0(n2396), .I1(VCC_net), 
            .CO(n42089));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(GND_net), .I1(n2397), .I2(VCC_net), 
            .I3(n42087), .O(n2456[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_4 (.CI(n40732), .I0(n1508), .I1(VCC_net), 
            .CO(n40733));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(GND_net), .I1(n1509), .I2(GND_net), 
            .I3(n40731), .O(n1565[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut_adj_1604 (.I0(n52405), .I1(n7_adj_5050), .I2(n1006), 
            .I3(n8_adj_5051), .O(n1037));
    defparam i5_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n40553));
    SB_CARRY mod_5_add_1071_3 (.CI(n40731), .I0(n1509), .I1(GND_net), 
            .CO(n40732));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(VCC_net), .O(n1565[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_15 (.CI(n42087), .I0(n2397), .I1(VCC_net), 
            .CO(n42088));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(GND_net), .I1(n2398), .I2(VCC_net), 
            .I3(n42086), .O(n2456[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_14 (.CI(n42086), .I0(n2398), .I1(VCC_net), 
            .CO(n42087));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(GND_net), .I1(n2399), .I2(VCC_net), 
            .I3(n42085), .O(n2456[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_13 (.CI(n42085), .I0(n2399), .I1(VCC_net), 
            .CO(n42086));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(GND_net), .I1(n2400), .I2(VCC_net), 
            .I3(n42084), .O(n2456[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_12 (.CI(n42084), .I0(n2400), .I1(VCC_net), 
            .CO(n42085));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(GND_net), .I1(n2401), .I2(VCC_net), 
            .I3(n42083), .O(n2456[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_11 (.CI(n42083), .I0(n2401), .I1(VCC_net), 
            .CO(n42084));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(GND_net), .I1(n2402), .I2(VCC_net), 
            .I3(n42082), .O(n2456[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_10 (.CI(n42082), .I0(n2402), .I1(VCC_net), 
            .CO(n42083));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(GND_net), .I1(n2403), .I2(VCC_net), 
            .I3(n42081), .O(n2456[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_9 (.CI(n42081), .I0(n2403), .I1(VCC_net), 
            .CO(n42082));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(GND_net), .I1(n2404), .I2(VCC_net), 
            .I3(n42080), .O(n2456[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_8 (.CI(n42080), .I0(n2404), .I1(VCC_net), 
            .CO(n42081));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(GND_net), .I1(n2405), .I2(VCC_net), 
            .I3(n42079), .O(n2456[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_7 (.CI(n42079), .I0(n2405), .I1(VCC_net), 
            .CO(n42080));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(GND_net), .I1(n2406), .I2(VCC_net), 
            .I3(n42078), .O(n2456[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_6 (.CI(n42078), .I0(n2406), .I1(VCC_net), 
            .CO(n42079));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(GND_net), .I1(n2407), .I2(VCC_net), 
            .I3(n42077), .O(n2456[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_5 (.CI(n42077), .I0(n2407), .I1(VCC_net), 
            .CO(n42078));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(GND_net), .I1(n2408), .I2(VCC_net), 
            .I3(n42076), .O(n2456[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_4 (.CI(n42076), .I0(n2408), .I1(VCC_net), 
            .CO(n42077));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(GND_net), .I1(n2409), .I2(GND_net), 
            .I3(n42075), .O(n2456[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_3 (.CI(n42075), .I0(n2409), .I1(GND_net), 
            .CO(n42076));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(VCC_net), .O(n2456[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(GND_net), 
            .CO(n42075));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2522), .I1(n2489), .I2(VCC_net), 
            .I3(n42074), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(GND_net), .I1(n2490), .I2(VCC_net), 
            .I3(n42073), .O(n2555[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_22 (.CI(n42073), .I0(n2490), .I1(VCC_net), 
            .CO(n42074));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(GND_net), .I1(n2491), .I2(VCC_net), 
            .I3(n42072), .O(n2555[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_21 (.CI(n42072), .I0(n2491), .I1(VCC_net), 
            .CO(n42073));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(GND_net), .I1(n2492), .I2(VCC_net), 
            .I3(n42071), .O(n2555[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_20 (.CI(n42071), .I0(n2492), .I1(VCC_net), 
            .CO(n42072));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(GND_net), .I1(n2493), .I2(VCC_net), 
            .I3(n42070), .O(n2555[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_19 (.CI(n42070), .I0(n2493), .I1(VCC_net), 
            .CO(n42071));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(GND_net), .I1(n2494), .I2(VCC_net), 
            .I3(n42069), .O(n2555[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_18 (.CI(n42069), .I0(n2494), .I1(VCC_net), 
            .CO(n42070));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(GND_net), .I1(n2495), .I2(VCC_net), 
            .I3(n42068), .O(n2555[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_17 (.CI(n42068), .I0(n2495), .I1(VCC_net), 
            .CO(n42069));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(GND_net), .I1(n2496), .I2(VCC_net), 
            .I3(n42067), .O(n2555[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_16 (.CI(n42067), .I0(n2496), .I1(VCC_net), 
            .CO(n42068));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(GND_net), .I1(n2497), .I2(VCC_net), 
            .I3(n42066), .O(n2555[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_15 (.CI(n42066), .I0(n2497), .I1(VCC_net), 
            .CO(n42067));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(GND_net), .I1(n2498), .I2(VCC_net), 
            .I3(n42065), .O(n2555[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_14 (.CI(n42065), .I0(n2498), .I1(VCC_net), 
            .CO(n42066));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(GND_net), .I1(n2499), .I2(VCC_net), 
            .I3(n42064), .O(n2555[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_13 (.CI(n42064), .I0(n2499), .I1(VCC_net), 
            .CO(n42065));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(GND_net), .I1(n2500), .I2(VCC_net), 
            .I3(n42063), .O(n2555[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_12 (.CI(n42063), .I0(n2500), .I1(VCC_net), 
            .CO(n42064));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(GND_net), .I1(n2501), .I2(VCC_net), 
            .I3(n42062), .O(n2555[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_11 (.CI(n42062), .I0(n2501), .I1(VCC_net), 
            .CO(n42063));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(GND_net), .I1(n2502), .I2(VCC_net), 
            .I3(n42061), .O(n2555[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_10 (.CI(n42061), .I0(n2502), .I1(VCC_net), 
            .CO(n42062));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(GND_net), .I1(n2503), .I2(VCC_net), 
            .I3(n42060), .O(n2555[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_9 (.CI(n42060), .I0(n2503), .I1(VCC_net), 
            .CO(n42061));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(GND_net), .I1(n2504), .I2(VCC_net), 
            .I3(n42059), .O(n2555[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_8 (.CI(n42059), .I0(n2504), .I1(VCC_net), 
            .CO(n42060));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(GND_net), .I1(n2505), .I2(VCC_net), 
            .I3(n42058), .O(n2555[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_7 (.CI(n42058), .I0(n2505), .I1(VCC_net), 
            .CO(n42059));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(GND_net), .I1(n2506), .I2(VCC_net), 
            .I3(n42057), .O(n2555[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_6 (.CI(n42057), .I0(n2506), .I1(VCC_net), 
            .CO(n42058));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(GND_net), .I1(n2507), .I2(VCC_net), 
            .I3(n42056), .O(n2555[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_5 (.CI(n42056), .I0(n2507), .I1(VCC_net), 
            .CO(n42057));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(GND_net), .I1(n2508), .I2(VCC_net), 
            .I3(n42055), .O(n2555[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_4 (.CI(n42055), .I0(n2508), .I1(VCC_net), 
            .CO(n42056));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(GND_net), .I1(n2509), .I2(GND_net), 
            .I3(n42054), .O(n2555[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_3 (.CI(n42054), .I0(n2509), .I1(GND_net), 
            .CO(n42055));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(VCC_net), .O(n2555[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(GND_net), 
            .CO(n42054));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2621), .I1(n2588), .I2(VCC_net), 
            .I3(n42053), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(GND_net), .I1(n2589), .I2(VCC_net), 
            .I3(n42052), .O(n2654[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_23 (.CI(n42052), .I0(n2589), .I1(VCC_net), 
            .CO(n42053));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(GND_net), .I1(n2590), .I2(VCC_net), 
            .I3(n42051), .O(n2654[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_22 (.CI(n42051), .I0(n2590), .I1(VCC_net), 
            .CO(n42052));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(GND_net), .I1(n2591), .I2(VCC_net), 
            .I3(n42050), .O(n2654[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_21 (.CI(n42050), .I0(n2591), .I1(VCC_net), 
            .CO(n42051));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(GND_net), .I1(n2592), .I2(VCC_net), 
            .I3(n42049), .O(n2654[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_20 (.CI(n42049), .I0(n2592), .I1(VCC_net), 
            .CO(n42050));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(GND_net), .I1(n2593), .I2(VCC_net), 
            .I3(n42048), .O(n2654[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_19 (.CI(n42048), .I0(n2593), .I1(VCC_net), 
            .CO(n42049));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(GND_net), .I1(n2594), .I2(VCC_net), 
            .I3(n42047), .O(n2654[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_18 (.CI(n42047), .I0(n2594), .I1(VCC_net), 
            .CO(n42048));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(GND_net), .I1(n2595), .I2(VCC_net), 
            .I3(n42046), .O(n2654[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_17 (.CI(n42046), .I0(n2595), .I1(VCC_net), 
            .CO(n42047));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(GND_net), .I1(n2596), .I2(VCC_net), 
            .I3(n42045), .O(n2654[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_16 (.CI(n42045), .I0(n2596), .I1(VCC_net), 
            .CO(n42046));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(GND_net), .I1(n2597), .I2(VCC_net), 
            .I3(n42044), .O(n2654[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_15 (.CI(n42044), .I0(n2597), .I1(VCC_net), 
            .CO(n42045));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(GND_net), .I1(n2598), .I2(VCC_net), 
            .I3(n42043), .O(n2654[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_14 (.CI(n42043), .I0(n2598), .I1(VCC_net), 
            .CO(n42044));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(GND_net), .I1(n2599), .I2(VCC_net), 
            .I3(n42042), .O(n2654[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_13 (.CI(n42042), .I0(n2599), .I1(VCC_net), 
            .CO(n42043));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(GND_net), .I1(n2600), .I2(VCC_net), 
            .I3(n42041), .O(n2654[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_12 (.CI(n42041), .I0(n2600), .I1(VCC_net), 
            .CO(n42042));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(GND_net), .I1(n2601), .I2(VCC_net), 
            .I3(n42040), .O(n2654[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_11 (.CI(n42040), .I0(n2601), .I1(VCC_net), 
            .CO(n42041));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(GND_net), .I1(n2602), .I2(VCC_net), 
            .I3(n42039), .O(n2654[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_10 (.CI(n42039), .I0(n2602), .I1(VCC_net), 
            .CO(n42040));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(GND_net), .I1(n2603), .I2(VCC_net), 
            .I3(n42038), .O(n2654[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_9 (.CI(n42038), .I0(n2603), .I1(VCC_net), 
            .CO(n42039));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(GND_net), .I1(n2604), .I2(VCC_net), 
            .I3(n42037), .O(n2654[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_8 (.CI(n42037), .I0(n2604), .I1(VCC_net), 
            .CO(n42038));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(GND_net), .I1(n2605), .I2(VCC_net), 
            .I3(n42036), .O(n2654[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_7 (.CI(n42036), .I0(n2605), .I1(VCC_net), 
            .CO(n42037));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(GND_net), .I1(n2606), .I2(VCC_net), 
            .I3(n42035), .O(n2654[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_6 (.CI(n42035), .I0(n2606), .I1(VCC_net), 
            .CO(n42036));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(GND_net), .I1(n2607), .I2(VCC_net), 
            .I3(n42034), .O(n2654[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_5 (.CI(n42034), .I0(n2607), .I1(VCC_net), 
            .CO(n42035));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(GND_net), .I1(n2608), .I2(VCC_net), 
            .I3(n42033), .O(n2654[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_4 (.CI(n42033), .I0(n2608), .I1(VCC_net), 
            .CO(n42034));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(GND_net), .I1(n2609), .I2(GND_net), 
            .I3(n42032), .O(n2654[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_3 (.CI(n42032), .I0(n2609), .I1(GND_net), 
            .CO(n42033));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(VCC_net), .O(n2654[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(GND_net), 
            .CO(n42032));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2720), .I1(n2687), .I2(VCC_net), 
            .I3(n42031), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(GND_net), .I1(n2688), .I2(VCC_net), 
            .I3(n42030), .O(n2753[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_24 (.CI(n42030), .I0(n2688), .I1(VCC_net), 
            .CO(n42031));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(GND_net), .I1(n2689), .I2(VCC_net), 
            .I3(n42029), .O(n2753[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_23 (.CI(n42029), .I0(n2689), .I1(VCC_net), 
            .CO(n42030));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(GND_net), .I1(n2690), .I2(VCC_net), 
            .I3(n42028), .O(n2753[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_22 (.CI(n42028), .I0(n2690), .I1(VCC_net), 
            .CO(n42029));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(GND_net), .I1(n2691), .I2(VCC_net), 
            .I3(n42027), .O(n2753[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_21 (.CI(n42027), .I0(n2691), .I1(VCC_net), 
            .CO(n42028));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(GND_net), .I1(n2692), .I2(VCC_net), 
            .I3(n42026), .O(n2753[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_20 (.CI(n42026), .I0(n2692), .I1(VCC_net), 
            .CO(n42027));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(GND_net), .I1(n2693), .I2(VCC_net), 
            .I3(n42025), .O(n2753[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_19 (.CI(n42025), .I0(n2693), .I1(VCC_net), 
            .CO(n42026));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(GND_net), .I1(n2694), .I2(VCC_net), 
            .I3(n42024), .O(n2753[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_18 (.CI(n42024), .I0(n2694), .I1(VCC_net), 
            .CO(n42025));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(GND_net), .I1(n2695), .I2(VCC_net), 
            .I3(n42023), .O(n2753[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_17 (.CI(n42023), .I0(n2695), .I1(VCC_net), 
            .CO(n42024));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(GND_net), .I1(n2696), .I2(VCC_net), 
            .I3(n42022), .O(n2753[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_16 (.CI(n42022), .I0(n2696), .I1(VCC_net), 
            .CO(n42023));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(GND_net), .I1(n2697), .I2(VCC_net), 
            .I3(n42021), .O(n2753[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_15 (.CI(n42021), .I0(n2697), .I1(VCC_net), 
            .CO(n42022));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(GND_net), .I1(n2698), .I2(VCC_net), 
            .I3(n42020), .O(n2753[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_14 (.CI(n42020), .I0(n2698), .I1(VCC_net), 
            .CO(n42021));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(GND_net), .I1(n2699), .I2(VCC_net), 
            .I3(n42019), .O(n2753[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_13 (.CI(n42019), .I0(n2699), .I1(VCC_net), 
            .CO(n42020));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(GND_net), .I1(n2700), .I2(VCC_net), 
            .I3(n42018), .O(n2753[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_12 (.CI(n42018), .I0(n2700), .I1(VCC_net), 
            .CO(n42019));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(GND_net), .I1(n2701), .I2(VCC_net), 
            .I3(n42017), .O(n2753[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_11 (.CI(n42017), .I0(n2701), .I1(VCC_net), 
            .CO(n42018));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(GND_net), .I1(n2702), .I2(VCC_net), 
            .I3(n42016), .O(n2753[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_10 (.CI(n42016), .I0(n2702), .I1(VCC_net), 
            .CO(n42017));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(GND_net), .I1(n2703), .I2(VCC_net), 
            .I3(n42015), .O(n2753[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_9 (.CI(n42015), .I0(n2703), .I1(VCC_net), 
            .CO(n42016));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(GND_net), .I1(n2704), .I2(VCC_net), 
            .I3(n42014), .O(n2753[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_8 (.CI(n42014), .I0(n2704), .I1(VCC_net), 
            .CO(n42015));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(GND_net), .I1(n2705), .I2(VCC_net), 
            .I3(n42013), .O(n2753[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_7 (.CI(n42013), .I0(n2705), .I1(VCC_net), 
            .CO(n42014));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(GND_net), .I1(n2706), .I2(VCC_net), 
            .I3(n42012), .O(n2753[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_6 (.CI(n42012), .I0(n2706), .I1(VCC_net), 
            .CO(n42013));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(GND_net), .I1(n2707), .I2(VCC_net), 
            .I3(n42011), .O(n2753[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_5 (.CI(n42011), .I0(n2707), .I1(VCC_net), 
            .CO(n42012));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(GND_net), .I1(n2708), .I2(VCC_net), 
            .I3(n42010), .O(n2753[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_4 (.CI(n42010), .I0(n2708), .I1(VCC_net), 
            .CO(n42011));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(GND_net), .I1(n2709), .I2(GND_net), 
            .I3(n42009), .O(n2753[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_3 (.CI(n42009), .I0(n2709), .I1(GND_net), 
            .CO(n42010));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(VCC_net), .O(n2753[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_2058__i1 (.Q(bit_ctr[1]), .C(CLK_c), .E(n6801), 
            .D(n133[1]), .R(n29446));   // verilog/neopixel.v(69[23:32])
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(GND_net), 
            .CO(n42009));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n42008), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n42007), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n42007), .I0(n2787), .I1(n2819), .CO(n42008));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n42006), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n42006), .I0(n2788), .I1(n2819), .CO(n42007));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n42005), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(GND_net), 
            .CO(n40731));
    SB_CARRY mod_5_add_1942_23 (.CI(n42005), .I0(n2789), .I1(n2819), .CO(n42006));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n42004), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n42004), .I0(n2790), .I1(n2819), .CO(n42005));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n42003), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n42003), .I0(n2791), .I1(n2819), .CO(n42004));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n42002), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n42002), .I0(n2792), .I1(n2819), .CO(n42003));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n42001), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n42001), .I0(n2793), .I1(n2819), .CO(n42002));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n42000), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n42000), .I0(n2794), .I1(n2819), .CO(n42001));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n41999), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n41999), .I0(n2795), .I1(n2819), .CO(n42000));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n41998), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n41998), .I0(n2796), .I1(n2819), .CO(n41999));
    SB_DFF timer_2057__i1 (.Q(timer[1]), .C(CLK_c), .D(n133_adj_5095[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i2 (.Q(timer[2]), .C(CLK_c), .D(n133_adj_5095[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i3 (.Q(timer[3]), .C(CLK_c), .D(n133_adj_5095[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i4 (.Q(timer[4]), .C(CLK_c), .D(n133_adj_5095[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i5 (.Q(timer[5]), .C(CLK_c), .D(n133_adj_5095[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i6 (.Q(timer[6]), .C(CLK_c), .D(n133_adj_5095[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i7 (.Q(timer[7]), .C(CLK_c), .D(n133_adj_5095[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i8 (.Q(timer[8]), .C(CLK_c), .D(n133_adj_5095[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i9 (.Q(timer[9]), .C(CLK_c), .D(n133_adj_5095[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i10 (.Q(timer[10]), .C(CLK_c), .D(n133_adj_5095[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i11 (.Q(timer[11]), .C(CLK_c), .D(n133_adj_5095[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i12 (.Q(timer[12]), .C(CLK_c), .D(n133_adj_5095[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i13 (.Q(timer[13]), .C(CLK_c), .D(n133_adj_5095[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i14 (.Q(timer[14]), .C(CLK_c), .D(n133_adj_5095[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i15 (.Q(timer[15]), .C(CLK_c), .D(n133_adj_5095[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i16 (.Q(timer[16]), .C(CLK_c), .D(n133_adj_5095[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i17 (.Q(timer[17]), .C(CLK_c), .D(n133_adj_5095[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i18 (.Q(timer[18]), .C(CLK_c), .D(n133_adj_5095[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i19 (.Q(timer[19]), .C(CLK_c), .D(n133_adj_5095[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i20 (.Q(timer[20]), .C(CLK_c), .D(n133_adj_5095[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i21 (.Q(timer[21]), .C(CLK_c), .D(n133_adj_5095[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i22 (.Q(timer[22]), .C(CLK_c), .D(n133_adj_5095[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i23 (.Q(timer[23]), .C(CLK_c), .D(n133_adj_5095[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i24 (.Q(timer[24]), .C(CLK_c), .D(n133_adj_5095[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i25 (.Q(timer[25]), .C(CLK_c), .D(n133_adj_5095[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i26 (.Q(timer[26]), .C(CLK_c), .D(n133_adj_5095[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i27 (.Q(timer[27]), .C(CLK_c), .D(n133_adj_5095[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i28 (.Q(timer[28]), .C(CLK_c), .D(n133_adj_5095[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i29 (.Q(timer[29]), .C(CLK_c), .D(n133_adj_5095[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i30 (.Q(timer[30]), .C(CLK_c), .D(n133_adj_5095[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i31 (.Q(timer[31]), .C(CLK_c), .D(n133_adj_5095[31]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i37615_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n53098));
    defparam i37615_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n41997), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(CLK_c), .E(VCC_net), .D(n29544));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(CLK_c), .D(n29539));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1942_15 (.CI(n41997), .I0(n2797), .I1(n2819), .CO(n41998));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n41996), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n41996), .I0(n2798), .I1(n2819), .CO(n41997));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n41995), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n41995), .I0(n2799), .I1(n2819), .CO(n41996));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n41994), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n41994), .I0(n2800), .I1(n2819), .CO(n41995));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n41993), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n41993), .I0(n2801), .I1(n2819), .CO(n41994));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n41992), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_10 (.CI(n41992), .I0(n2802), .I1(n2819), .CO(n41993));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n41991), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n41991), .I0(n2803), .I1(n2819), .CO(n41992));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n41990), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n41990), .I0(n2804), .I1(n2819), .CO(n41991));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n41989), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n41989), .I0(n2805), .I1(n2819), .CO(n41990));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n41988), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n41988), .I0(n2806), .I1(n2819), .CO(n41989));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n41987), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n41987), .I0(n2807), .I1(n2819), .CO(n41988));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n41986), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n41986), .I0(n2808), .I1(n2819), .CO(n41987));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n53098), 
            .I3(n41985), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n41985), .I0(n2809), .I1(n53098), .CO(n41986));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n53098), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n53098), 
            .CO(n41985));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n3017), .I1(n2984), .I2(VCC_net), 
            .I3(n41984), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(GND_net), .I1(n2985), .I2(VCC_net), 
            .I3(n41983), .O(n3050[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_27 (.CI(n41983), .I0(n2985), .I1(VCC_net), 
            .CO(n41984));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(GND_net), .I1(n2986), .I2(VCC_net), 
            .I3(n41982), .O(n3050[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_26 (.CI(n41982), .I0(n2986), .I1(VCC_net), 
            .CO(n41983));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(GND_net), .I1(n2987), .I2(VCC_net), 
            .I3(n41981), .O(n3050[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_25 (.CI(n41981), .I0(n2987), .I1(VCC_net), 
            .CO(n41982));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(GND_net), .I1(n2988), .I2(VCC_net), 
            .I3(n41980), .O(n3050[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_24 (.CI(n41980), .I0(n2988), .I1(VCC_net), 
            .CO(n41981));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(GND_net), .I1(n2989), .I2(VCC_net), 
            .I3(n41979), .O(n3050[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_23 (.CI(n41979), .I0(n2989), .I1(VCC_net), 
            .CO(n41980));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(GND_net), .I1(n2990), .I2(VCC_net), 
            .I3(n41978), .O(n3050[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_22 (.CI(n41978), .I0(n2990), .I1(VCC_net), 
            .CO(n41979));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(GND_net), .I1(n2991), .I2(VCC_net), 
            .I3(n41977), .O(n3050[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_21 (.CI(n41977), .I0(n2991), .I1(VCC_net), 
            .CO(n41978));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(GND_net), .I1(n2992), .I2(VCC_net), 
            .I3(n41976), .O(n3050[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_20 (.CI(n41976), .I0(n2992), .I1(VCC_net), 
            .CO(n41977));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(GND_net), .I1(n2993), .I2(VCC_net), 
            .I3(n41975), .O(n3050[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_19 (.CI(n41975), .I0(n2993), .I1(VCC_net), 
            .CO(n41976));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(GND_net), .I1(n2994), .I2(VCC_net), 
            .I3(n41974), .O(n3050[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_18 (.CI(n41974), .I0(n2994), .I1(VCC_net), 
            .CO(n41975));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(GND_net), .I1(n2995), .I2(VCC_net), 
            .I3(n41973), .O(n3050[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_17 (.CI(n41973), .I0(n2995), .I1(VCC_net), 
            .CO(n41974));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(GND_net), .I1(n2996), .I2(VCC_net), 
            .I3(n41972), .O(n3050[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_16 (.CI(n41972), .I0(n2996), .I1(VCC_net), 
            .CO(n41973));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(GND_net), .I1(n2997), .I2(VCC_net), 
            .I3(n41971), .O(n3050[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_15 (.CI(n41971), .I0(n2997), .I1(VCC_net), 
            .CO(n41972));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(GND_net), .I1(n2998), .I2(VCC_net), 
            .I3(n41970), .O(n3050[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_14 (.CI(n41970), .I0(n2998), .I1(VCC_net), 
            .CO(n41971));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(GND_net), .I1(n2999), .I2(VCC_net), 
            .I3(n41969), .O(n3050[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_13 (.CI(n41969), .I0(n2999), .I1(VCC_net), 
            .CO(n41970));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(GND_net), .I1(n3000), .I2(VCC_net), 
            .I3(n41968), .O(n3050[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_12 (.CI(n41968), .I0(n3000), .I1(VCC_net), 
            .CO(n41969));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(GND_net), .I1(n3001), .I2(VCC_net), 
            .I3(n41967), .O(n3050[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_11 (.CI(n41967), .I0(n3001), .I1(VCC_net), 
            .CO(n41968));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(GND_net), .I1(n3002), .I2(VCC_net), 
            .I3(n41966), .O(n3050[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_10 (.CI(n41966), .I0(n3002), .I1(VCC_net), 
            .CO(n41967));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(GND_net), .I1(n3003), .I2(VCC_net), 
            .I3(n41965), .O(n3050[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_9 (.CI(n41965), .I0(n3003), .I1(VCC_net), 
            .CO(n41966));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(GND_net), .I1(n3004), .I2(VCC_net), 
            .I3(n41964), .O(n3050[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_8 (.CI(n41964), .I0(n3004), .I1(VCC_net), 
            .CO(n41965));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(GND_net), .I1(n3005), .I2(VCC_net), 
            .I3(n41963), .O(n3050[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_7 (.CI(n41963), .I0(n3005), .I1(VCC_net), 
            .CO(n41964));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(GND_net), .I1(n3006), .I2(VCC_net), 
            .I3(n41962), .O(n3050[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_6 (.CI(n41962), .I0(n3006), .I1(VCC_net), 
            .CO(n41963));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(GND_net), .I1(n3007), .I2(VCC_net), 
            .I3(n41961), .O(n3050[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_5 (.CI(n41961), .I0(n3007), .I1(VCC_net), 
            .CO(n41962));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(GND_net), .I1(n3008), .I2(VCC_net), 
            .I3(n41960), .O(n3050[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_4 (.CI(n41960), .I0(n3008), .I1(VCC_net), 
            .CO(n41961));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(GND_net), .I1(n32309), .I2(GND_net), 
            .I3(n41959), .O(n3050[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_3 (.CI(n41959), .I0(n32309), .I1(GND_net), 
            .CO(n41960));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(VCC_net), .O(n3050[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(GND_net), 
            .CO(n41959));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3116), .I1(n3083), .I2(VCC_net), 
            .I3(n41958), .O(n50124)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(GND_net), .I1(n3084), .I2(VCC_net), 
            .I3(n41957), .O(n3149[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_28 (.CI(n41957), .I0(n3084), .I1(VCC_net), 
            .CO(n41958));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(GND_net), .I1(n3085), .I2(VCC_net), 
            .I3(n41956), .O(n3149[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_27 (.CI(n41956), .I0(n3085), .I1(VCC_net), 
            .CO(n41957));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(GND_net), .I1(n3086), .I2(VCC_net), 
            .I3(n41955), .O(n3149[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_26 (.CI(n41955), .I0(n3086), .I1(VCC_net), 
            .CO(n41956));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(GND_net), .I1(n3087), .I2(VCC_net), 
            .I3(n41954), .O(n3149[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_25 (.CI(n41954), .I0(n3087), .I1(VCC_net), 
            .CO(n41955));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(GND_net), .I1(n3088), .I2(VCC_net), 
            .I3(n41953), .O(n3149[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_24 (.CI(n41953), .I0(n3088), .I1(VCC_net), 
            .CO(n41954));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(GND_net), .I1(n3089), .I2(VCC_net), 
            .I3(n41952), .O(n3149[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_23 (.CI(n41952), .I0(n3089), .I1(VCC_net), 
            .CO(n41953));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(GND_net), .I1(n3090), .I2(VCC_net), 
            .I3(n41951), .O(n3149[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_22 (.CI(n41951), .I0(n3090), .I1(VCC_net), 
            .CO(n41952));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(GND_net), .I1(n3091), .I2(VCC_net), 
            .I3(n41950), .O(n3149[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_21 (.CI(n41950), .I0(n3091), .I1(VCC_net), 
            .CO(n41951));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(GND_net), .I1(n3092), .I2(VCC_net), 
            .I3(n41949), .O(n3149[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_20 (.CI(n41949), .I0(n3092), .I1(VCC_net), 
            .CO(n41950));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n52405), .I1(n52405), .I2(n1037), 
            .I3(n40547), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_19_lut (.I0(GND_net), .I1(n3093), .I2(VCC_net), 
            .I3(n41948), .O(n3149[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_19 (.CI(n41948), .I0(n3093), .I1(VCC_net), 
            .CO(n41949));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(GND_net), .I1(n3094), .I2(VCC_net), 
            .I3(n41947), .O(n3149[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_18 (.CI(n41947), .I0(n3094), .I1(VCC_net), 
            .CO(n41948));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(GND_net), .I1(n3095), .I2(VCC_net), 
            .I3(n41946), .O(n3149[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_17 (.CI(n41946), .I0(n3095), .I1(VCC_net), 
            .CO(n41947));
    SB_LUT4 mod_5_add_736_7_lut (.I0(n52398), .I1(n52398), .I2(n1037), 
            .I3(n40546), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_16_lut (.I0(GND_net), .I1(n3096), .I2(VCC_net), 
            .I3(n41945), .O(n3149[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_16 (.CI(n41945), .I0(n3096), .I1(VCC_net), 
            .CO(n41946));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(GND_net), .I1(n3097), .I2(VCC_net), 
            .I3(n41944), .O(n3149[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_15 (.CI(n41944), .I0(n3097), .I1(VCC_net), 
            .CO(n41945));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(GND_net), .I1(n3098), .I2(VCC_net), 
            .I3(n41943), .O(n3149[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_14 (.CI(n41943), .I0(n3098), .I1(VCC_net), 
            .CO(n41944));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(GND_net), .I1(n3099), .I2(VCC_net), 
            .I3(n41942), .O(n3149[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_13 (.CI(n41942), .I0(n3099), .I1(VCC_net), 
            .CO(n41943));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(GND_net), .I1(n3100), .I2(VCC_net), 
            .I3(n41941), .O(n3149[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_12 (.CI(n41941), .I0(n3100), .I1(VCC_net), 
            .CO(n41942));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(GND_net), .I1(n3101), .I2(VCC_net), 
            .I3(n41940), .O(n3149[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_11 (.CI(n41940), .I0(n3101), .I1(VCC_net), 
            .CO(n41941));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(GND_net), .I1(n3102), .I2(VCC_net), 
            .I3(n41939), .O(n3149[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_10 (.CI(n41939), .I0(n3102), .I1(VCC_net), 
            .CO(n41940));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(GND_net), .I1(n3103), .I2(VCC_net), 
            .I3(n41938), .O(n3149[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_9 (.CI(n41938), .I0(n3103), .I1(VCC_net), 
            .CO(n41939));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(GND_net), .I1(n3104), .I2(VCC_net), 
            .I3(n41937), .O(n3149[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_736_7 (.CI(n40546), .I0(n52398), .I1(n1037), .CO(n40547));
    SB_CARRY mod_5_add_2143_8 (.CI(n41937), .I0(n3104), .I1(VCC_net), 
            .CO(n41938));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(GND_net), .I1(n3105), .I2(VCC_net), 
            .I3(n41936), .O(n3149[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_7 (.CI(n41936), .I0(n3105), .I1(VCC_net), 
            .CO(n41937));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(GND_net), .I1(n3106), .I2(VCC_net), 
            .I3(n41935), .O(n3149[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_6 (.CI(n41935), .I0(n3106), .I1(VCC_net), 
            .CO(n41936));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(GND_net), .I1(n3107), .I2(VCC_net), 
            .I3(n41934), .O(n3149[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_5 (.CI(n41934), .I0(n3107), .I1(VCC_net), 
            .CO(n41935));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(GND_net), .I1(n3108), .I2(VCC_net), 
            .I3(n41933), .O(n3149[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_736_6_lut (.I0(n52396), .I1(n1006), .I2(n1037), 
            .I3(n40545), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n41933), .I0(n3108), .I1(VCC_net), 
            .CO(n41934));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(GND_net), .I1(n3109), .I2(GND_net), 
            .I3(n41932), .O(n3149[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_3 (.CI(n41932), .I0(n3109), .I1(GND_net), 
            .CO(n41933));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(VCC_net), .O(n3149[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(GND_net), 
            .CO(n41932));
    SB_CARRY mod_5_add_736_6 (.CI(n40545), .I0(n1006), .I1(n1037), .CO(n40546));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n52397), .I1(n1007), .I2(n1037), 
            .I3(n40544), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n40544), .I0(n1007), .I1(n1037), .CO(n40545));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n40543), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n40543), .I0(n1008), .I1(n1037), .CO(n40544));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n53099), 
            .I3(n40542), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n40542), .I0(n1009), .I1(n53099), .CO(n40543));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n53099), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n53099), 
            .CO(n40542));
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(CLK_c), .E(n46623), .D(\neo_pixel_transmitter.done_N_742 ), 
            .R(n48491));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i606_3_lut_3_lut_4_lut_3_lut (.I0(bit_ctr[27]), .I1(n26355), 
            .I2(n29324), .I3(GND_net), .O(n29362));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_3_lut_4_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(bit_ctr[27]), .I1(n26355), .I2(n29324), 
            .I3(GND_net), .O(n26353));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'h8585;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36199_3_lut_4_lut_3_lut (.I0(bit_ctr[27]), .I1(n26355), .I2(n29324), 
            .I3(GND_net), .O(n29316));   // verilog/neopixel.v(22[26:36])
    defparam i36199_3_lut_4_lut_3_lut.LUT_INIT = 16'h1919;
    SB_LUT4 i1_4_lut_4_lut (.I0(bit_ctr[26]), .I1(n26353), .I2(n29362), 
            .I3(n29316), .O(n2_adj_5049));   // verilog/neopixel.v(22[26:36])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i947_3_lut (.I0(n1309), .I1(n1367[23]), .I2(n1334), 
            .I3(GND_net), .O(n1408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i945_3_lut (.I0(n1307), .I1(n1367[25]), .I2(n1334), 
            .I3(GND_net), .O(n1406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i941_3_lut (.I0(n1303), .I1(n1367[29]), .I2(n1334), 
            .I3(GND_net), .O(n1402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i944_3_lut (.I0(n1306), .I1(n1367[26]), .I2(n1334), 
            .I3(GND_net), .O(n1405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i942_3_lut (.I0(n1304), .I1(n1367[28]), .I2(n1334), 
            .I3(GND_net), .O(n1403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i946_3_lut (.I0(n1308), .I1(n1367[24]), .I2(n1334), 
            .I3(GND_net), .O(n1407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i948_3_lut (.I0(bit_ctr[22]), .I1(n1367[22]), .I2(n1334), 
            .I3(GND_net), .O(n1409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i940_3_lut (.I0(n1302), .I1(n1367[30]), .I2(n1334), 
            .I3(GND_net), .O(n1401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i943_3_lut (.I0(n1305), .I1(n1367[27]), .I2(n1334), 
            .I3(GND_net), .O(n1404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_adj_1605 (.I0(n1404), .I1(n1401), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_5052));   // verilog/neopixel.v(22[26:36])
    defparam i2_2_lut_adj_1605.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1606 (.I0(bit_ctr[21]), .I1(n12_adj_5052), .I2(n1400), 
            .I3(n1409), .O(n16_adj_5053));   // verilog/neopixel.v(22[26:36])
    defparam i6_4_lut_adj_1606.LUT_INIT = 16'hfefc;
    SB_LUT4 i7_4_lut_adj_1607 (.I0(n1407), .I1(n1403), .I2(n1405), .I3(n1402), 
            .O(n17_adj_5054));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1608 (.I0(n17_adj_5054), .I1(n1406), .I2(n16_adj_5053), 
            .I3(n1408), .O(n1433));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_3_lut_adj_1609 (.I0(n1007), .I1(n971[30]), .I2(n2_adj_5049), 
            .I3(GND_net), .O(n8_adj_5051));
    defparam i2_2_lut_3_lut_adj_1609.LUT_INIT = 16'haeae;
    SB_LUT4 i35988_2_lut_3_lut (.I0(LED_c), .I1(\state_3__N_528[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n51333));
    defparam i35988_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i35983_3_lut_4_lut (.I0(n27768), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(n4), .O(n51314));
    defparam i35983_3_lut_4_lut.LUT_INIT = 16'hf3f7;
    SB_LUT4 i18798_3_lut (.I0(n32309), .I1(n3050[6]), .I2(n3017), .I3(GND_net), 
            .O(n3108));
    defparam i18798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2092_3_lut (.I0(n2998), .I1(n3050[17]), .I2(n3017), 
            .I3(GND_net), .O(n3097));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2093_3_lut (.I0(n2999), .I1(n3050[16]), .I2(n3017), 
            .I3(GND_net), .O(n3098));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2099_3_lut (.I0(n3005), .I1(n3050[10]), .I2(n3017), 
            .I3(GND_net), .O(n3104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2089_3_lut (.I0(n2995), .I1(n3050[20]), .I2(n3017), 
            .I3(GND_net), .O(n3094));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2088_3_lut (.I0(n2994), .I1(n3050[21]), .I2(n3017), 
            .I3(GND_net), .O(n3093));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2079_3_lut (.I0(n2985), .I1(n3050[30]), .I2(n3017), 
            .I3(GND_net), .O(n3084));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2096_3_lut (.I0(n3002), .I1(n3050[13]), .I2(n3017), 
            .I3(GND_net), .O(n3101));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2101_3_lut (.I0(n3007), .I1(n3050[8]), .I2(n3017), 
            .I3(GND_net), .O(n3106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2102_3_lut (.I0(n3008), .I1(n3050[7]), .I2(n3017), 
            .I3(GND_net), .O(n3107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2087_3_lut (.I0(n2993), .I1(n3050[22]), .I2(n3017), 
            .I3(GND_net), .O(n3092));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2085_3_lut (.I0(n2991), .I1(n3050[24]), .I2(n3017), 
            .I3(GND_net), .O(n3090));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2086_3_lut (.I0(n2992), .I1(n3050[23]), .I2(n3017), 
            .I3(GND_net), .O(n3091));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2084_3_lut (.I0(n2990), .I1(n3050[25]), .I2(n3017), 
            .I3(GND_net), .O(n3089));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18817_3_lut (.I0(bit_ctr[5]), .I1(n3050[5]), .I2(n3017), 
            .I3(GND_net), .O(n3109));
    defparam i18817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2094_3_lut (.I0(n3000), .I1(n3050[15]), .I2(n3017), 
            .I3(GND_net), .O(n3099));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2083_3_lut (.I0(n2989), .I1(n3050[26]), .I2(n3017), 
            .I3(GND_net), .O(n3088));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2081_3_lut (.I0(n2987), .I1(n3050[28]), .I2(n3017), 
            .I3(GND_net), .O(n3086));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2082_3_lut (.I0(n2988), .I1(n3050[27]), .I2(n3017), 
            .I3(GND_net), .O(n3087));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2080_3_lut (.I0(n2986), .I1(n3050[29]), .I2(n3017), 
            .I3(GND_net), .O(n3085));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2091_3_lut (.I0(n2997), .I1(n3050[18]), .I2(n3017), 
            .I3(GND_net), .O(n3096));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2098_3_lut (.I0(n3004), .I1(n3050[11]), .I2(n3017), 
            .I3(GND_net), .O(n3103));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2090_3_lut (.I0(n2996), .I1(n3050[19]), .I2(n3017), 
            .I3(GND_net), .O(n3095));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2026_3_lut (.I0(n2900), .I1(n2951[16]), .I2(n2918), 
            .I3(GND_net), .O(n2999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2034_3_lut (.I0(n2908), .I1(n2951[8]), .I2(n2918), 
            .I3(GND_net), .O(n3007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2018_3_lut (.I0(n2892), .I1(n2951[24]), .I2(n2918), 
            .I3(GND_net), .O(n2991));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2016_3_lut (.I0(n2890), .I1(n2951[26]), .I2(n2918), 
            .I3(GND_net), .O(n2989));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2017_3_lut (.I0(n2891), .I1(n2951[25]), .I2(n2918), 
            .I3(GND_net), .O(n2990));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2015_3_lut (.I0(n2889), .I1(n2951[27]), .I2(n2918), 
            .I3(GND_net), .O(n2988));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2025_3_lut (.I0(n2899), .I1(n2951[17]), .I2(n2918), 
            .I3(GND_net), .O(n2998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2028_3_lut (.I0(n2902), .I1(n2951[14]), .I2(n2918), 
            .I3(GND_net), .O(n3001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2023_3_lut (.I0(n2897), .I1(n2951[19]), .I2(n2918), 
            .I3(GND_net), .O(n2996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2030_3_lut (.I0(n2904), .I1(n2951[12]), .I2(n2918), 
            .I3(GND_net), .O(n3003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2032_3_lut (.I0(n2906), .I1(n2951[10]), .I2(n2918), 
            .I3(GND_net), .O(n3005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2021_3_lut (.I0(n2895), .I1(n2951[21]), .I2(n2918), 
            .I3(GND_net), .O(n2994));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2020_3_lut (.I0(n2894), .I1(n2951[22]), .I2(n2918), 
            .I3(GND_net), .O(n2993));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2027_3_lut (.I0(n2901), .I1(n2951[15]), .I2(n2918), 
            .I3(GND_net), .O(n3000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2019_3_lut (.I0(n2893), .I1(n2951[23]), .I2(n2918), 
            .I3(GND_net), .O(n2992));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18797_3_lut (.I0(bit_ctr[6]), .I1(n2951[6]), .I2(n2918), 
            .I3(GND_net), .O(n32309));
    defparam i18797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2022_3_lut (.I0(n2896), .I1(n2951[20]), .I2(n2918), 
            .I3(GND_net), .O(n2995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2024_3_lut (.I0(n2898), .I1(n2951[18]), .I2(n2918), 
            .I3(GND_net), .O(n2997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2029_3_lut (.I0(n2903), .I1(n2951[13]), .I2(n2918), 
            .I3(GND_net), .O(n3002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2035_3_lut (.I0(n2909), .I1(n2951[7]), .I2(n2918), 
            .I3(GND_net), .O(n3008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36342_3_lut_4_lut (.I0(n27768), .I1(n51824), .I2(start), 
            .I3(\state[1] ), .O(n51825));
    defparam i36342_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35981_2_lut_3_lut (.I0(one_wire_N_679[2]), .I1(one_wire_N_679[3]), 
            .I2(start), .I3(GND_net), .O(n51330));
    defparam i35981_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_i2031_3_lut (.I0(n2905), .I1(n2951[11]), .I2(n2918), 
            .I3(GND_net), .O(n3004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_3_lut_adj_1610 (.I0(n2896), .I1(bit_ctr[6]), .I2(n2909), 
            .I3(GND_net), .O(n32_adj_5055));
    defparam i7_3_lut_adj_1610.LUT_INIT = 16'heaea;
    SB_LUT4 i17_4_lut_adj_1611 (.I0(n2898), .I1(n2899), .I2(n2902), .I3(n2908), 
            .O(n42_adj_5056));
    defparam i17_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2886), .I2(n2885), .I3(GND_net), 
            .O(n38_adj_5057));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n36444), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n48491));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i18_4_lut_adj_1612 (.I0(n2905), .I1(n2904), .I2(n2907), .I3(n2897), 
            .O(n43_adj_5058));
    defparam i18_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1613 (.I0(n2891), .I1(n2893), .I2(n2892), .I3(n2894), 
            .O(n40_adj_5059));
    defparam i15_4_lut_adj_1613.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1614 (.I0(n2895), .I1(n42_adj_5056), .I2(n32_adj_5055), 
            .I3(n2903), .O(n46_adj_5060));
    defparam i21_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1615 (.I0(n2887), .I1(n2889), .I2(n2888), .I3(n2890), 
            .O(n39_adj_5061));
    defparam i14_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1616 (.I0(n43_adj_5058), .I1(n2900), .I2(n38_adj_5057), 
            .I3(n2901), .O(n47_adj_5062));
    defparam i22_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47_adj_5062), .I1(n39_adj_5061), .I2(n46_adj_5060), 
            .I3(n40_adj_5059), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2014_3_lut (.I0(n2888), .I1(n2951[28]), .I2(n2918), 
            .I3(GND_net), .O(n2987));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2013_3_lut (.I0(n2887), .I1(n2951[29]), .I2(n2918), 
            .I3(GND_net), .O(n2986));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2012_3_lut (.I0(n2886), .I1(n2951[30]), .I2(n2918), 
            .I3(GND_net), .O(n2985));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut_adj_1617 (.I0(n3004), .I1(n3008), .I2(n3002), .I3(n2997), 
            .O(n44_adj_5063));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1618 (.I0(bit_ctr[5]), .I1(n2995), .I2(n32309), 
            .I3(GND_net), .O(n33_adj_5064));   // verilog/neopixel.v(22[26:36])
    defparam i7_3_lut_adj_1618.LUT_INIT = 16'hecec;
    SB_LUT4 i14_4_lut_adj_1619 (.I0(n2985), .I1(n2986), .I2(n2984), .I3(n2987), 
            .O(n40_adj_5065));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1619.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1620 (.I0(n3005), .I1(n3003), .I2(n2996), .I3(n3006), 
            .O(n45_adj_5066));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1621 (.I0(n2992), .I1(n3000), .I2(n2993), .I3(n2994), 
            .O(n42_adj_5067));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1622 (.I0(n33_adj_5064), .I1(n44_adj_5063), .I2(n3001), 
            .I3(n2998), .O(n48_adj_5068));   // verilog/neopixel.v(22[26:36])
    defparam i22_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1623 (.I0(n2988), .I1(n2990), .I2(n2989), .I3(n2991), 
            .O(n41_adj_5069));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n45_adj_5066), .I1(n3007), .I2(n40_adj_5065), 
            .I3(n2999), .O(n49_adj_5070));   // verilog/neopixel.v(22[26:36])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n49_adj_5070), .I1(n41_adj_5069), .I2(n48_adj_5068), 
            .I3(n42_adj_5067), .O(n3017));   // verilog/neopixel.v(22[26:36])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2033_3_lut (.I0(n2907), .I1(n2951[9]), .I2(n2918), 
            .I3(GND_net), .O(n3006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2100_3_lut (.I0(n3006), .I1(n3050[9]), .I2(n3017), 
            .I3(GND_net), .O(n3105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2097_3_lut (.I0(n3003), .I1(n3050[12]), .I2(n3017), 
            .I3(GND_net), .O(n3102));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_2_lut (.I0(n3102), .I1(n3105), .I2(GND_net), .I3(GND_net), 
            .O(n36_adj_5071));
    defparam i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19_4_lut_adj_1624 (.I0(n3095), .I1(n3103), .I2(n3096), .I3(n3100), 
            .O(n46_adj_5072));
    defparam i19_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1625 (.I0(n3085), .I1(n3087), .I2(n3086), .I3(n3088), 
            .O(n42_adj_5073));
    defparam i15_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1626 (.I0(n3099), .I1(bit_ctr[4]), .I2(n3109), 
            .I3(GND_net), .O(n34_adj_5074));
    defparam i7_3_lut_adj_1626.LUT_INIT = 16'heaea;
    SB_LUT4 i16_4_lut_adj_1627 (.I0(n3089), .I1(n3091), .I2(n3090), .I3(n3092), 
            .O(n43_adj_5075));
    defparam i16_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1899_3_lut (.I0(n2709), .I1(n2753[9]), .I2(n2720), 
            .I3(GND_net), .O(n2808));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1882_3_lut (.I0(n2692), .I1(n2753[26]), .I2(n2720), 
            .I3(GND_net), .O(n2791));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1898_3_lut (.I0(n2708), .I1(n2753[10]), .I2(n2720), 
            .I3(GND_net), .O(n2807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1892_3_lut (.I0(n2702), .I1(n2753[16]), .I2(n2720), 
            .I3(GND_net), .O(n2801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23_4_lut_adj_1628 (.I0(n3107), .I1(n46_adj_5072), .I2(n36_adj_5071), 
            .I3(n3106), .O(n50));
    defparam i23_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1629 (.I0(n3101), .I1(n42_adj_5073), .I2(n3084), 
            .I3(n3083), .O(n48_adj_5076));
    defparam i21_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1630 (.I0(n43_adj_5075), .I1(n3093), .I2(n34_adj_5074), 
            .I3(n3094), .O(n49_adj_5077));
    defparam i22_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1631 (.I0(n3104), .I1(n3098), .I2(n3097), .I3(n3108), 
            .O(n47_adj_5078));
    defparam i20_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1632 (.I0(n47_adj_5078), .I1(n49_adj_5077), .I2(n48_adj_5076), 
            .I3(n50), .O(n3116));
    defparam i26_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2095_3_lut (.I0(n3001), .I1(n3050[14]), .I2(n3017), 
            .I3(GND_net), .O(n3100));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2162_3_lut (.I0(n3100), .I1(n3149[14]), .I2(n3116), 
            .I3(GND_net), .O(n29_adj_5079));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1888_3_lut (.I0(n2698), .I1(n2753[20]), .I2(n2720), 
            .I3(GND_net), .O(n2797));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2171_3_lut (.I0(n3109), .I1(n3149[5]), .I2(n3116), 
            .I3(GND_net), .O(n11_adj_5080));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1885_3_lut (.I0(n2695), .I1(n2753[23]), .I2(n2720), 
            .I3(GND_net), .O(n2794));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2167_3_lut (.I0(n3105), .I1(n3149[9]), .I2(n3116), 
            .I3(GND_net), .O(n19_adj_5081));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1893_3_lut (.I0(n2703), .I1(n2753[15]), .I2(n2720), 
            .I3(GND_net), .O(n2802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1886_3_lut (.I0(n2696), .I1(n2753[22]), .I2(n2720), 
            .I3(GND_net), .O(n2795));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1891_3_lut (.I0(n2701), .I1(n2753[17]), .I2(n2720), 
            .I3(GND_net), .O(n2800));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2163_3_lut (.I0(n3101), .I1(n3149[13]), .I2(n3116), 
            .I3(GND_net), .O(n27_adj_5082));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2165_3_lut (.I0(n3103), .I1(n3149[11]), .I2(n3116), 
            .I3(GND_net), .O(n23_adj_5083));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1890_3_lut (.I0(n2700), .I1(n2753[18]), .I2(n2720), 
            .I3(GND_net), .O(n2799));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2169_3_lut (.I0(n3107), .I1(n3149[7]), .I2(n3116), 
            .I3(GND_net), .O(n15_adj_5084));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1895_3_lut (.I0(n2705), .I1(n2753[13]), .I2(n2720), 
            .I3(GND_net), .O(n2804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1633 (.I0(n3102), .I1(n29_adj_5079), .I2(n3149[12]), 
            .I3(n3116), .O(n49547));
    defparam i1_4_lut_adj_1633.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1634 (.I0(n3098), .I1(n15_adj_5084), .I2(n3149[16]), 
            .I3(n3116), .O(n49549));
    defparam i1_4_lut_adj_1634.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1635 (.I0(n3096), .I1(n23_adj_5083), .I2(n3149[18]), 
            .I3(n3116), .O(n49543));
    defparam i1_4_lut_adj_1635.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1636 (.I0(n3108), .I1(n27_adj_5082), .I2(n3149[6]), 
            .I3(n3116), .O(n49541));
    defparam i1_4_lut_adj_1636.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2161_3_lut (.I0(n3099), .I1(n3149[15]), .I2(n3116), 
            .I3(GND_net), .O(n31_adj_5085));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1637 (.I0(n3106), .I1(n11_adj_5080), .I2(n3149[8]), 
            .I3(n3116), .O(n49539));
    defparam i1_4_lut_adj_1637.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1638 (.I0(n3104), .I1(n19_adj_5081), .I2(n3149[10]), 
            .I3(n3116), .O(n49551));
    defparam i1_4_lut_adj_1638.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1639 (.I0(n3097), .I1(n31_adj_5085), .I2(n3149[17]), 
            .I3(n3116), .O(n49545));
    defparam i1_4_lut_adj_1639.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2157_3_lut (.I0(n3095), .I1(n3149[19]), .I2(n3116), 
            .I3(GND_net), .O(n39_adj_5086));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1640 (.I0(n39_adj_5086), .I1(n49545), .I2(n49551), 
            .I3(n49539), .O(n49563));
    defparam i1_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1641 (.I0(n49541), .I1(n49543), .I2(n49549), 
            .I3(n49547), .O(n49561));
    defparam i1_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1642 (.I0(n49561), .I1(n49563), .I2(bit_ctr[3]), 
            .I3(n3209), .O(n49567));
    defparam i1_4_lut_adj_1642.LUT_INIT = 16'hfeee;
    SB_LUT4 mod_5_i1883_3_lut (.I0(n2693), .I1(n2753[25]), .I2(n2720), 
            .I3(GND_net), .O(n2792));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1879_3_lut (.I0(n2689), .I1(n2753[29]), .I2(n2720), 
            .I3(GND_net), .O(n2788));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1881_3_lut (.I0(n2691), .I1(n2753[27]), .I2(n2720), 
            .I3(GND_net), .O(n2790));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1643 (.I0(n49567), .I1(n3094), .I2(n3149[20]), 
            .I3(n3116), .O(n49569));
    defparam i1_4_lut_adj_1643.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1644 (.I0(n3093), .I1(n49569), .I2(n3149[21]), 
            .I3(n3116), .O(n49571));
    defparam i1_4_lut_adj_1644.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1645 (.I0(n3092), .I1(n49571), .I2(n3149[22]), 
            .I3(n3116), .O(n49573));
    defparam i1_4_lut_adj_1645.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i1894_3_lut (.I0(n2704), .I1(n2753[14]), .I2(n2720), 
            .I3(GND_net), .O(n2803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(n3091), .I1(n49573), .I2(n3149[23]), 
            .I3(n3116), .O(n49575));
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1647 (.I0(n3090), .I1(n49575), .I2(n3149[24]), 
            .I3(n3116), .O(n49577));
    defparam i1_4_lut_adj_1647.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1648 (.I0(n3089), .I1(n49577), .I2(n3149[25]), 
            .I3(n3116), .O(n49579));
    defparam i1_4_lut_adj_1648.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1649 (.I0(n3088), .I1(n49579), .I2(n3149[26]), 
            .I3(n3116), .O(n49581));
    defparam i1_4_lut_adj_1649.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i1897_3_lut (.I0(n2707), .I1(n2753[11]), .I2(n2720), 
            .I3(GND_net), .O(n2806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1884_3_lut (.I0(n2694), .I1(n2753[24]), .I2(n2720), 
            .I3(GND_net), .O(n2793));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1650 (.I0(n3087), .I1(n49581), .I2(n3149[27]), 
            .I3(n3116), .O(n49583));
    defparam i1_4_lut_adj_1650.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(n3086), .I1(n49583), .I2(n3149[28]), 
            .I3(n3116), .O(n49585));
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2147_3_lut (.I0(n3085), .I1(n3149[29]), .I2(n3116), 
            .I3(GND_net), .O(n59));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2146_3_lut (.I0(n3084), .I1(n3149[30]), .I2(n3116), 
            .I3(GND_net), .O(n61));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1889_3_lut (.I0(n2699), .I1(n2753[19]), .I2(n2720), 
            .I3(GND_net), .O(n2798));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1878_3_lut (.I0(n2688), .I1(n2753[30]), .I2(n2720), 
            .I3(GND_net), .O(n2787));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1896_3_lut (.I0(n2706), .I1(n2753[12]), .I2(n2720), 
            .I3(GND_net), .O(n2805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1880_3_lut (.I0(n2690), .I1(n2753[28]), .I2(n2720), 
            .I3(GND_net), .O(n2789));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1652 (.I0(n61), .I1(n50124), .I2(n59), .I3(n49585), 
            .O(n42492));
    defparam i1_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2172_3_lut (.I0(bit_ctr[4]), .I1(n3149[4]), .I2(n3116), 
            .I3(GND_net), .O(n3209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(\state[1] ), .I1(n36444), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n48405));
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'hf5fd;
    SB_LUT4 i1_4_lut_adj_1654 (.I0(n48405), .I1(n46580), .I2(\state[1] ), 
            .I3(n8), .O(n29252));
    defparam i1_4_lut_adj_1654.LUT_INIT = 16'ha0a8;
    SB_LUT4 i36182_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n42492), .I3(GND_net), 
            .O(color_bit_N_722[4]));
    defparam i36182_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i36349_3_lut (.I0(n53170), .I1(bit_ctr[3]), .I2(n42492), .I3(GND_net), 
            .O(n51343));
    defparam i36349_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i36786_4_lut (.I0(n53110), .I1(n53212), .I2(bit_ctr[3]), .I3(n42492), 
            .O(n52269));   // verilog/neopixel.v(22[26:36])
    defparam i36786_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 mod_5_i1900_3_lut (.I0(bit_ctr[8]), .I1(n2753[8]), .I2(n2720), 
            .I3(GND_net), .O(n2809));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1887_3_lut (.I0(n2697), .I1(n2753[21]), .I2(n2720), 
            .I3(GND_net), .O(n2796));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_3_lut_adj_1655 (.I0(bit_ctr[7]), .I1(n2796), .I2(n2809), 
            .I3(GND_net), .O(n31_adj_5087));
    defparam i7_3_lut_adj_1655.LUT_INIT = 16'hecec;
    SB_LUT4 i21765_4_lut (.I0(n52269), .I1(\state_3__N_528[1] ), .I2(n51343), 
            .I3(color_bit_N_722[4]), .O(state_3__N_528[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i21765_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i15_4_lut_adj_1656 (.I0(n2787), .I1(n2798), .I2(n2793), .I3(n2806), 
            .O(n39_adj_5088));
    defparam i15_4_lut_adj_1656.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1657 (.I0(n2789), .I1(n2805), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_5089));
    defparam i2_2_lut_adj_1657.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1658 (.I0(n2803), .I1(n2790), .I2(n2788), .I3(n2792), 
            .O(n38_adj_5090));
    defparam i14_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20_4_lut_adj_1659 (.I0(n39_adj_5088), .I1(n31_adj_5087), .I2(n2802), 
            .I3(n2794), .O(n44_adj_5091));
    defparam i20_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1660 (.I0(n2804), .I1(n2799), .I2(n2800), .I3(n2795), 
            .O(n42_adj_5092));
    defparam i18_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19_4_lut_adj_1661 (.I0(n2791), .I1(n38_adj_5090), .I2(n26_adj_5089), 
            .I3(n2808), .O(n43_adj_5093));
    defparam i19_4_lut_adj_1661.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1662 (.I0(n2797), .I1(n2801), .I2(n2786), .I3(n2807), 
            .O(n41_adj_5094));
    defparam i17_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1663 (.I0(n41_adj_5094), .I1(n43_adj_5093), .I2(n42_adj_5092), 
            .I3(n44_adj_5091), .O(n2819));
    defparam i23_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18814_3_lut_4_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[28]), .O(n29324));   // verilog/neopixel.v(18[12:19])
    defparam i18814_3_lut_4_lut.LUT_INIT = 16'hdb6d;
    SB_LUT4 i18816_3_lut_4_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[28]), .O(n26355));   // verilog/neopixel.v(18[12:19])
    defparam i18816_3_lut_4_lut.LUT_INIT = 16'hb6db;
    SB_LUT4 bit_ctr_1__bdd_4_lut_37673 (.I0(bit_ctr[1]), .I1(n50400), .I2(n50401), 
            .I3(bit_ctr[2]), .O(n53107));
    defparam bit_ctr_1__bdd_4_lut_37673.LUT_INIT = 16'he4aa;
    SB_LUT4 n53107_bdd_4_lut (.I0(n53107), .I1(n50398), .I2(n50397), .I3(bit_ctr[2]), 
            .O(n53110));
    defparam n53107_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=51, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, setpoint, motor_state, \Ki[11] , \Ki[14] , 
            \Ki[12] , \Ki[3] , \Ki[4] , \Ki[15] , \Kp[1] , \Kp[0] , 
            \Kp[2] , \Ki[5] , \Ki[13] , \Ki[0] , \Ki[1] , \Ki[6] , 
            \Ki[2] , \Kp[3] , \Kp[4] , \Kp[5] , \Kp[6] , IntegralLimit, 
            \Kp[7] , duty, clk32MHz, \Ki[7] , \Ki[8] , \Ki[9] , 
            \Ki[10] , VCC_net, PWMLimit, \Kp[8] , \Kp[9] , \Kp[10] , 
            \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , \Kp[15] ) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    input \Ki[11] ;
    input \Ki[14] ;
    input \Ki[12] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[15] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Ki[5] ;
    input \Ki[13] ;
    input \Ki[0] ;
    input \Ki[1] ;
    input \Ki[6] ;
    input \Ki[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input [23:0]IntegralLimit;
    input \Kp[7] ;
    output [23:0]duty;
    input clk32MHz;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input VCC_net;
    input [23:0]PWMLimit;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [12:0]n18193;
    wire [11:0]n18557;
    
    wire n177, n40805;
    wire [8:0]n19353;
    
    wire n47, n116, n40806, n40714;
    wire [7:0]n19533;
    wire [6:0]n19677;
    
    wire n630, n40713, n41005;
    wire [20:0]n11990;
    
    wire n41006, n35, n104, n40620, n40621, n40535;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    wire [23:0]n4096;
    
    wire n40536, n557, n40712;
    wire [23:0]n1;
    
    wire n40619;
    wire [21:0]n10300;
    
    wire n41004;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3672 ;
    
    wire n40534, n40618, n484, n40711;
    wire [10:0]n18869;
    
    wire n910, n40804, n40617, n837, n40803, n411, n40710, n41003, 
        n40616, n40533, n1099, n41002, n1026, n41001, \PID_CONTROLLER.integral_23__N_3720 , 
        n822, n1029, n764, n40802, n40532, n895, n271, n344, 
        n1102, n125, n56, n198, n417, n6;
    wire [3:0]n19933;
    wire [4:0]n19873;
    
    wire n968, n4;
    wire [2:0]n19973;
    wire [1:0]n19997;
    
    wire n490, n12_adj_4522, n8_adj_4523, n11_adj_4524, n6_adj_4525, 
        n40133, n18, n13_adj_4526, n4_adj_4527, n47634, n271_adj_4528, 
        n122, n53, n344_adj_4529, n1041, n195, n417_adj_4530, n6_adj_4531;
    wire [3:0]n19957;
    wire [4:0]n19908;
    
    wire n204, n338, n40709;
    wire [1:0]n20005;
    
    wire n131, n62, n4_adj_4534;
    wire [2:0]n19988;
    
    wire n691, n40801, n490_adj_4535, n12_adj_4536, n8_adj_4537, n11_adj_4538, 
        n6_adj_4539, n40174, n18_adj_4540, n13_adj_4541, n4_adj_4542, 
        n47516, n268, n107, n38, n77, n8_adj_4544, n1114, n341, 
        n180, n150, n223, n296, n53501, n414, n253;
    wire [23:0]n1_adj_4942;
    
    wire n560, n953, n41000, n618, n40800, n880, n40999, n40615, 
        n807, n40998, n265, n40708, n40531, n734, n40997, n545, 
        n40799, n192, n40707;
    wire [23:0]duty_23__N_3648;
    
    wire n40614, n40613, n40530, n661, n40996, n588, n40995, n50, 
        n119, n11_adj_4547, n51738, n53471, n51726, n472, n40798, 
        n515, n40994, n399, n40797, n40612, n442, n40993, n454;
    wire [5:0]n19789;
    
    wire n560_adj_4548, n40706, n369, n40992, n326, n40796, n487, 
        n40705, n40529, n40795, n527, n600, n101, n32, n40611, 
        n40704, n40528, n40610;
    wire [16:0]n16137;
    wire [15:0]n16749;
    
    wire n40887, n40527, n40991, n43, n19_adj_4550, n51673, n40990, 
        n40886, n53465, n40989, n174, n673, n247, n746, n40609, 
        n819, n40794, n40703, n40885;
    wire [19:0]n13852;
    
    wire n40988, n40526, n12_adj_4552, n51401, n320, n892, n53489, 
        n10_adj_4555, n40702, n40987, n17_adj_4556, n8_adj_4557;
    wire [5:0]n19837;
    
    wire n40793, n40792, n40986, n30, n40701, n40985, n965, n40884, 
        n40791, n53484, n51736, n52081, n393, n40984, n40525, 
        n40790, n40608, n40700, n40883, n40699, n40983, n466, 
        n1038, n40789, n40982, n40698, n40607, n40697, n40882, 
        n40524, n40606, n40981, n40881, n40605, n40523, n40522, 
        n40604, n198_adj_4559, n40696, n53479, n56_adj_4560, n125_adj_4561, 
        n749, n40880, n40521, n676, n40879, n956, n40980, n603, 
        n40878, n107_adj_4562, n883, n40979, n530, n40877, n38_adj_4563, 
        n40520, n810, n40978, n51410, n1111, n180_adj_4565, n253_adj_4567, 
        n737, n40977, n16_adj_4568, n45, n24_adj_4569, n40519, n53469, 
        n457, n40876, n326_adj_4570, n664, n40976, n539, n399_adj_4571, 
        n612, n685, n51951, n472_adj_4573;
    wire [23:0]n1_adj_4943;
    
    wire n545_adj_4576, n618_adj_4577, n691_adj_4578, n758, n591, 
        n40975, n764_adj_4580, n837_adj_4581, n910_adj_4582, n104_adj_4583, 
        n35_adj_4584, n831, n177_adj_4585, n250, n323, n396, n86, 
        n17_adj_4586, n384, n40875, n159, n469, n53495, n542, 
        n518, n40974, n615, n688, n445, n40973, n311, n40874, 
        n372, n40972, n238, n40873, n904, n761, n834, n232, 
        n977;
    wire [0:0]n10324;
    wire [21:0]n10831;
    
    wire n41572, n907, n980, n1050;
    wire [47:0]n106;
    
    wire n41571, n101_adj_4589, n32_adj_4590, n41570, n299, n40971;
    wire [23:0]duty_23__N_3772;
    wire [0:0]n9793;
    
    wire n40518, n41569, n41568, n41567, n41566, n41565, n1096, 
        n41564, n1023, n41563, n174_adj_4591, n950, n41562;
    wire [47:0]n155;
    
    wire n40517, n247_adj_4592, n305, n877, n41561, n804, n41560, 
        n165, n40872, n731, n41559, n320_adj_4593, n393_adj_4594, 
        n658, n41558, n585, n41557, n512, n41556, n439, n41555, 
        n366, n41554, n293, n41553, n220, n41552, n147_adj_4597, 
        n41551, n5_adj_4598, n74, n23_adj_4599, n92, n226, n40970, 
        n40516, n98, n52185, n29, n53460, n52278, n53457, n16_adj_4600, 
        n51390, n24_adj_4601, n6_adj_4602, n52131, n52132, n51732, 
        n51392, n8_adj_4603, n53455, n52117, n52112;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3723 ;
    
    wire n3_adj_4604, n4_adj_4605, n27, n52159, n29_adj_4606, n52160, 
        n33, n12_adj_4607, n15_adj_4608, n51684, n13_adj_4609, n10_adj_4610, 
        n35_adj_4611, n30_adj_4612, n31, n51690, n51686, n52239, 
        n40515, n466_adj_4613, n539_adj_4614;
    wire [14:0]n17293;
    
    wire n40871, n612_adj_4615, n685_adj_4616, n758_adj_4617, n153_adj_4618, 
        n40969, n40514, n831_adj_4619, n11_adj_4620, n80, n1117, 
        n40870;
    wire [9:0]n19133;
    
    wire n840, n40779;
    wire [20:0]n12475;
    
    wire n41523, n41522, n41521, n767, n40778, n41520, n41519, 
        n41518, n41517, n1099_adj_4621, n41516, n904_adj_4622, n1026_adj_4623, 
        n41515, n953_adj_4624, n41514, n880_adj_4625, n41513, n807_adj_4626, 
        n41512, n694, n40777, n734_adj_4627, n41511, n1044, n40869, 
        n661_adj_4628, n41510, n621, n40776;
    wire [18:0]n14693;
    
    wire n40968, n51775, n977_adj_4629, n1050_adj_4630, n588_adj_4631, 
        n41509, n98_adj_4632, n548, n40775, n29_adj_4633, n40967, 
        n171, n171_adj_4634, n244, n317, n515_adj_4635, n41508, 
        n40966, n390, n442_adj_4636, n41507, n369_adj_4637, n41506, 
        n971, n40868, n40965, n475, n40774, n898, n40867, n402, 
        n40773, n825, n40866, n40964, n329, n40772, n256, n40771, 
        n1105, n40963, n752, n40865, n1032, n40962, n296_adj_4638, 
        n41505, n223_adj_4639, n41504, n959, n40961, n679, n40864, 
        n150_adj_4640, n41503, n886, n40960, n8_adj_4641, n77_adj_4642;
    wire [19:0]n14292;
    
    wire n41502, n41501, n606, n40863, n52314, n41500, n183_adj_4643, 
        n40770, n533, n40862, n41, n110, n378, n41499, n41498, 
        n41497, n460, n40861, n813, n40959, n1102_adj_4647, n41496, 
        n1029_adj_4648, n41495, n463, n536, n609, n682, n451, 
        n956_adj_4649, n41494, n755, n883_adj_4651, n41493, n810_adj_4652, 
        n41492, n737_adj_4653, n41491, n664_adj_4654, n41490, n524, 
        n591_adj_4655, n41489, n40513, n387, n40860, n740, n40958, 
        n518_adj_4656, n41488, n667, n40957, n594, n40956, n828, 
        n445_adj_4657, n41487, n372_adj_4658, n41486, n299_adj_4659, 
        n41485, n37, n52315, n39, n52299, n7_adj_4660, n6_adj_4661, 
        n21_adj_4662, n52109, n23_adj_4663, n52110, n25_adj_4664, 
        n51697, n51675, n52119, n51773, n41_adj_4665, n52274, n51677, 
        n52257, n51781, n52259, n4_adj_4666, n52129, n52130, n51403, 
        n52282, n52114, n52320, n52321, n52293, n226_adj_4667, n41484, 
        n521, n40955, n153_adj_4668, n41483, n11_adj_4669, n80_adj_4670;
    wire [18:0]n15092;
    
    wire n41482, n40512, n314, n40859, n41481, n901, n51394, n52207, 
        n41480, n448, n40954, n241, n40858, n40, \PID_CONTROLLER.integral_23__N_3722 , 
        n52209, n41479, n168, n40857, n375, n40953, n41478, n40511, 
        n1105_adj_4671, n41477, n302, n40952, n1032_adj_4672, n41476, 
        n959_adj_4673, n41475, n229, n40951, n886_adj_4674, n41474, 
        n813_adj_4675, n41473, n40510, n156, n40950, n26_adj_4676, 
        n95, n14_adj_4677, n83;
    wire [7:0]n19613;
    wire [6:0]n19740;
    
    wire n630_adj_4678, n40856, n557_adj_4679, n40855, n39_adj_4680, 
        n41_adj_4681, n45_adj_4682, n37_adj_4683, n23_adj_4684, n25_adj_4685, 
        n43_adj_4686;
    wire [9:0]n19253;
    wire [8:0]n19452;
    
    wire n770, n40949, n29_adj_4687, n31_adj_4688, n35_adj_4689, n11_adj_4690, 
        n13_adj_4691, n15_adj_4692, n27_adj_4693, n697, n40948, n740_adj_4695, 
        n41472, n244_adj_4696, n597, n667_adj_4697, n41471, n624, 
        n40947, n33_adj_4699, n9_adj_4700, n974, n594_adj_4701, n41470, 
        n17_adj_4702, n670, n521_adj_4703, n41469, n551, n40946, 
        n1047, n19_adj_4704;
    wire [23:0]n257;
    
    wire n51636, n478, n40945, n448_adj_4705, n41468, n21_adj_4706, 
        n743, n1120, n317_adj_4707, n375_adj_4708, n41467, n51660, 
        n95_adj_4709, n26_adj_4710, n51654, n168_adj_4711, n12_adj_4712, 
        n302_adj_4713, n41466, n10_adj_4714, n30_adj_4715, n229_adj_4716, 
        n41465, n405, n40944, n51671, n51905, n156_adj_4717, n41464, 
        n51901, n52231, n52053, n52272, n16_adj_4718, n14_adj_4719, 
        n83_adj_4720, n6_adj_4721, n52155, n52156, n241_adj_4722, 
        n8_adj_4723, n24_adj_4724, n390_adj_4725, n484_adj_4727, n40854;
    wire [17:0]n15813;
    
    wire n41463, n314_adj_4728, n387_adj_4729, n51640, n460_adj_4731, 
        n6_adj_4732, n533_adj_4733, n51638, n52121, n51783, n4_adj_4734, 
        n332, n40943, n52153, n52154, n51650, n51648, n52241, 
        n51785, n52316, n52317, n463_adj_4735, n52297, n51642, n40509, 
        n52261, n41462, n51791, n52263, n606_adj_4737, n679_adj_4738, 
        duty_23__N_3771, n52069, n752_adj_4739, n52177, n825_adj_4741, 
        n41_adj_4742, n536_adj_4743, n816, n39_adj_4744, n45_adj_4745, 
        n898_adj_4747, n43_adj_4748, n29_adj_4749, n971_adj_4750, n31_adj_4752, 
        n37_adj_4753, n1044_adj_4754, n1117_adj_4755, n92_adj_4756, 
        n23_adj_4757, n23_adj_4758, n25_adj_4759, n41461, n35_adj_4760, 
        n33_adj_4762, n9_adj_4763, n609_adj_4764, n17_adj_4765, n19_adj_4766, 
        n21_adj_4768, n165_adj_4769, n682_adj_4770, n11_adj_4771, n13_adj_4772, 
        n889, n15_adj_4774, n41460, n27_adj_4776, n411_adj_4777, n40853, 
        n51624, n51618, n40508, n1108, n41459, n12_adj_4778, n238_adj_4779, 
        n1035, n41458, n259_adj_4780, n40942, n755_adj_4781, n962, 
        n41457, n338_adj_4782, n40852, n889_adj_4783, n41456, n186_adj_4784, 
        n40941, n40507, n816_adj_4785, n41455, n311_adj_4786, n743_adj_4787, 
        n41454, n10_adj_4788, n30_adj_4789, n670_adj_4790, n41453, 
        n265_adj_4791, n40851, n51873, n597_adj_4792, n41452, n51869, 
        n44, n113;
    wire [17:0]n15453;
    
    wire n40940, n524_adj_4793, n41451, n451_adj_4794, n41450, n40939, 
        n378_adj_4795, n41449, n192_adj_4796, n40850, n40506, n50_adj_4798, 
        n119_adj_4799, n305_adj_4800, n41448, n52225, n232_adj_4801, 
        n41447, n52037, n159_adj_4802, n41446, n40938;
    wire [13:0]n17773;
    
    wire n1120_adj_4803, n40849, n40505, n17_adj_4804, n86_adj_4805, 
        n1047_adj_4806, n40848;
    wire [16:0]n16460;
    
    wire n41445, n41444, n52270, n41443, n1111_adj_4807, n41442, 
        n16_adj_4808, n1038_adj_4809, n41441, n52149, n965_adj_4810, 
        n41440, n892_adj_4811, n41439, n384_adj_4812, n40937, n819_adj_4813, 
        n41438, n746_adj_4814, n41437, n673_adj_4815, n41436, n974_adj_4816, 
        n40847, n962_adj_4817, n828_adj_4818, n600_adj_4819, n41435, 
        n457_adj_4820, n527_adj_4821, n41434, n530_adj_4822, n40504, 
        n1035_adj_4823, n52150, n8_adj_4824, n24_adj_4825, n454_adj_4826, 
        n41433, n51604, n603_adj_4828, n676_adj_4829, n40672, n381, 
        n41432, n749_adj_4831, n822_adj_4832, n895_adj_4833, n968_adj_4834, 
        n51602, n52123, n51793, n4_adj_4835, n1041_adj_4836, n1114_adj_4837, 
        n52147, n52148, n51614, n51612, n52243, n51795, n308, 
        n41431, n235, n41430, n162, n41429, n52318, n52319, n52295, 
        n51606, n52265, n51801, n52267, n256_adj_4839, n40671, n20_adj_4841, 
        n89, n901_adj_4843, n40846;
    wire [23:0]duty_23__N_3747;
    
    wire n1108_adj_4844, n40936, n40670, n40503, n40669;
    wire [15:0]n17037;
    
    wire n41402, n41401, n41400, n41399, n41398, n41397, n41396, 
        n41395, n41394, n41393, n40668, n40935, n41392, n41391, 
        n40845, n40502, n40934, n41390, n41389, n40844, n41388, 
        n40933, n40667, n40843, n41387, n40842;
    wire [14:0]n17548;
    
    wire n41386, n41385, n41384, n40666, n40501, n41383, n41382, 
        n40665, n40932, n40841, n41381, n40500, n40664, n41380, 
        n41379, n41378, n40663, n40840, n40499, n41377, n41376, 
        n40662, n41375, n40498, n41374, n40661, n40839, n40497, 
        n41373, n41372, n40838;
    wire [13:0]n17997;
    
    wire n41371, n40931, n41370, n40930, n41369, n40660, n9_adj_4847, 
        n17_adj_4848, n40929, n40837, n40659, n41368, n41367, n40928, 
        n41366, n40658, n40496, n40927, n41365, n41364, n5_adj_4849, 
        n51388, n250_adj_4850, n40190, n41363, n41362, n40657, n40926, 
        n40656, n40655, n41361, n189_adj_4851, n41360, n41359, n41358, 
        n323_adj_4852, n262_adj_4853, n40836;
    wire [12:0]n18388;
    
    wire n41357, n396_adj_4854, n41356, n41355, n41354, n41353, 
        n41352, n335, n41351, n41350, n41349, n40654, n41348, 
        n469_adj_4855, n542_adj_4856, n408, n41347, n40925, n41346, 
        n116_adj_4857, n41345, n47_adj_4858, n40653, n40835;
    wire [11:0]n18725;
    
    wire n41344, n41343, n40834, n40924, n41342, n41341, n615_adj_4859, 
        n40833, n40652, n41340, n41339, n41338, n41337, n40923, 
        n41336, n41335, n189_adj_4860, n41334, n74_adj_4861, n5_adj_4862, 
        n481, n41333, n262_adj_4863, n40832;
    wire [10:0]n19012;
    
    wire n41332, n335_adj_4864, n41331, n147_adj_4865, n41330, n688_adj_4866, 
        n40831, n40651, n41329, n41328, n41327, n40650, n41326, 
        n40922, n40830, n40649, n40648, n554, n40921, n40829, 
        n41325, n40828, n220_adj_4867, n40920, n41324, n627, n41323, 
        n40647, n293_adj_4869, n41322, n366_adj_4871, n700, n761_adj_4872, 
        n40646, n40919, n110_adj_4873, n41_adj_4874, n408_adj_4875, 
        n183_adj_4876, n256_adj_4878, n329_adj_4879, n402_adj_4880, 
        n113_adj_4881, n44_adj_4882, n475_adj_4883, n834_adj_4884, n481_adj_4885, 
        n548_adj_4886, n621_adj_4887, n694_adj_4888, n186_adj_4889, 
        n439_adj_4890, n40918, n40645, n40827, n512_adj_4891, n767_adj_4892, 
        n840_adj_4893, n554_adj_4894, n907_adj_4895, n585_adj_4896, 
        n40826, n980_adj_4898, n40917, n627_adj_4899, n40644, n40916, 
        n40643, n40825, n40915, n40642, n40914, n40824, n41031, 
        n40913, n40823, n259_adj_4901, n700_adj_4902, n658_adj_4903, 
        n731_adj_4904, n804_adj_4905, n89_adj_4906, n20_adj_4907, n41030, 
        n41029, n40912, n41028, n40911, n40641, n40910, n41027, 
        n40822, n40640, n332_adj_4908, n40639, n405_adj_4910, n122_adj_4911, 
        n53_adj_4912, n195_adj_4913, n162_adj_4914, n877_adj_4915, n41026, 
        n235_adj_4918, n40638, n950_adj_4920, n268_adj_4921, n478_adj_4923, 
        n41025, n487_adj_4924, n40821, n41024, n770_adj_4925, n40730, 
        n697_adj_4926, n40729, n551_adj_4927, n381_adj_4928, n40909, 
        n1023_adj_4929, n341_adj_4930, n1096_adj_4931, n624_adj_4933, 
        n40637, n414_adj_4936, n40820, n308_adj_4937, n40908, n40636, 
        n40728, n40635, n41023, n40819, n41022, n40727, n40726, 
        n40634, n40818, n41021, n40907, n40633, n40632, n41020, 
        n40906, n40817, n40725, n11_adj_4938, n40631, n40724, n41019, 
        n41018, n41017, n40905, n40723, n9_adj_4939, n40630, n40904, 
        n40816, n40629, n41016, n40815, n40903, n41186, n41185, 
        n41015, n41014, n40722, n41184, n41183, n41182, n40902, 
        n40814, n41181, n41180, n41179, n41178, n40628, n41177, 
        n40901, n40813, n40721, n41013, n40627, n40541, n41012, 
        n40720, n40540, n41011, n40539, n40719, n40626, n40625, 
        n40812, n41010, n40538, n40900, n40537, n40899, n40718, 
        n40898, n40624, n41009, n40811, n40623, n41008, n51433, 
        n41007, n40717, n40810, n51428, n40809, n40716, n40622, 
        n40808, n40715, n40807, n51957, n51708, n51734, n4_adj_4940, 
        n40326, n40267, n51704, n40149, n4_adj_4941, n40224;
    
    SB_LUT4 add_6462_3_lut (.I0(GND_net), .I1(n18557[0]), .I2(n177), .I3(n40805), 
            .O(n18193[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n19353[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_3 (.CI(n40805), .I0(n18557[0]), .I1(n177), .CO(n40806));
    SB_CARRY add_6550_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n40714));
    SB_LUT4 add_6567_9_lut (.I0(GND_net), .I1(n19677[6]), .I2(n630), .I3(n40713), 
            .O(n19533[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_19 (.CI(n41005), .I0(n11990[16]), .I1(GND_net), 
            .CO(n41006));
    SB_LUT4 add_6462_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n18193[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_19 (.CI(n40620), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n40621));
    SB_CARRY add_904_19 (.CI(n40535), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n4096[17]), .CO(n40536));
    SB_LUT4 add_6567_8_lut (.I0(GND_net), .I1(n19677[5]), .I2(n557), .I3(n40712), 
            .O(n19533[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n40805));
    SB_CARRY add_6567_8 (.CI(n40712), .I0(n19677[5]), .I1(n557), .CO(n40713));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n40619), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4572_18_lut (.I0(GND_net), .I1(n11990[15]), .I2(GND_net), 
            .I3(n41004), .O(n10300[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_18 (.CI(n40619), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n40620));
    SB_LUT4 add_904_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n4096[16]), .I3(n40534), .O(\PID_CONTROLLER.integral_23__N_3672 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n40618), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_17 (.CI(n40618), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n40619));
    SB_CARRY add_904_18 (.CI(n40534), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n4096[16]), .CO(n40535));
    SB_LUT4 add_6567_7_lut (.I0(GND_net), .I1(n19677[4]), .I2(n484), .I3(n40711), 
            .O(n19533[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6487_13_lut (.I0(GND_net), .I1(n18869[10]), .I2(n910), 
            .I3(n40804), .O(n18557[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n40617), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6487_12_lut (.I0(GND_net), .I1(n18869[9]), .I2(n837), 
            .I3(n40803), .O(n18557[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_7 (.CI(n40711), .I0(n19677[4]), .I1(n484), .CO(n40712));
    SB_LUT4 add_6567_6_lut (.I0(GND_net), .I1(n19677[3]), .I2(n411), .I3(n40710), 
            .O(n19533[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_18 (.CI(n41004), .I0(n11990[15]), .I1(GND_net), 
            .CO(n41005));
    SB_LUT4 add_4572_17_lut (.I0(GND_net), .I1(n11990[14]), .I2(GND_net), 
            .I3(n41003), .O(n10300[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_16 (.CI(n40617), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n40618));
    SB_CARRY add_6567_6 (.CI(n40710), .I0(n19677[3]), .I1(n411), .CO(n40711));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n40616), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n4096[15]), .I3(n40533), .O(\PID_CONTROLLER.integral_23__N_3672 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_17 (.CI(n40533), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n4096[15]), .CO(n40534));
    SB_CARRY add_4572_17 (.CI(n41003), .I0(n11990[14]), .I1(GND_net), 
            .CO(n41004));
    SB_CARRY add_6487_12 (.CI(n40803), .I0(n18869[9]), .I1(n837), .CO(n40804));
    SB_LUT4 add_4572_16_lut (.I0(GND_net), .I1(n11990[13]), .I2(n1099), 
            .I3(n41002), .O(n10300[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_16 (.CI(n41002), .I0(n11990[13]), .I1(n1099), .CO(n41003));
    SB_LUT4 add_4572_15_lut (.I0(GND_net), .I1(n11990[12]), .I2(n1026), 
            .I3(n41001), .O(n10300[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_15 (.CI(n41001), .I0(n11990[12]), .I1(n1026), .CO(n41002));
    SB_LUT4 i22023_2_lut (.I0(n1[4]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22023_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22022_2_lut (.I0(n1[5]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22022_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6487_11_lut (.I0(GND_net), .I1(n18869[8]), .I2(n764), 
            .I3(n40802), .O(n18557[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22021_2_lut (.I0(n1[6]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22021_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_904_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n4096[14]), .I3(n40532), .O(\PID_CONTROLLER.integral_23__N_3672 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6), .I1(\Ki[4] ), .I2(n19933[2]), .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .O(n19873[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1510 (.I0(n4), .I1(\Ki[3] ), .I2(n19973[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), .O(n19933[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1510.LUT_INIT = 16'h965a;
    SB_LUT4 i26645_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n19997[0]));   // verilog/motorControl.v(34[25:36])
    defparam i26645_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1511 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [20]), .O(n12_adj_4522));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1511.LUT_INIT = 16'h9c50;
    SB_LUT4 i26758_4_lut (.I0(n19933[2]), .I1(\Ki[4] ), .I2(n6), .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .O(n8_adj_4523));   // verilog/motorControl.v(34[25:36])
    defparam i26758_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n11_adj_4524));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i26719_4_lut (.I0(n19973[1]), .I1(\Ki[3] ), .I2(n4), .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .O(n6_adj_4525));   // verilog/motorControl.v(34[25:36])
    defparam i26719_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i26647_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n40133));   // verilog/motorControl.v(34[25:36])
    defparam i26647_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4525), .I1(n11_adj_4524), .I2(n8_adj_4523), 
            .I3(n12_adj_4522), .O(n18));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [22]), .O(n13_adj_4526));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4526), .I1(n18), .I2(n40133), .I3(n4_adj_4527), 
            .O(n47634));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4528));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22020_2_lut (.I0(n1[7]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22020_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4529));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4530));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1512 (.I0(n6_adj_4531), .I1(\Kp[4] ), .I2(n19957[2]), 
            .I3(n1[18]), .O(n19908[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1512.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6567_5_lut (.I0(GND_net), .I1(n19677[2]), .I2(n338), .I3(n40709), 
            .O(n19533[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26683_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n20005[0]));   // verilog/motorControl.v(34[16:22])
    defparam i26683_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1513 (.I0(n4_adj_4534), .I1(\Kp[3] ), .I2(n19988[1]), 
            .I3(n1[19]), .O(n19957[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1513.LUT_INIT = 16'h965a;
    SB_CARRY add_6487_11 (.CI(n40802), .I0(n18869[8]), .I1(n764), .CO(n40803));
    SB_LUT4 add_6487_10_lut (.I0(GND_net), .I1(n18869[7]), .I2(n691), 
            .I3(n40801), .O(n18557[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4535));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1514 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n1[23]), 
            .I3(n1[20]), .O(n12_adj_4536));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1514.LUT_INIT = 16'h9c50;
    SB_LUT4 i26851_4_lut (.I0(n19957[2]), .I1(\Kp[4] ), .I2(n6_adj_4531), 
            .I3(n1[18]), .O(n8_adj_4537));   // verilog/motorControl.v(34[16:22])
    defparam i26851_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1515 (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n1[19]), 
            .I3(n1[21]), .O(n11_adj_4538));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut_adj_1515.LUT_INIT = 16'h6ca0;
    SB_LUT4 i26812_4_lut (.I0(n19988[1]), .I1(\Kp[3] ), .I2(n4_adj_4534), 
            .I3(n1[19]), .O(n6_adj_4539));   // verilog/motorControl.v(34[16:22])
    defparam i26812_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i26685_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n40174));   // verilog/motorControl.v(34[16:22])
    defparam i26685_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1516 (.I0(n6_adj_4539), .I1(n11_adj_4538), .I2(n8_adj_4537), 
            .I3(n12_adj_4536), .O(n18_adj_4540));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut_adj_1516.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1517 (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n1[18]), 
            .I3(n1[22]), .O(n13_adj_4541));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut_adj_1517.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1518 (.I0(n13_adj_4541), .I1(n18_adj_4540), .I2(n40174), 
            .I3(n4_adj_4542), .O(n47516));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_CARRY sub_3_add_2_15 (.CI(n40616), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n40617));
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22019_2_lut (.I0(n1[8]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22019_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4544));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22018_2_lut (.I0(n1[9]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22018_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22017_2_lut (.I0(n1[10]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22017_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_175_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n53501));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_175_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22016_2_lut (.I0(n1[11]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22016_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6487_10 (.CI(n40801), .I0(n18869[7]), .I1(n691), .CO(n40802));
    SB_CARRY add_6567_5 (.CI(n40709), .I0(n19677[2]), .I1(n338), .CO(n40710));
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4572_14_lut (.I0(GND_net), .I1(n11990[11]), .I2(n953), 
            .I3(n41000), .O(n10300[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6487_9_lut (.I0(GND_net), .I1(n18869[6]), .I2(n618), .I3(n40800), 
            .O(n18557[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_14 (.CI(n41000), .I0(n11990[11]), .I1(n953), .CO(n41001));
    SB_CARRY add_904_16 (.CI(n40532), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n4096[14]), .CO(n40533));
    SB_LUT4 add_4572_13_lut (.I0(GND_net), .I1(n11990[10]), .I2(n880), 
            .I3(n40999), .O(n10300[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n40615), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_13 (.CI(n40999), .I0(n11990[10]), .I1(n880), .CO(n41000));
    SB_LUT4 add_4572_12_lut (.I0(GND_net), .I1(n11990[9]), .I2(n807), 
            .I3(n40998), .O(n10300[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_9 (.CI(n40800), .I0(n18869[6]), .I1(n618), .CO(n40801));
    SB_CARRY add_4572_12 (.CI(n40998), .I0(n11990[9]), .I1(n807), .CO(n40999));
    SB_LUT4 add_6567_4_lut (.I0(GND_net), .I1(n19677[1]), .I2(n265), .I3(n40708), 
            .O(n19533[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n4096[13]), .I3(n40531), .O(\PID_CONTROLLER.integral_23__N_3672 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4572_11_lut (.I0(GND_net), .I1(n11990[8]), .I2(n734), 
            .I3(n40997), .O(n10300[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_14 (.CI(n40615), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n40616));
    SB_LUT4 add_6487_8_lut (.I0(GND_net), .I1(n18869[5]), .I2(n545), .I3(n40799), 
            .O(n18557[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_4 (.CI(n40708), .I0(n19677[1]), .I1(n265), .CO(n40709));
    SB_LUT4 add_6567_3_lut (.I0(GND_net), .I1(n19677[0]), .I2(n192), .I3(n40707), 
            .O(n19533[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_8 (.CI(n40799), .I0(n18869[5]), .I1(n545), .CO(n40800));
    SB_CARRY add_6567_3 (.CI(n40707), .I0(n19677[0]), .I1(n192), .CO(n40708));
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3648[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_4572_11 (.CI(n40997), .I0(n11990[8]), .I1(n734), .CO(n40998));
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n40614), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY sub_3_add_2_13 (.CI(n40614), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n40615));
    SB_CARRY add_904_15 (.CI(n40531), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n4096[13]), .CO(n40532));
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n40613), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n4096[12]), .I3(n40530), .O(\PID_CONTROLLER.integral_23__N_3672 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4572_10_lut (.I0(GND_net), .I1(n11990[7]), .I2(n661), 
            .I3(n40996), .O(n10300[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_10 (.CI(n40996), .I0(n11990[7]), .I1(n661), .CO(n40997));
    SB_LUT4 add_4572_9_lut (.I0(GND_net), .I1(n11990[6]), .I2(n588), .I3(n40995), 
            .O(n10300[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6567_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n19533[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_12 (.CI(n40613), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n40614));
    SB_LUT4 i36256_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n53501), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4547), .O(n51738));
    defparam i36256_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_145_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n53471));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_145_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36244_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n53471), 
            .I2(IntegralLimit[14]), .I3(n51738), .O(n51726));
    defparam i36244_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY add_4572_9 (.CI(n40995), .I0(n11990[6]), .I1(n588), .CO(n40996));
    SB_LUT4 add_6487_7_lut (.I0(GND_net), .I1(n18869[4]), .I2(n472), .I3(n40798), 
            .O(n18557[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4572_8_lut (.I0(GND_net), .I1(n11990[5]), .I2(n515), .I3(n40994), 
            .O(n10300[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n40707));
    SB_CARRY add_4572_8 (.CI(n40994), .I0(n11990[5]), .I1(n515), .CO(n40995));
    SB_CARRY add_6487_7 (.CI(n40798), .I0(n18869[4]), .I1(n472), .CO(n40799));
    SB_LUT4 add_6487_6_lut (.I0(GND_net), .I1(n18869[3]), .I2(n399), .I3(n40797), 
            .O(n18557[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n40612), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_14 (.CI(n40530), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n4096[12]), .CO(n40531));
    SB_LUT4 add_4572_7_lut (.I0(GND_net), .I1(n11990[4]), .I2(n442), .I3(n40993), 
            .O(n10300[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_7 (.CI(n40993), .I0(n11990[4]), .I1(n442), .CO(n40994));
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6582_8_lut (.I0(GND_net), .I1(n19789[5]), .I2(n560_adj_4548), 
            .I3(n40706), .O(n19677[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4572_6_lut (.I0(GND_net), .I1(n11990[3]), .I2(n369), .I3(n40992), 
            .O(n10300[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_6 (.CI(n40797), .I0(n18869[3]), .I1(n399), .CO(n40798));
    SB_CARRY sub_3_add_2_11 (.CI(n40612), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n40613));
    SB_LUT4 add_6487_5_lut (.I0(GND_net), .I1(n18869[2]), .I2(n326), .I3(n40796), 
            .O(n18557[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_5 (.CI(n40796), .I0(n18869[2]), .I1(n326), .CO(n40797));
    SB_LUT4 add_6582_7_lut (.I0(GND_net), .I1(n19789[4]), .I2(n487), .I3(n40705), 
            .O(n19677[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_904_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n4096[11]), .I3(n40529), .O(\PID_CONTROLLER.integral_23__N_3672 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_6 (.CI(n40992), .I0(n11990[3]), .I1(n369), .CO(n40993));
    SB_CARRY add_6582_7 (.CI(n40705), .I0(n19789[4]), .I1(n487), .CO(n40706));
    SB_LUT4 add_6487_4_lut (.I0(GND_net), .I1(n18869[1]), .I2(n253), .I3(n40795), 
            .O(n18557[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_4 (.CI(n40795), .I0(n18869[1]), .I1(n253), .CO(n40796));
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n40611), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_13 (.CI(n40529), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n4096[11]), .CO(n40530));
    SB_CARRY sub_3_add_2_10 (.CI(n40611), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n40612));
    SB_LUT4 add_6582_6_lut (.I0(GND_net), .I1(n19789[3]), .I2(n414), .I3(n40704), 
            .O(n19677[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n4096[10]), .I3(n40528), .O(\PID_CONTROLLER.integral_23__N_3672 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n40610), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_18_lut (.I0(GND_net), .I1(n16749[15]), .I2(GND_net), 
            .I3(n40887), .O(n16137[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_12 (.CI(n40528), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n4096[10]), .CO(n40529));
    SB_LUT4 add_904_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n4096[9]), .I3(n40527), .O(\PID_CONTROLLER.integral_23__N_3672 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_9 (.CI(n40610), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n40611));
    SB_LUT4 add_4572_5_lut (.I0(GND_net), .I1(n11990[2]), .I2(n296), .I3(n40991), 
            .O(n10300[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_5 (.CI(n40991), .I0(n11990[2]), .I1(n296), .CO(n40992));
    SB_LUT4 i36191_2_lut (.I0(n43), .I1(n19_adj_4550), .I2(GND_net), .I3(GND_net), 
            .O(n51673));
    defparam i36191_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_4572_4_lut (.I0(GND_net), .I1(n11990[1]), .I2(n223), .I3(n40990), 
            .O(n10300[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_17_lut (.I0(GND_net), .I1(n16749[14]), .I2(GND_net), 
            .I3(n40886), .O(n16137[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_139_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n53465));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_139_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6582_6 (.CI(n40704), .I0(n19789[3]), .I1(n414), .CO(n40705));
    SB_CARRY add_4572_4 (.CI(n40990), .I0(n11990[1]), .I1(n223), .CO(n40991));
    SB_LUT4 add_4572_3_lut (.I0(GND_net), .I1(n11990[0]), .I2(n150), .I3(n40989), 
            .O(n10300[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_11 (.CI(n40527), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n4096[9]), .CO(n40528));
    SB_CARRY add_6342_17 (.CI(n40886), .I0(n16749[14]), .I1(GND_net), 
            .CO(n40887));
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n40609), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6487_3_lut (.I0(GND_net), .I1(n18869[0]), .I2(n180), .I3(n40794), 
            .O(n18557[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_3 (.CI(n40989), .I0(n11990[0]), .I1(n150), .CO(n40990));
    SB_LUT4 add_6582_5_lut (.I0(GND_net), .I1(n19789[2]), .I2(n341), .I3(n40703), 
            .O(n19677[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_16_lut (.I0(GND_net), .I1(n16749[13]), .I2(n1114), 
            .I3(n40885), .O(n16137[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4572_2_lut (.I0(GND_net), .I1(n8_adj_4544), .I2(n77), 
            .I3(GND_net), .O(n10300[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_3 (.CI(n40794), .I0(n18869[0]), .I1(n180), .CO(n40795));
    SB_CARRY add_6582_5 (.CI(n40703), .I0(n19789[2]), .I1(n341), .CO(n40704));
    SB_LUT4 add_6487_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n18557[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_2 (.CI(GND_net), .I0(n8_adj_4544), .I1(n77), .CO(n40989));
    SB_CARRY add_6487_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n40794));
    SB_LUT4 add_5251_22_lut (.I0(GND_net), .I1(n13852[19]), .I2(GND_net), 
            .I3(n40988), .O(n11990[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n4096[8]), .I3(n40526), .O(\PID_CONTROLLER.integral_23__N_3672 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_8 (.CI(n40609), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n40610));
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4552));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35919_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n51401));
    defparam i35919_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_163_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n53489));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_163_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4555));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6582_4_lut (.I0(GND_net), .I1(n19789[1]), .I2(n268), .I3(n40702), 
            .O(n19677[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6582_4 (.CI(n40702), .I0(n19789[1]), .I1(n268), .CO(n40703));
    SB_LUT4 add_5251_21_lut (.I0(GND_net), .I1(n13852[18]), .I2(GND_net), 
            .I3(n40987), .O(n11990[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_16 (.CI(n40885), .I0(n16749[13]), .I1(n1114), .CO(n40886));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4556), .I3(GND_net), 
            .O(n8_adj_4557));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_6601_7_lut (.I0(GND_net), .I1(n47516), .I2(n490_adj_4535), 
            .I3(n40793), .O(n19837[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_21 (.CI(n40987), .I0(n13852[18]), .I1(GND_net), 
            .CO(n40988));
    SB_CARRY add_904_10 (.CI(n40526), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n4096[8]), .CO(n40527));
    SB_LUT4 add_6601_6_lut (.I0(GND_net), .I1(n19908[3]), .I2(n417_adj_4530), 
            .I3(n40792), .O(n19837[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5251_20_lut (.I0(GND_net), .I1(n13852[17]), .I2(GND_net), 
            .I3(n40986), .O(n11990[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_20 (.CI(n40986), .I0(n13852[17]), .I1(GND_net), 
            .CO(n40987));
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4552), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6582_3_lut (.I0(GND_net), .I1(n19789[0]), .I2(n195), .I3(n40701), 
            .O(n19677[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6582_3 (.CI(n40701), .I0(n19789[0]), .I1(n195), .CO(n40702));
    SB_LUT4 add_5251_19_lut (.I0(GND_net), .I1(n13852[16]), .I2(GND_net), 
            .I3(n40985), .O(n11990[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5251_19 (.CI(n40985), .I0(n13852[16]), .I1(GND_net), 
            .CO(n40986));
    SB_CARRY add_6601_6 (.CI(n40792), .I0(n19908[3]), .I1(n417_adj_4530), 
            .CO(n40793));
    SB_LUT4 add_6342_15_lut (.I0(GND_net), .I1(n16749[12]), .I2(n1041), 
            .I3(n40884), .O(n16137[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6601_5_lut (.I0(GND_net), .I1(n19908[2]), .I2(n344_adj_4529), 
            .I3(n40791), .O(n19837[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36598_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n53484), 
            .I2(IntegralLimit[11]), .I3(n51736), .O(n52081));
    defparam i36598_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5251_18_lut (.I0(GND_net), .I1(n13852[15]), .I2(GND_net), 
            .I3(n40984), .O(n11990[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n4096[7]), .I3(n40525), .O(\PID_CONTROLLER.integral_23__N_3672 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_18 (.CI(n40984), .I0(n13852[15]), .I1(GND_net), 
            .CO(n40985));
    SB_LUT4 add_6582_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n19677[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_5 (.CI(n40791), .I0(n19908[2]), .I1(n344_adj_4529), 
            .CO(n40792));
    SB_LUT4 add_6601_4_lut (.I0(GND_net), .I1(n19908[1]), .I2(n271_adj_4528), 
            .I3(n40790), .O(n19837[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6582_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n40701));
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n40608), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_15 (.CI(n40884), .I0(n16749[12]), .I1(n1041), .CO(n40885));
    SB_LUT4 add_6595_7_lut (.I0(GND_net), .I1(n47634), .I2(n490), .I3(n40700), 
            .O(n19789[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_14_lut (.I0(GND_net), .I1(n16749[11]), .I2(n968), 
            .I3(n40883), .O(n16137[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6595_6_lut (.I0(GND_net), .I1(n19873[3]), .I2(n417), .I3(n40699), 
            .O(n19789[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6595_6 (.CI(n40699), .I0(n19873[3]), .I1(n417), .CO(n40700));
    SB_CARRY add_6601_4 (.CI(n40790), .I0(n19908[1]), .I1(n271_adj_4528), 
            .CO(n40791));
    SB_CARRY sub_3_add_2_7 (.CI(n40608), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n40609));
    SB_CARRY add_6342_14 (.CI(n40883), .I0(n16749[11]), .I1(n968), .CO(n40884));
    SB_LUT4 add_5251_17_lut (.I0(GND_net), .I1(n13852[14]), .I2(GND_net), 
            .I3(n40983), .O(n11990[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5251_17 (.CI(n40983), .I0(n13852[14]), .I1(GND_net), 
            .CO(n40984));
    SB_CARRY add_904_9 (.CI(n40525), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n4096[7]), .CO(n40526));
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6601_3_lut (.I0(GND_net), .I1(n19908[0]), .I2(n198), .I3(n40789), 
            .O(n19837[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_3 (.CI(n40789), .I0(n19908[0]), .I1(n198), .CO(n40790));
    SB_LUT4 add_6601_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n19837[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5251_16_lut (.I0(GND_net), .I1(n13852[13]), .I2(n1102), 
            .I3(n40982), .O(n11990[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6595_5_lut (.I0(GND_net), .I1(n19873[2]), .I2(n344), .I3(n40698), 
            .O(n19789[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n40607), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_16 (.CI(n40982), .I0(n13852[13]), .I1(n1102), .CO(n40983));
    SB_CARRY add_6595_5 (.CI(n40698), .I0(n19873[2]), .I1(n344), .CO(n40699));
    SB_CARRY sub_3_add_2_6 (.CI(n40607), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n40608));
    SB_LUT4 add_6595_4_lut (.I0(GND_net), .I1(n19873[1]), .I2(n271), .I3(n40697), 
            .O(n19789[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_13_lut (.I0(GND_net), .I1(n16749[10]), .I2(n895), 
            .I3(n40882), .O(n16137[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n40789));
    SB_LUT4 add_904_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n4096[6]), .I3(n40524), .O(\PID_CONTROLLER.integral_23__N_3672 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6595_4 (.CI(n40697), .I0(n19873[1]), .I1(n271), .CO(n40698));
    SB_CARRY add_6342_13 (.CI(n40882), .I0(n16749[10]), .I1(n895), .CO(n40883));
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n40606), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5251_15_lut (.I0(GND_net), .I1(n13852[12]), .I2(n1029), 
            .I3(n40981), .O(n11990[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_5 (.CI(n40606), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n40607));
    SB_CARRY add_904_8 (.CI(n40524), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n4096[6]), .CO(n40525));
    SB_LUT4 add_6342_12_lut (.I0(GND_net), .I1(n16749[9]), .I2(n822), 
            .I3(n40881), .O(n16137[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n40605), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n4096[5]), .I3(n40523), .O(\PID_CONTROLLER.integral_23__N_3672 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_7 (.CI(n40523), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n4096[5]), .CO(n40524));
    SB_LUT4 add_904_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n4096[4]), .I3(n40522), .O(\PID_CONTROLLER.integral_23__N_3672 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_4 (.CI(n40605), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n40606));
    SB_CARRY add_904_6 (.CI(n40522), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n4096[4]), .CO(n40523));
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n40604), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6595_3_lut (.I0(GND_net), .I1(n19873[0]), .I2(n198_adj_4559), 
            .I3(n40696), .O(n19789[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_153_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n53479));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_153_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_3_add_2_3 (.CI(n40604), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n40605));
    SB_CARRY add_6595_3 (.CI(n40696), .I0(n19873[0]), .I1(n198_adj_4559), 
            .CO(n40697));
    SB_CARRY add_6342_12 (.CI(n40881), .I0(n16749[9]), .I1(n822), .CO(n40882));
    SB_LUT4 add_6595_2_lut (.I0(GND_net), .I1(n56_adj_4560), .I2(n125_adj_4561), 
            .I3(GND_net), .O(n19789[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_11_lut (.I0(GND_net), .I1(n16749[8]), .I2(n749), 
            .I3(n40880), .O(n16137[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6595_2 (.CI(GND_net), .I0(n56_adj_4560), .I1(n125_adj_4561), 
            .CO(n40696));
    SB_LUT4 add_904_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n4096[3]), .I3(n40521), .O(\PID_CONTROLLER.integral_23__N_3672 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_15 (.CI(n40981), .I0(n13852[12]), .I1(n1029), .CO(n40982));
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n40604));
    SB_CARRY add_6342_11 (.CI(n40880), .I0(n16749[8]), .I1(n749), .CO(n40881));
    SB_LUT4 add_6342_10_lut (.I0(GND_net), .I1(n16749[7]), .I2(n676), 
            .I3(n40879), .O(n16137[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5251_14_lut (.I0(GND_net), .I1(n13852[11]), .I2(n956), 
            .I3(n40980), .O(n11990[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_10 (.CI(n40879), .I0(n16749[7]), .I1(n676), .CO(n40880));
    SB_LUT4 add_6342_9_lut (.I0(GND_net), .I1(n16749[6]), .I2(n603), .I3(n40878), 
            .O(n16137[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_9 (.CI(n40878), .I0(n16749[6]), .I1(n603), .CO(n40879));
    SB_CARRY add_5251_14 (.CI(n40980), .I0(n13852[11]), .I1(n956), .CO(n40981));
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4562));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5251_13_lut (.I0(GND_net), .I1(n13852[10]), .I2(n883), 
            .I3(n40979), .O(n11990[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_8_lut (.I0(GND_net), .I1(n16749[5]), .I2(n530), .I3(n40877), 
            .O(n16137[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4563));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5251_13 (.CI(n40979), .I0(n13852[10]), .I1(n883), .CO(n40980));
    SB_CARRY add_904_5 (.CI(n40521), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n4096[3]), .CO(n40522));
    SB_LUT4 add_904_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n4096[2]), .I3(n40520), .O(\PID_CONTROLLER.integral_23__N_3672 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5251_12_lut (.I0(GND_net), .I1(n13852[9]), .I2(n810), 
            .I3(n40978), .O(n11990[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35928_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n53479), 
            .I2(IntegralLimit[13]), .I3(n52081), .O(n51410));
    defparam i35928_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_5251_12 (.CI(n40978), .I0(n13852[9]), .I1(n810), .CO(n40979));
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4565));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4567));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6342_8 (.CI(n40877), .I0(n16749[5]), .I1(n530), .CO(n40878));
    SB_CARRY add_904_4 (.CI(n40520), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n4096[2]), .CO(n40521));
    SB_LUT4 add_5251_11_lut (.I0(GND_net), .I1(n13852[8]), .I2(n737), 
            .I3(n40977), .O(n11990[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4568), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_4569));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_904_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n4096[1]), .I3(n40519), .O(\PID_CONTROLLER.integral_23__N_3672 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_3 (.CI(n40519), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n4096[1]), .CO(n40520));
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_143_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n53469));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_143_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5251_11 (.CI(n40977), .I0(n13852[8]), .I1(n737), .CO(n40978));
    SB_LUT4 add_6342_7_lut (.I0(GND_net), .I1(n16749[4]), .I2(n457), .I3(n40876), 
            .O(n16137[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4570));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5251_10_lut (.I0(GND_net), .I1(n13852[7]), .I2(n664), 
            .I3(n40976), .O(n11990[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4571));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6342_7 (.CI(n40876), .I0(n16749[4]), .I1(n457), .CO(n40877));
    SB_LUT4 i36468_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n53469), 
            .I2(IntegralLimit[15]), .I3(n51410), .O(n51951));
    defparam i36468_4_lut.LUT_INIT = 16'hffde;
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_5251_10 (.CI(n40976), .I0(n13852[7]), .I1(n664), .CO(n40977));
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3648[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3648[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3648[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3648[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3648[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3648[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3648[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3648[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3648[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3648[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3648[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3648[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3648[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3648[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3648[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3648[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3648[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3648[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3648[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3648[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3648[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3648[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3648[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4573));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4576));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4577));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4578));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5251_9_lut (.I0(GND_net), .I1(n13852[6]), .I2(n591), .I3(n40975), 
            .O(n11990[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n4096[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3672 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4580));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4581));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4582));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4583));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4584));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4585));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5251_9 (.CI(n40975), .I0(n13852[6]), .I1(n591), .CO(n40976));
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4586));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6342_6_lut (.I0(GND_net), .I1(n16749[3]), .I2(n384), .I3(n40875), 
            .O(n16137[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_904_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n4096[0]), .CO(n40519));
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_169_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n53495));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_169_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5251_8_lut (.I0(GND_net), .I1(n13852[5]), .I2(n518), .I3(n40974), 
            .O(n11990[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6342_6 (.CI(n40875), .I0(n16749[3]), .I1(n384), .CO(n40876));
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5251_8 (.CI(n40974), .I0(n13852[5]), .I1(n518), .CO(n40975));
    SB_LUT4 add_5251_7_lut (.I0(GND_net), .I1(n13852[4]), .I2(n445), .I3(n40973), 
            .O(n11990[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_5_lut (.I0(GND_net), .I1(n16749[2]), .I2(n311), .I3(n40874), 
            .O(n16137[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_7 (.CI(n40973), .I0(n13852[4]), .I1(n445), .CO(n40974));
    SB_LUT4 add_5251_6_lut (.I0(GND_net), .I1(n13852[3]), .I2(n372), .I3(n40972), 
            .O(n11990[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_5 (.CI(n40874), .I0(n16749[2]), .I1(n311), .CO(n40875));
    SB_LUT4 add_6342_4_lut (.I0(GND_net), .I1(n16749[1]), .I2(n238), .I3(n40873), 
            .O(n16137[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_6 (.CI(n40972), .I0(n13852[3]), .I1(n372), .CO(n40973));
    SB_CARRY add_6342_4 (.CI(n40873), .I0(n16749[1]), .I1(n238), .CO(n40874));
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n1[23]), .I1(n10831[21]), .I2(GND_net), 
            .I3(n41572), .O(n10324[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n10831[20]), .I2(GND_net), 
            .I3(n41571), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4589));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4590));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_23 (.CI(n41571), .I0(n10831[20]), .I1(GND_net), 
            .CO(n41572));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n10831[19]), .I2(GND_net), 
            .I3(n41570), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5251_5_lut (.I0(GND_net), .I1(n13852[2]), .I2(n299), .I3(n40971), 
            .O(n11990[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n10324[0]), .I2(n9793[0]), 
            .I3(n40518), .O(duty_23__N_3772[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n41570), .I0(n10831[19]), .I1(GND_net), 
            .CO(n41571));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n10831[18]), .I2(GND_net), 
            .I3(n41569), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n41569), .I0(n10831[18]), .I1(GND_net), 
            .CO(n41570));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n10831[17]), .I2(GND_net), 
            .I3(n41568), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_20 (.CI(n41568), .I0(n10831[17]), .I1(GND_net), 
            .CO(n41569));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n10831[16]), .I2(GND_net), 
            .I3(n41567), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n41567), .I0(n10831[16]), .I1(GND_net), 
            .CO(n41568));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n10831[15]), .I2(GND_net), 
            .I3(n41566), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n41566), .I0(n10831[15]), .I1(GND_net), 
            .CO(n41567));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n10831[14]), .I2(GND_net), 
            .I3(n41565), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n41565), .I0(n10831[14]), .I1(GND_net), 
            .CO(n41566));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n10831[13]), .I2(n1096), 
            .I3(n41564), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n41564), .I0(n10831[13]), .I1(n1096), 
            .CO(n41565));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n10831[12]), .I2(n1023), 
            .I3(n41563), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4591));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_15 (.CI(n41563), .I0(n10831[12]), .I1(n1023), 
            .CO(n41564));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n10831[11]), .I2(n950), 
            .I3(n41562), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n40517), .O(duty_23__N_3772[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n41562), .I0(n10831[11]), .I1(n950), 
            .CO(n41563));
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4592));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n10831[10]), .I2(n877), 
            .I3(n41561), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n41561), .I0(n10831[10]), .I1(n877), 
            .CO(n41562));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n10831[9]), .I2(n804), 
            .I3(n41560), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_3_lut (.I0(GND_net), .I1(n16749[0]), .I2(n165), .I3(n40872), 
            .O(n16137[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n41560), .I0(n10831[9]), .I1(n804), 
            .CO(n41561));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n10831[8]), .I2(n731), 
            .I3(n41559), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n41559), .I0(n10831[8]), .I1(n731), 
            .CO(n41560));
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4593));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4594));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n10831[7]), .I2(n658), 
            .I3(n41558), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n41558), .I0(n10831[7]), .I1(n658), 
            .CO(n41559));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n10831[6]), .I2(n585), 
            .I3(n41557), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n41557), .I0(n10831[6]), .I1(n585), 
            .CO(n41558));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n10831[5]), .I2(n512), 
            .I3(n41556), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_5 (.CI(n40971), .I0(n13852[2]), .I1(n299), .CO(n40972));
    SB_CARRY mult_10_add_1225_8 (.CI(n41556), .I0(n10831[5]), .I1(n512), 
            .CO(n41557));
    SB_CARRY add_6342_3 (.CI(n40872), .I0(n16749[0]), .I1(n165), .CO(n40873));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n10831[4]), .I2(n439), 
            .I3(n41555), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n41555), .I0(n10831[4]), .I1(n439), 
            .CO(n41556));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n10831[3]), .I2(n366), 
            .I3(n41554), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n41554), .I0(n10831[3]), .I1(n366), 
            .CO(n41555));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n10831[2]), .I2(n293), 
            .I3(n41553), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n41553), .I0(n10831[2]), .I1(n293), 
            .CO(n41554));
    SB_CARRY add_12_24 (.CI(n40517), .I0(n106[22]), .I1(n155[22]), .CO(n40518));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n10831[1]), .I2(n220), 
            .I3(n41552), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n41552), .I0(n10831[1]), .I1(n220), 
            .CO(n41553));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n10831[0]), .I2(n147_adj_4597), 
            .I3(n41551), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n41551), .I0(n10831[0]), .I1(n147_adj_4597), 
            .CO(n41552));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4598), .I2(n74), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_2_lut (.I0(GND_net), .I1(n23_adj_4599), .I2(n92), 
            .I3(GND_net), .O(n16137[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4598), .I1(n74), 
            .CO(n41551));
    SB_LUT4 add_5251_4_lut (.I0(GND_net), .I1(n13852[1]), .I2(n226), .I3(n40970), 
            .O(n11990[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n40516), .O(duty_23__N_3772[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36702_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n53495), 
            .I2(IntegralLimit[17]), .I3(n51951), .O(n52185));
    defparam i36702_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_12_23 (.CI(n40516), .I0(n106[21]), .I1(n155[21]), .CO(n40517));
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6342_2 (.CI(GND_net), .I0(n23_adj_4599), .I1(n92), .CO(n40872));
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_134_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n53460));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_134_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36795_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n53460), 
            .I2(IntegralLimit[19]), .I3(n52185), .O(n52278));
    defparam i36795_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_131_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n53457));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_131_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4600));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35908_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n51390));
    defparam i35908_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4600), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4601));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4602));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36648_3_lut (.I0(n6_adj_4602), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n52131));   // verilog/motorControl.v(31[10:34])
    defparam i36648_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36649_3_lut (.I0(n52131), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n52132));   // verilog/motorControl.v(31[10:34])
    defparam i36649_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35910_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n53479), 
            .I2(IntegralLimit[21]), .I3(n51732), .O(n51392));
    defparam i35910_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i36634_4_lut (.I0(n24_adj_4601), .I1(n8_adj_4603), .I2(n53455), 
            .I3(n51390), .O(n52117));   // verilog/motorControl.v(31[10:34])
    defparam i36634_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36629_3_lut (.I0(n52132), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n52112));   // verilog/motorControl.v(31[10:34])
    defparam i36629_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3723 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4604), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4605));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i36676_3_lut (.I0(n4_adj_4605), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n52159));   // verilog/motorControl.v(31[38:63])
    defparam i36676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36677_3_lut (.I0(n52159), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4606), .I3(GND_net), .O(n52160));   // verilog/motorControl.v(31[38:63])
    defparam i36677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4607));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i36202_2_lut (.I0(n33), .I1(n15_adj_4608), .I2(GND_net), .I3(GND_net), 
            .O(n51684));
    defparam i36202_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4609), .I3(GND_net), 
            .O(n10_adj_4610));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4607), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4611), .I3(GND_net), 
            .O(n30_adj_4612));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i36204_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4606), .I3(n51690), 
            .O(n51686));
    defparam i36204_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36756_4_lut (.I0(n30_adj_4612), .I1(n10_adj_4610), .I2(n35_adj_4611), 
            .I3(n51684), .O(n52239));   // verilog/motorControl.v(31[38:63])
    defparam i36756_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n40515), .O(duty_23__N_3772[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5251_4 (.CI(n40970), .I0(n13852[1]), .I1(n226), .CO(n40971));
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4613));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4614));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6375_17_lut (.I0(GND_net), .I1(n17293[14]), .I2(GND_net), 
            .I3(n40871), .O(n16749[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4616));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4617));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5251_3_lut (.I0(GND_net), .I1(n13852[0]), .I2(n153_adj_4618), 
            .I3(n40969), .O(n11990[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_22 (.CI(n40515), .I0(n106[20]), .I1(n155[20]), .CO(n40516));
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n40514), .O(duty_23__N_3772[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4619));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5251_3 (.CI(n40969), .I0(n13852[0]), .I1(n153_adj_4618), 
            .CO(n40970));
    SB_LUT4 add_5251_2_lut (.I0(GND_net), .I1(n11_adj_4620), .I2(n80), 
            .I3(GND_net), .O(n11990[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5251_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_16_lut (.I0(GND_net), .I1(n17293[13]), .I2(n1117), 
            .I3(n40870), .O(n16749[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6510_12_lut (.I0(GND_net), .I1(n19133[9]), .I2(n840), 
            .I3(n40779), .O(n18869[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4595_23_lut (.I0(GND_net), .I1(n12475[20]), .I2(GND_net), 
            .I3(n41523), .O(n10831[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4595_22_lut (.I0(GND_net), .I1(n12475[19]), .I2(GND_net), 
            .I3(n41522), .O(n10831[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_22 (.CI(n41522), .I0(n12475[19]), .I1(GND_net), 
            .CO(n41523));
    SB_LUT4 add_4595_21_lut (.I0(GND_net), .I1(n12475[18]), .I2(GND_net), 
            .I3(n41521), .O(n10831[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6510_11_lut (.I0(GND_net), .I1(n19133[8]), .I2(n767), 
            .I3(n40778), .O(n18869[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_21 (.CI(n41521), .I0(n12475[18]), .I1(GND_net), 
            .CO(n41522));
    SB_LUT4 add_4595_20_lut (.I0(GND_net), .I1(n12475[17]), .I2(GND_net), 
            .I3(n41520), .O(n10831[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_20 (.CI(n41520), .I0(n12475[17]), .I1(GND_net), 
            .CO(n41521));
    SB_LUT4 add_4595_19_lut (.I0(GND_net), .I1(n12475[16]), .I2(GND_net), 
            .I3(n41519), .O(n10831[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_19 (.CI(n41519), .I0(n12475[16]), .I1(GND_net), 
            .CO(n41520));
    SB_LUT4 add_4595_18_lut (.I0(GND_net), .I1(n12475[15]), .I2(GND_net), 
            .I3(n41518), .O(n10831[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_18 (.CI(n41518), .I0(n12475[15]), .I1(GND_net), 
            .CO(n41519));
    SB_LUT4 add_4595_17_lut (.I0(GND_net), .I1(n12475[14]), .I2(GND_net), 
            .I3(n41517), .O(n10831[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_17 (.CI(n41517), .I0(n12475[14]), .I1(GND_net), 
            .CO(n41518));
    SB_LUT4 add_4595_16_lut (.I0(GND_net), .I1(n12475[13]), .I2(n1099_adj_4621), 
            .I3(n41516), .O(n10831[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4622));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4595_16 (.CI(n41516), .I0(n12475[13]), .I1(n1099_adj_4621), 
            .CO(n41517));
    SB_LUT4 add_4595_15_lut (.I0(GND_net), .I1(n12475[12]), .I2(n1026_adj_4623), 
            .I3(n41515), .O(n10831[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_11 (.CI(n40778), .I0(n19133[8]), .I1(n767), .CO(n40779));
    SB_CARRY add_4595_15 (.CI(n41515), .I0(n12475[12]), .I1(n1026_adj_4623), 
            .CO(n41516));
    SB_LUT4 add_4595_14_lut (.I0(GND_net), .I1(n12475[11]), .I2(n953_adj_4624), 
            .I3(n41514), .O(n10831[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_14 (.CI(n41514), .I0(n12475[11]), .I1(n953_adj_4624), 
            .CO(n41515));
    SB_LUT4 add_4595_13_lut (.I0(GND_net), .I1(n12475[10]), .I2(n880_adj_4625), 
            .I3(n41513), .O(n10831[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_13 (.CI(n41513), .I0(n12475[10]), .I1(n880_adj_4625), 
            .CO(n41514));
    SB_LUT4 add_4595_12_lut (.I0(GND_net), .I1(n12475[9]), .I2(n807_adj_4626), 
            .I3(n41512), .O(n10831[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_12 (.CI(n41512), .I0(n12475[9]), .I1(n807_adj_4626), 
            .CO(n41513));
    SB_LUT4 add_6510_10_lut (.I0(GND_net), .I1(n19133[7]), .I2(n694), 
            .I3(n40777), .O(n18869[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4595_11_lut (.I0(GND_net), .I1(n12475[8]), .I2(n734_adj_4627), 
            .I3(n41511), .O(n10831[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_11 (.CI(n41511), .I0(n12475[8]), .I1(n734_adj_4627), 
            .CO(n41512));
    SB_CARRY add_6375_16 (.CI(n40870), .I0(n17293[13]), .I1(n1117), .CO(n40871));
    SB_LUT4 add_6375_15_lut (.I0(GND_net), .I1(n17293[12]), .I2(n1044), 
            .I3(n40869), .O(n16749[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_15 (.CI(n40869), .I0(n17293[12]), .I1(n1044), .CO(n40870));
    SB_LUT4 add_4595_10_lut (.I0(GND_net), .I1(n12475[7]), .I2(n661_adj_4628), 
            .I3(n41510), .O(n10831[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_10 (.CI(n40777), .I0(n19133[7]), .I1(n694), .CO(n40778));
    SB_CARRY add_5251_2 (.CI(GND_net), .I0(n11_adj_4620), .I1(n80), .CO(n40969));
    SB_LUT4 add_6510_9_lut (.I0(GND_net), .I1(n19133[6]), .I2(n621), .I3(n40776), 
            .O(n18869[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_21_lut (.I0(GND_net), .I1(n14693[18]), .I2(GND_net), 
            .I3(n40968), .O(n13852[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_9 (.CI(n40776), .I0(n19133[6]), .I1(n621), .CO(n40777));
    SB_LUT4 i36293_3_lut (.I0(n52160), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n51775));   // verilog/motorControl.v(31[38:63])
    defparam i36293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4629));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4630));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4595_10 (.CI(n41510), .I0(n12475[7]), .I1(n661_adj_4628), 
            .CO(n41511));
    SB_LUT4 add_4595_9_lut (.I0(GND_net), .I1(n12475[6]), .I2(n588_adj_4631), 
            .I3(n41509), .O(n10831[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4632));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6510_8_lut (.I0(GND_net), .I1(n19133[5]), .I2(n548), .I3(n40775), 
            .O(n18869[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4633));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6230_20_lut (.I0(GND_net), .I1(n14693[17]), .I2(GND_net), 
            .I3(n40967), .O(n13852[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4634));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6510_8 (.CI(n40775), .I0(n19133[5]), .I1(n548), .CO(n40776));
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4595_9 (.CI(n41509), .I0(n12475[6]), .I1(n588_adj_4631), 
            .CO(n41510));
    SB_CARRY add_6230_20 (.CI(n40967), .I0(n14693[17]), .I1(GND_net), 
            .CO(n40968));
    SB_LUT4 add_4595_8_lut (.I0(GND_net), .I1(n12475[5]), .I2(n515_adj_4635), 
            .I3(n41508), .O(n10831[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_19_lut (.I0(GND_net), .I1(n14693[16]), .I2(GND_net), 
            .I3(n40966), .O(n13852[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_8 (.CI(n41508), .I0(n12475[5]), .I1(n515_adj_4635), 
            .CO(n41509));
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4595_7_lut (.I0(GND_net), .I1(n12475[4]), .I2(n442_adj_4636), 
            .I3(n41507), .O(n10831[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_7 (.CI(n41507), .I0(n12475[4]), .I1(n442_adj_4636), 
            .CO(n41508));
    SB_LUT4 add_4595_6_lut (.I0(GND_net), .I1(n12475[3]), .I2(n369_adj_4637), 
            .I3(n41506), .O(n10831[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_6 (.CI(n41506), .I0(n12475[3]), .I1(n369_adj_4637), 
            .CO(n41507));
    SB_CARRY add_6230_19 (.CI(n40966), .I0(n14693[16]), .I1(GND_net), 
            .CO(n40967));
    SB_LUT4 add_6375_14_lut (.I0(GND_net), .I1(n17293[11]), .I2(n971), 
            .I3(n40868), .O(n16749[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_18_lut (.I0(GND_net), .I1(n14693[15]), .I2(GND_net), 
            .I3(n40965), .O(n13852[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_14 (.CI(n40868), .I0(n17293[11]), .I1(n971), .CO(n40869));
    SB_LUT4 add_6510_7_lut (.I0(GND_net), .I1(n19133[4]), .I2(n475), .I3(n40774), 
            .O(n18869[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_7 (.CI(n40774), .I0(n19133[4]), .I1(n475), .CO(n40775));
    SB_LUT4 add_6375_13_lut (.I0(GND_net), .I1(n17293[10]), .I2(n898), 
            .I3(n40867), .O(n16749[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_13 (.CI(n40867), .I0(n17293[10]), .I1(n898), .CO(n40868));
    SB_CARRY add_6230_18 (.CI(n40965), .I0(n14693[15]), .I1(GND_net), 
            .CO(n40966));
    SB_LUT4 add_6510_6_lut (.I0(GND_net), .I1(n19133[3]), .I2(n402), .I3(n40773), 
            .O(n18869[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_12_lut (.I0(GND_net), .I1(n17293[9]), .I2(n825), 
            .I3(n40866), .O(n16749[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_17_lut (.I0(GND_net), .I1(n14693[14]), .I2(GND_net), 
            .I3(n40964), .O(n13852[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_6 (.CI(n40773), .I0(n19133[3]), .I1(n402), .CO(n40774));
    SB_LUT4 add_6510_5_lut (.I0(GND_net), .I1(n19133[2]), .I2(n329), .I3(n40772), 
            .O(n18869[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_5 (.CI(n40772), .I0(n19133[2]), .I1(n329), .CO(n40773));
    SB_LUT4 add_6510_4_lut (.I0(GND_net), .I1(n19133[1]), .I2(n256), .I3(n40771), 
            .O(n18869[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_17 (.CI(n40964), .I0(n14693[14]), .I1(GND_net), 
            .CO(n40965));
    SB_CARRY add_6510_4 (.CI(n40771), .I0(n19133[1]), .I1(n256), .CO(n40772));
    SB_LUT4 add_6230_16_lut (.I0(GND_net), .I1(n14693[13]), .I2(n1105), 
            .I3(n40963), .O(n13852[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_16 (.CI(n40963), .I0(n14693[13]), .I1(n1105), .CO(n40964));
    SB_CARRY add_6375_12 (.CI(n40866), .I0(n17293[9]), .I1(n825), .CO(n40867));
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6375_11_lut (.I0(GND_net), .I1(n17293[8]), .I2(n752), 
            .I3(n40865), .O(n16749[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_15_lut (.I0(GND_net), .I1(n14693[12]), .I2(n1032), 
            .I3(n40962), .O(n13852[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_11 (.CI(n40865), .I0(n17293[8]), .I1(n752), .CO(n40866));
    SB_LUT4 add_4595_5_lut (.I0(GND_net), .I1(n12475[2]), .I2(n296_adj_4638), 
            .I3(n41505), .O(n10831[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_15 (.CI(n40962), .I0(n14693[12]), .I1(n1032), .CO(n40963));
    SB_CARRY add_4595_5 (.CI(n41505), .I0(n12475[2]), .I1(n296_adj_4638), 
            .CO(n41506));
    SB_LUT4 add_4595_4_lut (.I0(GND_net), .I1(n12475[1]), .I2(n223_adj_4639), 
            .I3(n41504), .O(n10831[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_14_lut (.I0(GND_net), .I1(n14693[11]), .I2(n959), 
            .I3(n40961), .O(n13852[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_10_lut (.I0(GND_net), .I1(n17293[7]), .I2(n679), 
            .I3(n40864), .O(n16749[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_10 (.CI(n40864), .I0(n17293[7]), .I1(n679), .CO(n40865));
    SB_CARRY add_4595_4 (.CI(n41504), .I0(n12475[1]), .I1(n223_adj_4639), 
            .CO(n41505));
    SB_LUT4 add_4595_3_lut (.I0(GND_net), .I1(n12475[0]), .I2(n150_adj_4640), 
            .I3(n41503), .O(n10831[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_14 (.CI(n40961), .I0(n14693[11]), .I1(n959), .CO(n40962));
    SB_CARRY add_4595_3 (.CI(n41503), .I0(n12475[0]), .I1(n150_adj_4640), 
            .CO(n41504));
    SB_LUT4 add_6230_13_lut (.I0(GND_net), .I1(n14693[10]), .I2(n886), 
            .I3(n40960), .O(n13852[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4595_2_lut (.I0(GND_net), .I1(n8_adj_4641), .I2(n77_adj_4642), 
            .I3(GND_net), .O(n10831[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_2 (.CI(GND_net), .I0(n8_adj_4641), .I1(n77_adj_4642), 
            .CO(n41503));
    SB_LUT4 add_5274_22_lut (.I0(GND_net), .I1(n14292[19]), .I2(GND_net), 
            .I3(n41502), .O(n12475[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5274_21_lut (.I0(GND_net), .I1(n14292[18]), .I2(GND_net), 
            .I3(n41501), .O(n12475[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_9_lut (.I0(GND_net), .I1(n17293[6]), .I2(n606), .I3(n40863), 
            .O(n16749[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_9 (.CI(n40863), .I0(n17293[6]), .I1(n606), .CO(n40864));
    SB_CARRY add_5274_21 (.CI(n41501), .I0(n14292[18]), .I1(GND_net), 
            .CO(n41502));
    SB_LUT4 i36831_4_lut (.I0(n51775), .I1(n52239), .I2(n35_adj_4611), 
            .I3(n51686), .O(n52314));   // verilog/motorControl.v(31[38:63])
    defparam i36831_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5274_20_lut (.I0(GND_net), .I1(n14292[17]), .I2(GND_net), 
            .I3(n41500), .O(n12475[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6510_3_lut (.I0(GND_net), .I1(n19133[0]), .I2(n183_adj_4643), 
            .I3(n40770), .O(n18869[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6375_8_lut (.I0(GND_net), .I1(n17293[5]), .I2(n533), .I3(n40862), 
            .O(n16749[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6510_3 (.CI(n40770), .I0(n19133[0]), .I1(n183_adj_4643), 
            .CO(n40771));
    SB_CARRY add_6375_8 (.CI(n40862), .I0(n17293[5]), .I1(n533), .CO(n40863));
    SB_LUT4 add_6510_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n18869[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_21 (.CI(n40514), .I0(n106[19]), .I1(n155[19]), .CO(n40515));
    SB_CARRY add_6230_13 (.CI(n40960), .I0(n14693[10]), .I1(n886), .CO(n40961));
    SB_CARRY add_5274_20 (.CI(n41500), .I0(n14292[17]), .I1(GND_net), 
            .CO(n41501));
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5274_19_lut (.I0(GND_net), .I1(n14292[16]), .I2(GND_net), 
            .I3(n41499), .O(n12475[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5274_19 (.CI(n41499), .I0(n14292[16]), .I1(GND_net), 
            .CO(n41500));
    SB_LUT4 add_5274_18_lut (.I0(GND_net), .I1(n14292[15]), .I2(GND_net), 
            .I3(n41498), .O(n12475[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6510_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n40770));
    SB_CARRY add_5274_18 (.CI(n41498), .I0(n14292[15]), .I1(GND_net), 
            .CO(n41499));
    SB_LUT4 add_5274_17_lut (.I0(GND_net), .I1(n14292[14]), .I2(GND_net), 
            .I3(n41497), .O(n12475[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_7_lut (.I0(GND_net), .I1(n17293[4]), .I2(n460), .I3(n40861), 
            .O(n16749[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_17 (.CI(n41497), .I0(n14292[14]), .I1(GND_net), 
            .CO(n41498));
    SB_LUT4 add_6230_12_lut (.I0(GND_net), .I1(n14693[9]), .I2(n813), 
            .I3(n40959), .O(n13852[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5274_16_lut (.I0(GND_net), .I1(n14292[13]), .I2(n1102_adj_4647), 
            .I3(n41496), .O(n12475[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_16 (.CI(n41496), .I0(n14292[13]), .I1(n1102_adj_4647), 
            .CO(n41497));
    SB_LUT4 add_5274_15_lut (.I0(GND_net), .I1(n14292[12]), .I2(n1029_adj_4648), 
            .I3(n41495), .O(n12475[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_15 (.CI(n41495), .I0(n14292[12]), .I1(n1029_adj_4648), 
            .CO(n41496));
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5274_14_lut (.I0(GND_net), .I1(n14292[11]), .I2(n956_adj_4649), 
            .I3(n41494), .O(n12475[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5274_14 (.CI(n41494), .I0(n14292[11]), .I1(n956_adj_4649), 
            .CO(n41495));
    SB_LUT4 add_5274_13_lut (.I0(GND_net), .I1(n14292[10]), .I2(n883_adj_4651), 
            .I3(n41493), .O(n12475[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_13 (.CI(n41493), .I0(n14292[10]), .I1(n883_adj_4651), 
            .CO(n41494));
    SB_LUT4 add_5274_12_lut (.I0(GND_net), .I1(n14292[9]), .I2(n810_adj_4652), 
            .I3(n41492), .O(n12475[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_12 (.CI(n41492), .I0(n14292[9]), .I1(n810_adj_4652), 
            .CO(n41493));
    SB_LUT4 add_5274_11_lut (.I0(GND_net), .I1(n14292[8]), .I2(n737_adj_4653), 
            .I3(n41491), .O(n12475[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_11 (.CI(n41491), .I0(n14292[8]), .I1(n737_adj_4653), 
            .CO(n41492));
    SB_LUT4 add_5274_10_lut (.I0(GND_net), .I1(n14292[7]), .I2(n664_adj_4654), 
            .I3(n41490), .O(n12475[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_12 (.CI(n40959), .I0(n14693[9]), .I1(n813), .CO(n40960));
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6375_7 (.CI(n40861), .I0(n17293[4]), .I1(n460), .CO(n40862));
    SB_CARRY add_5274_10 (.CI(n41490), .I0(n14292[7]), .I1(n664_adj_4654), 
            .CO(n41491));
    SB_LUT4 add_5274_9_lut (.I0(GND_net), .I1(n14292[6]), .I2(n591_adj_4655), 
            .I3(n41489), .O(n12475[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n40513), .O(duty_23__N_3772[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_6_lut (.I0(GND_net), .I1(n17293[3]), .I2(n387), .I3(n40860), 
            .O(n16749[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_11_lut (.I0(GND_net), .I1(n14693[8]), .I2(n740), 
            .I3(n40958), .O(n13852[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_11 (.CI(n40958), .I0(n14693[8]), .I1(n740), .CO(n40959));
    SB_CARRY add_5274_9 (.CI(n41489), .I0(n14292[6]), .I1(n591_adj_4655), 
            .CO(n41490));
    SB_LUT4 add_5274_8_lut (.I0(GND_net), .I1(n14292[5]), .I2(n518_adj_4656), 
            .I3(n41488), .O(n12475[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_10_lut (.I0(GND_net), .I1(n14693[7]), .I2(n667), 
            .I3(n40957), .O(n13852[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_10 (.CI(n40957), .I0(n14693[7]), .I1(n667), .CO(n40958));
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6230_9_lut (.I0(GND_net), .I1(n14693[6]), .I2(n594), .I3(n40956), 
            .O(n13852[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_8 (.CI(n41488), .I0(n14292[5]), .I1(n518_adj_4656), 
            .CO(n41489));
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6375_6 (.CI(n40860), .I0(n17293[3]), .I1(n387), .CO(n40861));
    SB_LUT4 add_5274_7_lut (.I0(GND_net), .I1(n14292[4]), .I2(n445_adj_4657), 
            .I3(n41487), .O(n12475[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_9 (.CI(n40956), .I0(n14693[6]), .I1(n594), .CO(n40957));
    SB_CARRY add_5274_7 (.CI(n41487), .I0(n14292[4]), .I1(n445_adj_4657), 
            .CO(n41488));
    SB_CARRY add_12_20 (.CI(n40513), .I0(n106[18]), .I1(n155[18]), .CO(n40514));
    SB_LUT4 add_5274_6_lut (.I0(GND_net), .I1(n14292[3]), .I2(n372_adj_4658), 
            .I3(n41486), .O(n12475[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_6 (.CI(n41486), .I0(n14292[3]), .I1(n372_adj_4658), 
            .CO(n41487));
    SB_LUT4 add_5274_5_lut (.I0(GND_net), .I1(n14292[2]), .I2(n299_adj_4659), 
            .I3(n41485), .O(n12475[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_5 (.CI(n41485), .I0(n14292[2]), .I1(n299_adj_4659), 
            .CO(n41486));
    SB_LUT4 i36832_3_lut (.I0(n52314), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n52315));   // verilog/motorControl.v(31[38:63])
    defparam i36832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36816_3_lut (.I0(n52315), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n52299));   // verilog/motorControl.v(31[38:63])
    defparam i36816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4660), .I3(GND_net), 
            .O(n6_adj_4661));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i36626_3_lut (.I0(n6_adj_4661), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4662), .I3(GND_net), .O(n52109));   // verilog/motorControl.v(31[38:63])
    defparam i36626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36627_3_lut (.I0(n52109), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4663), .I3(GND_net), .O(n52110));   // verilog/motorControl.v(31[38:63])
    defparam i36627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36193_4_lut (.I0(n43), .I1(n25_adj_4664), .I2(n23_adj_4663), 
            .I3(n51697), .O(n51675));
    defparam i36193_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36636_4_lut (.I0(n24_adj_4569), .I1(n8_adj_4557), .I2(n45), 
            .I3(n51673), .O(n52119));   // verilog/motorControl.v(31[38:63])
    defparam i36636_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36291_3_lut (.I0(n52110), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4664), .I3(GND_net), .O(n51773));   // verilog/motorControl.v(31[38:63])
    defparam i36291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36195_4_lut (.I0(n43), .I1(n41_adj_4665), .I2(n39), .I3(n52274), 
            .O(n51677));
    defparam i36195_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36774_4_lut (.I0(n51773), .I1(n52119), .I2(n45), .I3(n51675), 
            .O(n52257));   // verilog/motorControl.v(31[38:63])
    defparam i36774_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36299_3_lut (.I0(n52299), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4665), .I3(GND_net), .O(n51781));   // verilog/motorControl.v(31[38:63])
    defparam i36299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36776_4_lut (.I0(n51781), .I1(n52257), .I2(n45), .I3(n51677), 
            .O(n52259));   // verilog/motorControl.v(31[38:63])
    defparam i36776_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4666));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i36646_3_lut (.I0(n4_adj_4666), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n52129));   // verilog/motorControl.v(31[10:34])
    defparam i36646_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36647_3_lut (.I0(n52129), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n52130));   // verilog/motorControl.v(31[10:34])
    defparam i36647_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35921_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n53465), 
            .I2(IntegralLimit[16]), .I3(n51726), .O(n51403));
    defparam i35921_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i36799_4_lut (.I0(n30), .I1(n10_adj_4555), .I2(n53489), .I3(n51401), 
            .O(n52282));   // verilog/motorControl.v(31[10:34])
    defparam i36799_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36631_3_lut (.I0(n52130), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n52114));   // verilog/motorControl.v(31[10:34])
    defparam i36631_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36837_4_lut (.I0(n52114), .I1(n52282), .I2(n53489), .I3(n51403), 
            .O(n52320));   // verilog/motorControl.v(31[10:34])
    defparam i36837_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36838_3_lut (.I0(n52320), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n52321));   // verilog/motorControl.v(31[10:34])
    defparam i36838_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36810_3_lut (.I0(n52321), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n52293));   // verilog/motorControl.v(31[10:34])
    defparam i36810_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5274_4_lut (.I0(GND_net), .I1(n14292[1]), .I2(n226_adj_4667), 
            .I3(n41484), .O(n12475[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_4 (.CI(n41484), .I0(n14292[1]), .I1(n226_adj_4667), 
            .CO(n41485));
    SB_LUT4 add_6230_8_lut (.I0(GND_net), .I1(n14693[5]), .I2(n521), .I3(n40955), 
            .O(n13852[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5274_3_lut (.I0(GND_net), .I1(n14292[0]), .I2(n153_adj_4668), 
            .I3(n41483), .O(n12475[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_3 (.CI(n41483), .I0(n14292[0]), .I1(n153_adj_4668), 
            .CO(n41484));
    SB_LUT4 add_5274_2_lut (.I0(GND_net), .I1(n11_adj_4669), .I2(n80_adj_4670), 
            .I3(GND_net), .O(n12475[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5274_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5274_2 (.CI(GND_net), .I0(n11_adj_4669), .I1(n80_adj_4670), 
            .CO(n41483));
    SB_LUT4 add_6250_21_lut (.I0(GND_net), .I1(n15092[18]), .I2(GND_net), 
            .I3(n41482), .O(n14292[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n40512), .O(duty_23__N_3772[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_5_lut (.I0(GND_net), .I1(n17293[2]), .I2(n314), .I3(n40859), 
            .O(n16749[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_20_lut (.I0(GND_net), .I1(n15092[17]), .I2(GND_net), 
            .I3(n41481), .O(n14292[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_8 (.CI(n40955), .I0(n14693[5]), .I1(n521), .CO(n40956));
    SB_CARRY add_12_19 (.CI(n40512), .I0(n106[17]), .I1(n155[17]), .CO(n40513));
    SB_CARRY add_6375_5 (.CI(n40859), .I0(n17293[2]), .I1(n314), .CO(n40860));
    SB_CARRY add_6250_20 (.CI(n41481), .I0(n15092[17]), .I1(GND_net), 
            .CO(n41482));
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35912_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n53457), 
            .I2(IntegralLimit[21]), .I3(n52278), .O(n51394));
    defparam i35912_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_129_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n53455));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_129_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36724_4_lut (.I0(n52112), .I1(n52117), .I2(n53455), .I3(n51392), 
            .O(n52207));   // verilog/motorControl.v(31[10:34])
    defparam i36724_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_6250_19_lut (.I0(GND_net), .I1(n15092[16]), .I2(GND_net), 
            .I3(n41480), .O(n14292[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_7_lut (.I0(GND_net), .I1(n14693[4]), .I2(n448), .I3(n40954), 
            .O(n13852[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_7 (.CI(n40954), .I0(n14693[4]), .I1(n448), .CO(n40955));
    SB_LUT4 add_6375_4_lut (.I0(GND_net), .I1(n17293[1]), .I2(n241), .I3(n40858), 
            .O(n16749[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36808_3_lut (.I0(n52293), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(31[10:34])
    defparam i36808_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36777_3_lut (.I0(n52259), .I1(\PID_CONTROLLER.integral_23__N_3723 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3722 ));   // verilog/motorControl.v(31[38:63])
    defparam i36777_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36726_4_lut (.I0(n40), .I1(n52207), .I2(n53455), .I3(n51394), 
            .O(n52209));   // verilog/motorControl.v(31[10:34])
    defparam i36726_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_6250_19 (.CI(n41480), .I0(n15092[16]), .I1(GND_net), 
            .CO(n41481));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_850_4_lut  (.I0(n52209), .I1(\PID_CONTROLLER.integral_23__N_3722 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3720 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_850_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22015_2_lut (.I0(n1[12]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22015_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6250_18_lut (.I0(GND_net), .I1(n15092[15]), .I2(GND_net), 
            .I3(n41479), .O(n14292[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_4 (.CI(n40858), .I0(n17293[1]), .I1(n241), .CO(n40859));
    SB_LUT4 add_6375_3_lut (.I0(GND_net), .I1(n17293[0]), .I2(n168), .I3(n40857), 
            .O(n16749[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_18 (.CI(n41479), .I0(n15092[15]), .I1(GND_net), 
            .CO(n41480));
    SB_LUT4 add_6230_6_lut (.I0(GND_net), .I1(n14693[3]), .I2(n375), .I3(n40953), 
            .O(n13852[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_17_lut (.I0(GND_net), .I1(n15092[14]), .I2(GND_net), 
            .I3(n41478), .O(n14292[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n40511), .O(duty_23__N_3772[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_3 (.CI(n40857), .I0(n17293[0]), .I1(n168), .CO(n40858));
    SB_CARRY add_6250_17 (.CI(n41478), .I0(n15092[14]), .I1(GND_net), 
            .CO(n41479));
    SB_LUT4 add_6250_16_lut (.I0(GND_net), .I1(n15092[13]), .I2(n1105_adj_4671), 
            .I3(n41477), .O(n14292[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_18 (.CI(n40511), .I0(n106[16]), .I1(n155[16]), .CO(n40512));
    SB_CARRY add_6250_16 (.CI(n41477), .I0(n15092[13]), .I1(n1105_adj_4671), 
            .CO(n41478));
    SB_CARRY add_6230_6 (.CI(n40953), .I0(n14693[3]), .I1(n375), .CO(n40954));
    SB_LUT4 add_6230_5_lut (.I0(GND_net), .I1(n14693[2]), .I2(n302), .I3(n40952), 
            .O(n13852[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_15_lut (.I0(GND_net), .I1(n15092[12]), .I2(n1032_adj_4672), 
            .I3(n41476), .O(n14292[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_5 (.CI(n40952), .I0(n14693[2]), .I1(n302), .CO(n40953));
    SB_CARRY add_6250_15 (.CI(n41476), .I0(n15092[12]), .I1(n1032_adj_4672), 
            .CO(n41477));
    SB_LUT4 add_6250_14_lut (.I0(GND_net), .I1(n15092[11]), .I2(n959_adj_4673), 
            .I3(n41475), .O(n14292[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_4_lut (.I0(GND_net), .I1(n14693[1]), .I2(n229), .I3(n40951), 
            .O(n13852[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_14 (.CI(n41475), .I0(n15092[11]), .I1(n959_adj_4673), 
            .CO(n41476));
    SB_LUT4 add_6250_13_lut (.I0(GND_net), .I1(n15092[10]), .I2(n886_adj_4674), 
            .I3(n41474), .O(n14292[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_13 (.CI(n41474), .I0(n15092[10]), .I1(n886_adj_4674), 
            .CO(n41475));
    SB_LUT4 add_6250_12_lut (.I0(GND_net), .I1(n15092[9]), .I2(n813_adj_4675), 
            .I3(n41473), .O(n14292[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n40510), .O(duty_23__N_3772[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_4 (.CI(n40951), .I0(n14693[1]), .I1(n229), .CO(n40952));
    SB_CARRY add_6250_12 (.CI(n41473), .I0(n15092[9]), .I1(n813_adj_4675), 
            .CO(n41474));
    SB_LUT4 add_6230_3_lut (.I0(GND_net), .I1(n14693[0]), .I2(n156), .I3(n40950), 
            .O(n13852[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_2_lut (.I0(GND_net), .I1(n26_adj_4676), .I2(n95), 
            .I3(GND_net), .O(n16749[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_2 (.CI(GND_net), .I0(n26_adj_4676), .I1(n95), .CO(n40857));
    SB_CARRY add_6230_3 (.CI(n40950), .I0(n14693[0]), .I1(n156), .CO(n40951));
    SB_LUT4 add_6230_2_lut (.I0(GND_net), .I1(n14_adj_4677), .I2(n83), 
            .I3(GND_net), .O(n13852[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6575_9_lut (.I0(GND_net), .I1(n19740[6]), .I2(n630_adj_4678), 
            .I3(n40856), .O(n19613[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6575_8_lut (.I0(GND_net), .I1(n19740[5]), .I2(n557_adj_4679), 
            .I3(n40855), .O(n19613[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3772[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4680));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3772[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4681));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3772[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4682));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6230_2 (.CI(GND_net), .I0(n14_adj_4677), .I1(n83), .CO(n40950));
    SB_LUT4 duty_23__I_851_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3772[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4683));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3772[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4684));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3772[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4685));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4686));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6541_11_lut (.I0(GND_net), .I1(n19452[8]), .I2(n770), 
            .I3(n40949), .O(n19253[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3772[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4687));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3772[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4688));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3772[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4689));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3772[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4690));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3772[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4691));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3772[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4692));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3772[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4693));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6541_10_lut (.I0(GND_net), .I1(n19452[7]), .I2(n697), 
            .I3(n40948), .O(n19253[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_11_lut (.I0(GND_net), .I1(n15092[8]), .I2(n740_adj_4695), 
            .I3(n41472), .O(n14292[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_11 (.CI(n41472), .I0(n15092[8]), .I1(n740_adj_4695), 
            .CO(n41473));
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4696));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6541_10 (.CI(n40948), .I0(n19452[7]), .I1(n697), .CO(n40949));
    SB_LUT4 add_6250_10_lut (.I0(GND_net), .I1(n15092[7]), .I2(n667_adj_4697), 
            .I3(n41471), .O(n14292[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6541_9_lut (.I0(GND_net), .I1(n19452[6]), .I2(n624), .I3(n40947), 
            .O(n19253[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_9 (.CI(n40947), .I0(n19452[6]), .I1(n624), .CO(n40948));
    SB_CARRY add_12_17 (.CI(n40510), .I0(n106[15]), .I1(n155[15]), .CO(n40511));
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_851_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4699));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3772[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4700));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6250_10 (.CI(n41471), .I0(n15092[7]), .I1(n667_adj_4697), 
            .CO(n41472));
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6250_9_lut (.I0(GND_net), .I1(n15092[6]), .I2(n594_adj_4701), 
            .I3(n41470), .O(n14292[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_9 (.CI(n41470), .I0(n15092[6]), .I1(n594_adj_4701), 
            .CO(n41471));
    SB_LUT4 duty_23__I_851_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3772[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4702));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6250_8_lut (.I0(GND_net), .I1(n15092[5]), .I2(n521_adj_4703), 
            .I3(n41469), .O(n14292[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6541_8_lut (.I0(GND_net), .I1(n19452[5]), .I2(n551), .I3(n40946), 
            .O(n19253[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3772[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4704));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36154_3_lut_4_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3772[2]), .O(n51636));   // verilog/motorControl.v(38[19:35])
    defparam i36154_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_6541_8 (.CI(n40946), .I0(n19452[5]), .I1(n551), .CO(n40947));
    SB_CARRY add_6250_8 (.CI(n41469), .I0(n15092[5]), .I1(n521_adj_4703), 
            .CO(n41470));
    SB_LUT4 add_6541_7_lut (.I0(GND_net), .I1(n19452[4]), .I2(n478), .I3(n40945), 
            .O(n19253[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_7_lut (.I0(GND_net), .I1(n15092[4]), .I2(n448_adj_4705), 
            .I3(n41468), .O(n14292[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3772[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4706));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6250_7 (.CI(n41468), .I0(n15092[4]), .I1(n448_adj_4705), 
            .CO(n41469));
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4707));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6250_6_lut (.I0(GND_net), .I1(n15092[3]), .I2(n375_adj_4708), 
            .I3(n41467), .O(n14292[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_6 (.CI(n41467), .I0(n15092[3]), .I1(n375_adj_4708), 
            .CO(n41468));
    SB_LUT4 i36178_4_lut (.I0(n21_adj_4706), .I1(n19_adj_4704), .I2(n17_adj_4702), 
            .I3(n9_adj_4700), .O(n51660));
    defparam i36178_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4709));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4710));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36172_4_lut (.I0(n27_adj_4693), .I1(n15_adj_4692), .I2(n13_adj_4691), 
            .I3(n11_adj_4690), .O(n51654));
    defparam i36172_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4711));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i12_3_lut (.I0(duty_23__N_3772[7]), .I1(duty_23__N_3772[16]), 
            .I2(n33_adj_4699), .I3(GND_net), .O(n12_adj_4712));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6250_5_lut (.I0(GND_net), .I1(n15092[2]), .I2(n302_adj_4713), 
            .I3(n41466), .O(n14292[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_5 (.CI(n41466), .I0(n15092[2]), .I1(n302_adj_4713), 
            .CO(n41467));
    SB_CARRY add_6575_8 (.CI(n40855), .I0(n19740[5]), .I1(n557_adj_4679), 
            .CO(n40856));
    SB_LUT4 duty_23__I_851_i10_3_lut (.I0(duty_23__N_3772[5]), .I1(duty_23__N_3772[6]), 
            .I2(n13_adj_4691), .I3(GND_net), .O(n10_adj_4714));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i30_3_lut (.I0(n12_adj_4712), .I1(duty_23__N_3772[17]), 
            .I2(n35_adj_4689), .I3(GND_net), .O(n30_adj_4715));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6250_4_lut (.I0(GND_net), .I1(n15092[1]), .I2(n229_adj_4716), 
            .I3(n41465), .O(n14292[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_4 (.CI(n41465), .I0(n15092[1]), .I1(n229_adj_4716), 
            .CO(n41466));
    SB_CARRY add_6541_7 (.CI(n40945), .I0(n19452[4]), .I1(n478), .CO(n40946));
    SB_LUT4 add_6541_6_lut (.I0(GND_net), .I1(n19452[3]), .I2(n405), .I3(n40944), 
            .O(n19253[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36422_4_lut (.I0(n13_adj_4691), .I1(n11_adj_4690), .I2(n9_adj_4700), 
            .I3(n51671), .O(n51905));
    defparam i36422_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_6250_3_lut (.I0(GND_net), .I1(n15092[0]), .I2(n156_adj_4717), 
            .I3(n41464), .O(n14292[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36418_4_lut (.I0(n19_adj_4704), .I1(n17_adj_4702), .I2(n15_adj_4692), 
            .I3(n51905), .O(n51901));
    defparam i36418_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_6250_3 (.CI(n41464), .I0(n15092[0]), .I1(n156_adj_4717), 
            .CO(n41465));
    SB_LUT4 i36748_4_lut (.I0(n25_adj_4685), .I1(n23_adj_4684), .I2(n21_adj_4706), 
            .I3(n51901), .O(n52231));
    defparam i36748_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36570_4_lut (.I0(n31_adj_4688), .I1(n29_adj_4687), .I2(n27_adj_4693), 
            .I3(n52231), .O(n52053));
    defparam i36570_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36789_4_lut (.I0(n37_adj_4683), .I1(n35_adj_4689), .I2(n33_adj_4699), 
            .I3(n52053), .O(n52272));
    defparam i36789_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 duty_23__I_851_i16_3_lut (.I0(duty_23__N_3772[9]), .I1(duty_23__N_3772[21]), 
            .I2(n43_adj_4686), .I3(GND_net), .O(n16_adj_4718));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6250_2_lut (.I0(GND_net), .I1(n14_adj_4719), .I2(n83_adj_4720), 
            .I3(GND_net), .O(n14292[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36672_3_lut (.I0(n6_adj_4721), .I1(duty_23__N_3772[10]), .I2(n21_adj_4706), 
            .I3(GND_net), .O(n52155));   // verilog/motorControl.v(36[10:25])
    defparam i36672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36673_3_lut (.I0(n52155), .I1(duty_23__N_3772[11]), .I2(n23_adj_4684), 
            .I3(GND_net), .O(n52156));   // verilog/motorControl.v(36[10:25])
    defparam i36673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4722));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6541_6 (.CI(n40944), .I0(n19452[3]), .I1(n405), .CO(n40945));
    SB_LUT4 duty_23__I_851_i8_3_lut (.I0(duty_23__N_3772[4]), .I1(duty_23__N_3772[8]), 
            .I2(n17_adj_4702), .I3(GND_net), .O(n8_adj_4723));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i24_3_lut (.I0(n16_adj_4718), .I1(duty_23__N_3772[22]), 
            .I2(n45_adj_4682), .I3(GND_net), .O(n24_adj_4724));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4725));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6575_7_lut (.I0(GND_net), .I1(n19740[4]), .I2(n484_adj_4727), 
            .I3(n40854), .O(n19613[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_2 (.CI(GND_net), .I0(n14_adj_4719), .I1(n83_adj_4720), 
            .CO(n41464));
    SB_LUT4 add_6289_20_lut (.I0(GND_net), .I1(n15813[17]), .I2(GND_net), 
            .I3(n41463), .O(n15092[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4728));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4729));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36158_4_lut (.I0(n43_adj_4686), .I1(n25_adj_4685), .I2(n23_adj_4684), 
            .I3(n51660), .O(n51640));
    defparam i36158_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4731));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4732));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4733));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36638_4_lut (.I0(n24_adj_4724), .I1(n8_adj_4723), .I2(n45_adj_4682), 
            .I3(n51638), .O(n52121));   // verilog/motorControl.v(36[10:25])
    defparam i36638_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36301_3_lut (.I0(n52156), .I1(duty_23__N_3772[12]), .I2(n25_adj_4685), 
            .I3(GND_net), .O(n51783));   // verilog/motorControl.v(36[10:25])
    defparam i36301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(duty_23__N_3772[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4734));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 add_6541_5_lut (.I0(GND_net), .I1(n19452[2]), .I2(n332), .I3(n40943), 
            .O(n19253[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36670_3_lut (.I0(n4_adj_4734), .I1(duty_23__N_3772[13]), .I2(n27_adj_4693), 
            .I3(GND_net), .O(n52153));   // verilog/motorControl.v(36[10:25])
    defparam i36670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36671_3_lut (.I0(n52153), .I1(duty_23__N_3772[14]), .I2(n29_adj_4687), 
            .I3(GND_net), .O(n52154));   // verilog/motorControl.v(36[10:25])
    defparam i36671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36168_4_lut (.I0(n33_adj_4699), .I1(n31_adj_4688), .I2(n29_adj_4687), 
            .I3(n51654), .O(n51650));
    defparam i36168_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36758_4_lut (.I0(n30_adj_4715), .I1(n10_adj_4714), .I2(n35_adj_4689), 
            .I3(n51648), .O(n52241));   // verilog/motorControl.v(36[10:25])
    defparam i36758_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_6575_7 (.CI(n40854), .I0(n19740[4]), .I1(n484_adj_4727), 
            .CO(n40855));
    SB_LUT4 i36303_3_lut (.I0(n52154), .I1(duty_23__N_3772[15]), .I2(n31_adj_4688), 
            .I3(GND_net), .O(n51785));   // verilog/motorControl.v(36[10:25])
    defparam i36303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36833_4_lut (.I0(n51785), .I1(n52241), .I2(n35_adj_4689), 
            .I3(n51650), .O(n52316));   // verilog/motorControl.v(36[10:25])
    defparam i36833_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36834_3_lut (.I0(n52316), .I1(duty_23__N_3772[18]), .I2(n37_adj_4683), 
            .I3(GND_net), .O(n52317));   // verilog/motorControl.v(36[10:25])
    defparam i36834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4735));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36814_3_lut (.I0(n52317), .I1(duty_23__N_3772[19]), .I2(n39_adj_4680), 
            .I3(GND_net), .O(n52297));   // verilog/motorControl.v(36[10:25])
    defparam i36814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36160_4_lut (.I0(n43_adj_4686), .I1(n41_adj_4681), .I2(n39_adj_4680), 
            .I3(n52272), .O(n51642));
    defparam i36160_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36189_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(PWMLimit[2]), .O(n51671));   // verilog/motorControl.v(36[10:25])
    defparam i36189_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n40509), .O(duty_23__N_3772[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36778_4_lut (.I0(n51783), .I1(n52121), .I2(n45_adj_4682), 
            .I3(n51640), .O(n52261));   // verilog/motorControl.v(36[10:25])
    defparam i36778_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_6289_19_lut (.I0(GND_net), .I1(n15813[16]), .I2(GND_net), 
            .I3(n41462), .O(n15092[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36309_3_lut (.I0(n52297), .I1(duty_23__N_3772[20]), .I2(n41_adj_4681), 
            .I3(GND_net), .O(n51791));   // verilog/motorControl.v(36[10:25])
    defparam i36309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36780_4_lut (.I0(n51791), .I1(n52261), .I2(n45_adj_4682), 
            .I3(n51642), .O(n52263));   // verilog/motorControl.v(36[10:25])
    defparam i36780_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4737));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4738));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36781_3_lut (.I0(n52263), .I1(PWMLimit[23]), .I2(duty_23__N_3772[23]), 
            .I3(GND_net), .O(duty_23__N_3771));   // verilog/motorControl.v(36[10:25])
    defparam i36781_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36791_4_lut (.I0(n37), .I1(n35_adj_4611), .I2(n33), .I3(n52069), 
            .O(n52274));
    defparam i36791_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4739));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36586_4_lut (.I0(n31), .I1(n29_adj_4606), .I2(n27), .I3(n52177), 
            .O(n52069));
    defparam i36586_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4741));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4742));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4743));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4744));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4745));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4747));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4748));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4749));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4750));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4752));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4753));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4754));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4755));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4756));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4757));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4758));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6289_19 (.CI(n41462), .I0(n15813[16]), .I1(GND_net), 
            .CO(n41463));
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4759));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_12_16 (.CI(n40509), .I0(n106[14]), .I1(n155[14]), .CO(n40510));
    SB_LUT4 add_6289_18_lut (.I0(GND_net), .I1(n15813[15]), .I2(GND_net), 
            .I3(n41461), .O(n15092[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4760));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4762));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4763));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4765));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4766));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4768));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4769));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4771));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4772));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6289_18 (.CI(n41461), .I0(n15813[15]), .I1(GND_net), 
            .CO(n41462));
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4774));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6289_17_lut (.I0(GND_net), .I1(n15813[14]), .I2(GND_net), 
            .I3(n41460), .O(n15092[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4776));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6575_6_lut (.I0(GND_net), .I1(n19740[3]), .I2(n411_adj_4777), 
            .I3(n40853), .O(n19613[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36142_4_lut (.I0(n21_adj_4768), .I1(n19_adj_4766), .I2(n17_adj_4765), 
            .I3(n9_adj_4763), .O(n51624));
    defparam i36142_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6289_17 (.CI(n41460), .I0(n15813[14]), .I1(GND_net), 
            .CO(n41461));
    SB_LUT4 i36136_4_lut (.I0(n27_adj_4776), .I1(n15_adj_4774), .I2(n13_adj_4772), 
            .I3(n11_adj_4771), .O(n51618));
    defparam i36136_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n40508), .O(duty_23__N_3772[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_15 (.CI(n40508), .I0(n106[13]), .I1(n155[13]), .CO(n40509));
    SB_CARRY add_6541_5 (.CI(n40943), .I0(n19452[2]), .I1(n332), .CO(n40944));
    SB_LUT4 add_6289_16_lut (.I0(GND_net), .I1(n15813[13]), .I2(n1108), 
            .I3(n41459), .O(n15092[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_16 (.CI(n41459), .I0(n15813[13]), .I1(n1108), .CO(n41460));
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4762), 
            .I3(GND_net), .O(n12_adj_4778));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4779));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6289_15_lut (.I0(GND_net), .I1(n15813[12]), .I2(n1035), 
            .I3(n41458), .O(n15092[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_15 (.CI(n41458), .I0(n15813[12]), .I1(n1035), .CO(n41459));
    SB_CARRY add_6575_6 (.CI(n40853), .I0(n19740[3]), .I1(n411_adj_4777), 
            .CO(n40854));
    SB_LUT4 add_6541_4_lut (.I0(GND_net), .I1(n19452[1]), .I2(n259_adj_4780), 
            .I3(n40942), .O(n19253[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4781));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6289_14_lut (.I0(GND_net), .I1(n15813[11]), .I2(n962), 
            .I3(n41457), .O(n15092[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_14 (.CI(n41457), .I0(n15813[11]), .I1(n962), .CO(n41458));
    SB_LUT4 add_6575_5_lut (.I0(GND_net), .I1(n19740[2]), .I2(n338_adj_4782), 
            .I3(n40852), .O(n19613[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_13_lut (.I0(GND_net), .I1(n15813[10]), .I2(n889_adj_4783), 
            .I3(n41456), .O(n15092[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_4 (.CI(n40942), .I0(n19452[1]), .I1(n259_adj_4780), 
            .CO(n40943));
    SB_CARRY add_6289_13 (.CI(n41456), .I0(n15813[10]), .I1(n889_adj_4783), 
            .CO(n41457));
    SB_LUT4 add_6541_3_lut (.I0(GND_net), .I1(n19452[0]), .I2(n186_adj_4784), 
            .I3(n40941), .O(n19253[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n40507), .O(duty_23__N_3772[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6575_5 (.CI(n40852), .I0(n19740[2]), .I1(n338_adj_4782), 
            .CO(n40853));
    SB_LUT4 add_6289_12_lut (.I0(GND_net), .I1(n15813[9]), .I2(n816_adj_4785), 
            .I3(n41455), .O(n15092[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4786));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6289_12 (.CI(n41455), .I0(n15813[9]), .I1(n816_adj_4785), 
            .CO(n41456));
    SB_LUT4 add_6289_11_lut (.I0(GND_net), .I1(n15813[8]), .I2(n743_adj_4787), 
            .I3(n41454), .O(n15092[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4772), 
            .I3(GND_net), .O(n10_adj_4788));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6541_3 (.CI(n40941), .I0(n19452[0]), .I1(n186_adj_4784), 
            .CO(n40942));
    SB_CARRY add_6289_11 (.CI(n41454), .I0(n15813[8]), .I1(n743_adj_4787), 
            .CO(n41455));
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4778), .I1(n257[17]), .I2(n35_adj_4760), 
            .I3(GND_net), .O(n30_adj_4789));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6289_10_lut (.I0(GND_net), .I1(n15813[7]), .I2(n670_adj_4790), 
            .I3(n41453), .O(n15092[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_10 (.CI(n41453), .I0(n15813[7]), .I1(n670_adj_4790), 
            .CO(n41454));
    SB_LUT4 add_6575_4_lut (.I0(GND_net), .I1(n19740[1]), .I2(n265_adj_4791), 
            .I3(n40851), .O(n19613[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36390_4_lut (.I0(n13_adj_4772), .I1(n11_adj_4771), .I2(n9_adj_4763), 
            .I3(n51636), .O(n51873));
    defparam i36390_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_6289_9_lut (.I0(GND_net), .I1(n15813[6]), .I2(n597_adj_4792), 
            .I3(n41452), .O(n15092[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36386_4_lut (.I0(n19_adj_4766), .I1(n17_adj_4765), .I2(n15_adj_4774), 
            .I3(n51873), .O(n51869));
    defparam i36386_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_6541_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n19253[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n40941));
    SB_CARRY add_6289_9 (.CI(n41452), .I0(n15813[6]), .I1(n597_adj_4792), 
            .CO(n41453));
    SB_LUT4 add_6270_20_lut (.I0(GND_net), .I1(n15453[17]), .I2(GND_net), 
            .I3(n40940), .O(n14693[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n40507), .I0(n106[12]), .I1(n155[12]), .CO(n40508));
    SB_LUT4 add_6289_8_lut (.I0(GND_net), .I1(n15813[5]), .I2(n524_adj_4793), 
            .I3(n41451), .O(n15092[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_8 (.CI(n41451), .I0(n15813[5]), .I1(n524_adj_4793), 
            .CO(n41452));
    SB_CARRY add_6575_4 (.CI(n40851), .I0(n19740[1]), .I1(n265_adj_4791), 
            .CO(n40852));
    SB_LUT4 add_6289_7_lut (.I0(GND_net), .I1(n15813[4]), .I2(n451_adj_4794), 
            .I3(n41450), .O(n15092[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6270_19_lut (.I0(GND_net), .I1(n15453[16]), .I2(GND_net), 
            .I3(n40939), .O(n14693[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_7 (.CI(n41450), .I0(n15813[4]), .I1(n451_adj_4794), 
            .CO(n41451));
    SB_LUT4 add_6289_6_lut (.I0(GND_net), .I1(n15813[3]), .I2(n378_adj_4795), 
            .I3(n41449), .O(n15092[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6575_3_lut (.I0(GND_net), .I1(n19740[0]), .I2(n192_adj_4796), 
            .I3(n40850), .O(n19613[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n40506), .O(duty_23__N_3772[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6575_3 (.CI(n40850), .I0(n19740[0]), .I1(n192_adj_4796), 
            .CO(n40851));
    SB_CARRY add_6289_6 (.CI(n41449), .I0(n15813[3]), .I1(n378_adj_4795), 
            .CO(n41450));
    SB_LUT4 add_6575_2_lut (.I0(GND_net), .I1(n50_adj_4798), .I2(n119_adj_4799), 
            .I3(GND_net), .O(n19613[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_5_lut (.I0(GND_net), .I1(n15813[2]), .I2(n305_adj_4800), 
            .I3(n41448), .O(n15092[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36742_4_lut (.I0(n25_adj_4759), .I1(n23_adj_4758), .I2(n21_adj_4768), 
            .I3(n51869), .O(n52225));
    defparam i36742_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_6289_5 (.CI(n41448), .I0(n15813[2]), .I1(n305_adj_4800), 
            .CO(n41449));
    SB_CARRY add_6575_2 (.CI(GND_net), .I0(n50_adj_4798), .I1(n119_adj_4799), 
            .CO(n40850));
    SB_LUT4 add_6289_4_lut (.I0(GND_net), .I1(n15813[1]), .I2(n232_adj_4801), 
            .I3(n41447), .O(n15092[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_19 (.CI(n40939), .I0(n15453[16]), .I1(GND_net), 
            .CO(n40940));
    SB_CARRY add_6289_4 (.CI(n41447), .I0(n15813[1]), .I1(n232_adj_4801), 
            .CO(n41448));
    SB_LUT4 i36554_4_lut (.I0(n31_adj_4752), .I1(n29_adj_4749), .I2(n27_adj_4776), 
            .I3(n52225), .O(n52037));
    defparam i36554_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_6289_3_lut (.I0(GND_net), .I1(n15813[0]), .I2(n159_adj_4802), 
            .I3(n41446), .O(n15092[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_3 (.CI(n41446), .I0(n15813[0]), .I1(n159_adj_4802), 
            .CO(n41447));
    SB_LUT4 add_6270_18_lut (.I0(GND_net), .I1(n15453[15]), .I2(GND_net), 
            .I3(n40938), .O(n14693[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_13 (.CI(n40506), .I0(n106[11]), .I1(n155[11]), .CO(n40507));
    SB_LUT4 add_6406_16_lut (.I0(GND_net), .I1(n17773[13]), .I2(n1120_adj_4803), 
            .I3(n40849), .O(n17293[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n40505), .O(duty_23__N_3772[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_2_lut (.I0(GND_net), .I1(n17_adj_4804), .I2(n86_adj_4805), 
            .I3(GND_net), .O(n15092[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_2 (.CI(GND_net), .I0(n17_adj_4804), .I1(n86_adj_4805), 
            .CO(n41446));
    SB_LUT4 add_6406_15_lut (.I0(GND_net), .I1(n17773[12]), .I2(n1047_adj_4806), 
            .I3(n40848), .O(n17293[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_19_lut (.I0(GND_net), .I1(n16460[16]), .I2(GND_net), 
            .I3(n41445), .O(n15813[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_18_lut (.I0(GND_net), .I1(n16460[15]), .I2(GND_net), 
            .I3(n41444), .O(n15813[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_18 (.CI(n41444), .I0(n16460[15]), .I1(GND_net), 
            .CO(n41445));
    SB_LUT4 i36787_4_lut (.I0(n37_adj_4753), .I1(n35_adj_4760), .I2(n33_adj_4762), 
            .I3(n52037), .O(n52270));
    defparam i36787_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_6325_17_lut (.I0(GND_net), .I1(n16460[14]), .I2(GND_net), 
            .I3(n41443), .O(n15813[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_17 (.CI(n41443), .I0(n16460[14]), .I1(GND_net), 
            .CO(n41444));
    SB_LUT4 add_6325_16_lut (.I0(GND_net), .I1(n16460[13]), .I2(n1111_adj_4807), 
            .I3(n41442), .O(n15813[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4748), 
            .I3(GND_net), .O(n16_adj_4808));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6325_16 (.CI(n41442), .I0(n16460[13]), .I1(n1111_adj_4807), 
            .CO(n41443));
    SB_LUT4 add_6325_15_lut (.I0(GND_net), .I1(n16460[12]), .I2(n1038_adj_4809), 
            .I3(n41441), .O(n15813[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36666_3_lut (.I0(n6_adj_4732), .I1(n257[10]), .I2(n21_adj_4768), 
            .I3(GND_net), .O(n52149));   // verilog/motorControl.v(38[19:35])
    defparam i36666_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6325_15 (.CI(n41441), .I0(n16460[12]), .I1(n1038_adj_4809), 
            .CO(n41442));
    SB_CARRY add_6270_18 (.CI(n40938), .I0(n15453[15]), .I1(GND_net), 
            .CO(n40939));
    SB_LUT4 add_6325_14_lut (.I0(GND_net), .I1(n16460[11]), .I2(n965_adj_4810), 
            .I3(n41440), .O(n15813[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_14 (.CI(n41440), .I0(n16460[11]), .I1(n965_adj_4810), 
            .CO(n41441));
    SB_LUT4 add_6325_13_lut (.I0(GND_net), .I1(n16460[10]), .I2(n892_adj_4811), 
            .I3(n41439), .O(n15813[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_13 (.CI(n41439), .I0(n16460[10]), .I1(n892_adj_4811), 
            .CO(n41440));
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4812));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6270_17_lut (.I0(GND_net), .I1(n15453[14]), .I2(GND_net), 
            .I3(n40937), .O(n14693[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_12_lut (.I0(GND_net), .I1(n16460[9]), .I2(n819_adj_4813), 
            .I3(n41438), .O(n15813[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_12 (.CI(n41438), .I0(n16460[9]), .I1(n819_adj_4813), 
            .CO(n41439));
    SB_LUT4 add_6325_11_lut (.I0(GND_net), .I1(n16460[8]), .I2(n746_adj_4814), 
            .I3(n41437), .O(n15813[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n40505), .I0(n106[10]), .I1(n155[10]), .CO(n40506));
    SB_CARRY add_6325_11 (.CI(n41437), .I0(n16460[8]), .I1(n746_adj_4814), 
            .CO(n41438));
    SB_LUT4 add_6325_10_lut (.I0(GND_net), .I1(n16460[7]), .I2(n673_adj_4815), 
            .I3(n41436), .O(n15813[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_15 (.CI(n40848), .I0(n17773[12]), .I1(n1047_adj_4806), 
            .CO(n40849));
    SB_LUT4 add_6406_14_lut (.I0(GND_net), .I1(n17773[11]), .I2(n974_adj_4816), 
            .I3(n40847), .O(n17293[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_10 (.CI(n41436), .I0(n16460[7]), .I1(n673_adj_4815), 
            .CO(n41437));
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4817));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4818));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6325_9_lut (.I0(GND_net), .I1(n16460[6]), .I2(n600_adj_4819), 
            .I3(n41435), .O(n15813[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4820));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6325_9 (.CI(n41435), .I0(n16460[6]), .I1(n600_adj_4819), 
            .CO(n41436));
    SB_LUT4 add_6325_8_lut (.I0(GND_net), .I1(n16460[5]), .I2(n527_adj_4821), 
            .I3(n41434), .O(n15813[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6325_8 (.CI(n41434), .I0(n16460[5]), .I1(n527_adj_4821), 
            .CO(n41435));
    SB_LUT4 duty_23__I_851_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(GND_net), .O(n6_adj_4721));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n40504), 
            .O(duty_23__N_3772[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4823));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36667_3_lut (.I0(n52149), .I1(n257[11]), .I2(n23_adj_4758), 
            .I3(GND_net), .O(n52150));   // verilog/motorControl.v(38[19:35])
    defparam i36667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4765), 
            .I3(GND_net), .O(n8_adj_4824));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4808), .I1(n257[22]), .I2(n45_adj_4745), 
            .I3(GND_net), .O(n24_adj_4825));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6325_7_lut (.I0(GND_net), .I1(n16460[4]), .I2(n454_adj_4826), 
            .I3(n41433), .O(n15813[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_7 (.CI(n41433), .I0(n16460[4]), .I1(n454_adj_4826), 
            .CO(n41434));
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36122_4_lut (.I0(n43_adj_4748), .I1(n25_adj_4759), .I2(n23_adj_4758), 
            .I3(n51624), .O(n51604));
    defparam i36122_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4828));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4829));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[23]), 
            .I3(n40672), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_6_lut (.I0(GND_net), .I1(n16460[3]), .I2(n381), .I3(n41432), 
            .O(n15813[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4831));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4832));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4833));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36640_4_lut (.I0(n24_adj_4825), .I1(n8_adj_4824), .I2(n45_adj_4745), 
            .I3(n51602), .O(n52123));   // verilog/motorControl.v(38[19:35])
    defparam i36640_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36311_3_lut (.I0(n52150), .I1(n257[12]), .I2(n25_adj_4759), 
            .I3(GND_net), .O(n51793));   // verilog/motorControl.v(38[19:35])
    defparam i36311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(n257[1]), 
            .I2(duty_23__N_3772[1]), .I3(n257[0]), .O(n4_adj_4835));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4836));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4837));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36664_3_lut (.I0(n4_adj_4835), .I1(n257[13]), .I2(n27_adj_4776), 
            .I3(GND_net), .O(n52147));   // verilog/motorControl.v(38[19:35])
    defparam i36664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36665_3_lut (.I0(n52147), .I1(n257[14]), .I2(n29_adj_4749), 
            .I3(GND_net), .O(n52148));   // verilog/motorControl.v(38[19:35])
    defparam i36665_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6325_6 (.CI(n41432), .I0(n16460[3]), .I1(n381), .CO(n41433));
    SB_LUT4 i36132_4_lut (.I0(n33_adj_4762), .I1(n31_adj_4752), .I2(n29_adj_4749), 
            .I3(n51618), .O(n51614));
    defparam i36132_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36760_4_lut (.I0(n30_adj_4789), .I1(n10_adj_4788), .I2(n35_adj_4760), 
            .I3(n51612), .O(n52243));   // verilog/motorControl.v(38[19:35])
    defparam i36760_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36313_3_lut (.I0(n52148), .I1(n257[15]), .I2(n31_adj_4752), 
            .I3(GND_net), .O(n51795));   // verilog/motorControl.v(38[19:35])
    defparam i36313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6325_5_lut (.I0(GND_net), .I1(n16460[2]), .I2(n308), .I3(n41431), 
            .O(n15813[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_5 (.CI(n41431), .I0(n16460[2]), .I1(n308), .CO(n41432));
    SB_LUT4 add_6325_4_lut (.I0(GND_net), .I1(n16460[1]), .I2(n235), .I3(n41430), 
            .O(n15813[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_4 (.CI(n41430), .I0(n16460[1]), .I1(n235), .CO(n41431));
    SB_LUT4 add_6325_3_lut (.I0(GND_net), .I1(n16460[0]), .I2(n162), .I3(n41429), 
            .O(n15813[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36835_4_lut (.I0(n51795), .I1(n52243), .I2(n35_adj_4760), 
            .I3(n51614), .O(n52318));   // verilog/motorControl.v(38[19:35])
    defparam i36835_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36836_3_lut (.I0(n52318), .I1(n257[18]), .I2(n37_adj_4753), 
            .I3(GND_net), .O(n52319));   // verilog/motorControl.v(38[19:35])
    defparam i36836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36812_3_lut (.I0(n52319), .I1(n257[19]), .I2(n39_adj_4744), 
            .I3(GND_net), .O(n52295));   // verilog/motorControl.v(38[19:35])
    defparam i36812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36124_4_lut (.I0(n43_adj_4748), .I1(n41_adj_4742), .I2(n39_adj_4744), 
            .I3(n52270), .O(n51606));
    defparam i36124_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36782_4_lut (.I0(n51793), .I1(n52123), .I2(n45_adj_4745), 
            .I3(n51604), .O(n52265));   // verilog/motorControl.v(38[19:35])
    defparam i36782_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_6325_3 (.CI(n41429), .I0(n16460[0]), .I1(n162), .CO(n41430));
    SB_LUT4 i36319_3_lut (.I0(n52295), .I1(n257[20]), .I2(n41_adj_4742), 
            .I3(GND_net), .O(n51801));   // verilog/motorControl.v(38[19:35])
    defparam i36319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36784_4_lut (.I0(n51801), .I1(n52265), .I2(n45_adj_4745), 
            .I3(n51606), .O(n52267));   // verilog/motorControl.v(38[19:35])
    defparam i36784_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36785_3_lut (.I0(n52267), .I1(duty_23__N_3772[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256_adj_4839));   // verilog/motorControl.v(38[19:35])
    defparam i36785_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[22]), 
            .I3(n40671), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_2_lut (.I0(GND_net), .I1(n20_adj_4841), .I2(n89), 
            .I3(GND_net), .O(n15813[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_17 (.CI(n40937), .I0(n15453[14]), .I1(GND_net), 
            .CO(n40938));
    SB_CARRY add_6325_2 (.CI(GND_net), .I0(n20_adj_4841), .I1(n89), .CO(n41429));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n40671), .I0(GND_net), .I1(n1_adj_4943[22]), 
            .CO(n40672));
    SB_CARRY add_6406_14 (.CI(n40847), .I0(n17773[11]), .I1(n974_adj_4816), 
            .CO(n40848));
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6406_13_lut (.I0(GND_net), .I1(n17773[10]), .I2(n901_adj_4843), 
            .I3(n40846), .O(n17293[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3772[0]), .I1(n257[0]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6270_16_lut (.I0(GND_net), .I1(n15453[13]), .I2(n1108_adj_4844), 
            .I3(n40936), .O(n14693[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3747[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[21]), 
            .I3(n40670), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4844));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n40670), .I0(GND_net), .I1(n1_adj_4943[21]), 
            .CO(n40671));
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4843));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4841));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_11 (.CI(n40504), .I0(n106[9]), .I1(n155[9]), .CO(n40505));
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n40503), 
            .O(duty_23__N_3772[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i26698_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [19]), .I3(\Ki[1] ), 
            .O(n19933[0]));   // verilog/motorControl.v(34[25:36])
    defparam i26698_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[20]), 
            .I3(n40669), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_18_lut (.I0(GND_net), .I1(n17037[15]), .I2(GND_net), 
            .I3(n41402), .O(n16460[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_17_lut (.I0(GND_net), .I1(n17037[14]), .I2(GND_net), 
            .I3(n41401), .O(n16460[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_17 (.CI(n41401), .I0(n17037[14]), .I1(GND_net), 
            .CO(n41402));
    SB_LUT4 add_6359_16_lut (.I0(GND_net), .I1(n17037[13]), .I2(n1114_adj_4837), 
            .I3(n41400), .O(n16460[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_16 (.CI(n41400), .I0(n17037[13]), .I1(n1114_adj_4837), 
            .CO(n41401));
    SB_LUT4 add_6359_15_lut (.I0(GND_net), .I1(n17037[12]), .I2(n1041_adj_4836), 
            .I3(n41399), .O(n16460[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_15 (.CI(n41399), .I0(n17037[12]), .I1(n1041_adj_4836), 
            .CO(n41400));
    SB_LUT4 add_6359_14_lut (.I0(GND_net), .I1(n17037[11]), .I2(n968_adj_4834), 
            .I3(n41398), .O(n16460[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_14 (.CI(n41398), .I0(n17037[11]), .I1(n968_adj_4834), 
            .CO(n41399));
    SB_LUT4 add_6359_13_lut (.I0(GND_net), .I1(n17037[10]), .I2(n895_adj_4833), 
            .I3(n41397), .O(n16460[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_13 (.CI(n41397), .I0(n17037[10]), .I1(n895_adj_4833), 
            .CO(n41398));
    SB_LUT4 add_6359_12_lut (.I0(GND_net), .I1(n17037[9]), .I2(n822_adj_4832), 
            .I3(n41396), .O(n16460[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_12 (.CI(n41396), .I0(n17037[9]), .I1(n822_adj_4832), 
            .CO(n41397));
    SB_LUT4 add_6359_11_lut (.I0(GND_net), .I1(n17037[8]), .I2(n749_adj_4831), 
            .I3(n41395), .O(n16460[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_11 (.CI(n41395), .I0(n17037[8]), .I1(n749_adj_4831), 
            .CO(n41396));
    SB_LUT4 add_6359_10_lut (.I0(GND_net), .I1(n17037[7]), .I2(n676_adj_4829), 
            .I3(n41394), .O(n16460[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n40669), .I0(GND_net), .I1(n1_adj_4943[20]), 
            .CO(n40670));
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6359_10 (.CI(n41394), .I0(n17037[7]), .I1(n676_adj_4829), 
            .CO(n41395));
    SB_LUT4 add_6359_9_lut (.I0(GND_net), .I1(n17037[6]), .I2(n603_adj_4828), 
            .I3(n41393), .O(n16460[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4943[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[19]), 
            .I3(n40668), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n40668), .I0(GND_net), .I1(n1_adj_4943[19]), 
            .CO(n40669));
    SB_CARRY add_6270_16 (.CI(n40936), .I0(n15453[13]), .I1(n1108_adj_4844), 
            .CO(n40937));
    SB_CARRY add_6406_13 (.CI(n40846), .I0(n17773[10]), .I1(n901_adj_4843), 
            .CO(n40847));
    SB_LUT4 add_6270_15_lut (.I0(GND_net), .I1(n15453[12]), .I2(n1035_adj_4823), 
            .I3(n40935), .O(n14693[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_9 (.CI(n41393), .I0(n17037[6]), .I1(n603_adj_4828), 
            .CO(n41394));
    SB_LUT4 add_6359_8_lut (.I0(GND_net), .I1(n17037[5]), .I2(n530_adj_4822), 
            .I3(n41392), .O(n16460[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_10 (.CI(n40503), .I0(n106[8]), .I1(n155[8]), .CO(n40504));
    SB_CARRY add_6359_8 (.CI(n41392), .I0(n17037[5]), .I1(n530_adj_4822), 
            .CO(n41393));
    SB_LUT4 add_6359_7_lut (.I0(GND_net), .I1(n17037[4]), .I2(n457_adj_4820), 
            .I3(n41391), .O(n16460[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_7 (.CI(n41391), .I0(n17037[4]), .I1(n457_adj_4820), 
            .CO(n41392));
    SB_LUT4 add_6406_12_lut (.I0(GND_net), .I1(n17773[9]), .I2(n828_adj_4818), 
            .I3(n40845), .O(n17293[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_15 (.CI(n40935), .I0(n15453[12]), .I1(n1035_adj_4823), 
            .CO(n40936));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n40502), 
            .O(duty_23__N_3772[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6270_14_lut (.I0(GND_net), .I1(n15453[11]), .I2(n962_adj_4817), 
            .I3(n40934), .O(n14693[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_14 (.CI(n40934), .I0(n15453[11]), .I1(n962_adj_4817), 
            .CO(n40935));
    SB_CARRY add_6406_12 (.CI(n40845), .I0(n17773[9]), .I1(n828_adj_4818), 
            .CO(n40846));
    SB_LUT4 add_6359_6_lut (.I0(GND_net), .I1(n17037[3]), .I2(n384_adj_4812), 
            .I3(n41390), .O(n16460[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_6 (.CI(n41390), .I0(n17037[3]), .I1(n384_adj_4812), 
            .CO(n41391));
    SB_LUT4 add_6359_5_lut (.I0(GND_net), .I1(n17037[2]), .I2(n311_adj_4786), 
            .I3(n41389), .O(n16460[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_5 (.CI(n41389), .I0(n17037[2]), .I1(n311_adj_4786), 
            .CO(n41390));
    SB_LUT4 add_6406_11_lut (.I0(GND_net), .I1(n17773[8]), .I2(n755_adj_4781), 
            .I3(n40844), .O(n17293[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_4_lut (.I0(GND_net), .I1(n17037[1]), .I2(n238_adj_4779), 
            .I3(n41388), .O(n16460[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4826));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6270_13_lut (.I0(GND_net), .I1(n15453[10]), .I2(n889), 
            .I3(n40933), .O(n14693[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_4 (.CI(n41388), .I0(n17037[1]), .I1(n238_adj_4779), 
            .CO(n41389));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[18]), 
            .I3(n40667), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4821));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n40667), .I0(GND_net), .I1(n1_adj_4943[18]), 
            .CO(n40668));
    SB_CARRY add_6406_11 (.CI(n40844), .I0(n17773[8]), .I1(n755_adj_4781), 
            .CO(n40845));
    SB_CARRY add_6270_13 (.CI(n40933), .I0(n15453[10]), .I1(n889), .CO(n40934));
    SB_LUT4 add_6406_10_lut (.I0(GND_net), .I1(n17773[7]), .I2(n682_adj_4770), 
            .I3(n40843), .O(n17293[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_10 (.CI(n40843), .I0(n17773[7]), .I1(n682_adj_4770), 
            .CO(n40844));
    SB_CARRY add_12_9 (.CI(n40502), .I0(n106[7]), .I1(n155[7]), .CO(n40503));
    SB_LUT4 add_6359_3_lut (.I0(GND_net), .I1(n17037[0]), .I2(n165_adj_4769), 
            .I3(n41387), .O(n16460[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6406_9_lut (.I0(GND_net), .I1(n17773[6]), .I2(n609_adj_4764), 
            .I3(n40842), .O(n17293[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_3 (.CI(n41387), .I0(n17037[0]), .I1(n165_adj_4769), 
            .CO(n41388));
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6359_2_lut (.I0(GND_net), .I1(n23_adj_4757), .I2(n92_adj_4756), 
            .I3(GND_net), .O(n16460[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_2 (.CI(GND_net), .I0(n23_adj_4757), .I1(n92_adj_4756), 
            .CO(n41387));
    SB_LUT4 add_6391_17_lut (.I0(GND_net), .I1(n17548[14]), .I2(GND_net), 
            .I3(n41386), .O(n17037[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_16_lut (.I0(GND_net), .I1(n17548[13]), .I2(n1117_adj_4755), 
            .I3(n41385), .O(n17037[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_16 (.CI(n41385), .I0(n17548[13]), .I1(n1117_adj_4755), 
            .CO(n41386));
    SB_LUT4 add_6391_15_lut (.I0(GND_net), .I1(n17548[12]), .I2(n1044_adj_4754), 
            .I3(n41384), .O(n17037[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22014_2_lut (.I0(n1[13]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22014_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[17]), 
            .I3(n40666), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n40501), 
            .O(duty_23__N_3772[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_15 (.CI(n41384), .I0(n17548[12]), .I1(n1044_adj_4754), 
            .CO(n41385));
    SB_LUT4 add_6391_14_lut (.I0(GND_net), .I1(n17548[11]), .I2(n971_adj_4750), 
            .I3(n41383), .O(n17037[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_14 (.CI(n41383), .I0(n17548[11]), .I1(n971_adj_4750), 
            .CO(n41384));
    SB_CARRY unary_minus_16_add_3_19 (.CI(n40666), .I0(GND_net), .I1(n1_adj_4943[17]), 
            .CO(n40667));
    SB_LUT4 add_6391_13_lut (.I0(GND_net), .I1(n17548[10]), .I2(n898_adj_4747), 
            .I3(n41382), .O(n17037[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[16]), 
            .I3(n40665), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_13 (.CI(n41382), .I0(n17548[10]), .I1(n898_adj_4747), 
            .CO(n41383));
    SB_LUT4 add_6270_12_lut (.I0(GND_net), .I1(n15453[9]), .I2(n816), 
            .I3(n40932), .O(n14693[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n40665), .I0(GND_net), .I1(n1_adj_4943[16]), 
            .CO(n40666));
    SB_CARRY add_6406_9 (.CI(n40842), .I0(n17773[6]), .I1(n609_adj_4764), 
            .CO(n40843));
    SB_LUT4 add_6406_8_lut (.I0(GND_net), .I1(n17773[5]), .I2(n536_adj_4743), 
            .I3(n40841), .O(n17293[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_8 (.CI(n40841), .I0(n17773[5]), .I1(n536_adj_4743), 
            .CO(n40842));
    SB_CARRY add_12_8 (.CI(n40501), .I0(n106[6]), .I1(n155[6]), .CO(n40502));
    SB_LUT4 add_6391_12_lut (.I0(GND_net), .I1(n17548[9]), .I2(n825_adj_4741), 
            .I3(n41381), .O(n17037[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n40500), 
            .O(duty_23__N_3772[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_12 (.CI(n41381), .I0(n17548[9]), .I1(n825_adj_4741), 
            .CO(n41382));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[15]), 
            .I3(n40664), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_11_lut (.I0(GND_net), .I1(n17548[8]), .I2(n752_adj_4739), 
            .I3(n41380), .O(n17037[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n40664), .I0(GND_net), .I1(n1_adj_4943[15]), 
            .CO(n40665));
    SB_CARRY add_6391_11 (.CI(n41380), .I0(n17548[8]), .I1(n752_adj_4739), 
            .CO(n41381));
    SB_LUT4 add_6391_10_lut (.I0(GND_net), .I1(n17548[7]), .I2(n679_adj_4738), 
            .I3(n41379), .O(n17037[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_10 (.CI(n41379), .I0(n17548[7]), .I1(n679_adj_4738), 
            .CO(n41380));
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6391_9_lut (.I0(GND_net), .I1(n17548[6]), .I2(n606_adj_4737), 
            .I3(n41378), .O(n17037[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[14]), 
            .I3(n40663), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n40500), .I0(n106[5]), .I1(n155[5]), .CO(n40501));
    SB_LUT4 add_6406_7_lut (.I0(GND_net), .I1(n17773[4]), .I2(n463_adj_4735), 
            .I3(n40840), .O(n17293[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n40663), .I0(GND_net), .I1(n1_adj_4943[14]), 
            .CO(n40664));
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4815));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6391_9 (.CI(n41378), .I0(n17548[6]), .I1(n606_adj_4737), 
            .CO(n41379));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n40499), 
            .O(duty_23__N_3772[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_8_lut (.I0(GND_net), .I1(n17548[5]), .I2(n533_adj_4733), 
            .I3(n41377), .O(n17037[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_8 (.CI(n41377), .I0(n17548[5]), .I1(n533_adj_4733), 
            .CO(n41378));
    SB_LUT4 add_6391_7_lut (.I0(GND_net), .I1(n17548[4]), .I2(n460_adj_4731), 
            .I3(n41376), .O(n17037[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_6 (.CI(n40499), .I0(n106[4]), .I1(n155[4]), .CO(n40500));
    SB_CARRY add_6391_7 (.CI(n41376), .I0(n17548[4]), .I1(n460_adj_4731), 
            .CO(n41377));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[13]), 
            .I3(n40662), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_6_lut (.I0(GND_net), .I1(n17548[3]), .I2(n387_adj_4729), 
            .I3(n41375), .O(n17037[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n40498), 
            .O(duty_23__N_3772[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n40662), .I0(GND_net), .I1(n1_adj_4943[13]), 
            .CO(n40663));
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4814));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6391_6 (.CI(n41375), .I0(n17548[3]), .I1(n387_adj_4729), 
            .CO(n41376));
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4811));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6391_5_lut (.I0(GND_net), .I1(n17548[2]), .I2(n314_adj_4728), 
            .I3(n41374), .O(n17037[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_7 (.CI(n40840), .I0(n17773[4]), .I1(n463_adj_4735), 
            .CO(n40841));
    SB_CARRY add_12_5 (.CI(n40498), .I0(n106[3]), .I1(n155[3]), .CO(n40499));
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4809));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[12]), 
            .I3(n40661), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6406_6_lut (.I0(GND_net), .I1(n17773[3]), .I2(n390_adj_4725), 
            .I3(n40839), .O(n17293[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_5 (.CI(n41374), .I0(n17548[2]), .I1(n314_adj_4728), 
            .CO(n41375));
    SB_CARRY add_6270_12 (.CI(n40932), .I0(n15453[9]), .I1(n816), .CO(n40933));
    SB_CARRY add_6406_6 (.CI(n40839), .I0(n17773[3]), .I1(n390_adj_4725), 
            .CO(n40840));
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n40497), 
            .O(duty_23__N_3772[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_4_lut (.I0(GND_net), .I1(n17548[1]), .I2(n241_adj_4722), 
            .I3(n41373), .O(n17037[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_4 (.CI(n41373), .I0(n17548[1]), .I1(n241_adj_4722), 
            .CO(n41374));
    SB_LUT4 add_6391_3_lut (.I0(GND_net), .I1(n17548[0]), .I2(n168_adj_4711), 
            .I3(n41372), .O(n17037[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_3 (.CI(n41372), .I0(n17548[0]), .I1(n168_adj_4711), 
            .CO(n41373));
    SB_LUT4 add_6391_2_lut (.I0(GND_net), .I1(n26_adj_4710), .I2(n95_adj_4709), 
            .I3(GND_net), .O(n17037[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4807));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4806));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4805));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6391_2 (.CI(GND_net), .I0(n26_adj_4710), .I1(n95_adj_4709), 
            .CO(n41372));
    SB_LUT4 add_6406_5_lut (.I0(GND_net), .I1(n17773[2]), .I2(n317_adj_4707), 
            .I3(n40838), .O(n17293[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_16_lut (.I0(GND_net), .I1(n17997[13]), .I2(n1120), 
            .I3(n41371), .O(n17548[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_4 (.CI(n40497), .I0(n106[2]), .I1(n155[2]), .CO(n40498));
    SB_CARRY unary_minus_16_add_3_14 (.CI(n40661), .I0(GND_net), .I1(n1_adj_4943[12]), 
            .CO(n40662));
    SB_LUT4 add_6270_11_lut (.I0(GND_net), .I1(n15453[8]), .I2(n743), 
            .I3(n40931), .O(n14693[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_15_lut (.I0(GND_net), .I1(n17997[12]), .I2(n1047), 
            .I3(n41370), .O(n17548[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_11 (.CI(n40931), .I0(n15453[8]), .I1(n743), .CO(n40932));
    SB_LUT4 add_6270_10_lut (.I0(GND_net), .I1(n15453[7]), .I2(n670), 
            .I3(n40930), .O(n14693[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_15 (.CI(n41370), .I0(n17997[12]), .I1(n1047), .CO(n41371));
    SB_LUT4 add_6421_14_lut (.I0(GND_net), .I1(n17997[11]), .I2(n974), 
            .I3(n41369), .O(n17548[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_14 (.CI(n41369), .I0(n17997[11]), .I1(n974), .CO(n41370));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[11]), 
            .I3(n40660), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4847));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4547));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n40660), .I0(GND_net), .I1(n1_adj_4943[11]), 
            .CO(n40661));
    SB_CARRY add_6406_5 (.CI(n40838), .I0(n17773[2]), .I1(n317_adj_4707), 
            .CO(n40839));
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4804));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4848));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6270_10 (.CI(n40930), .I0(n15453[7]), .I1(n670), .CO(n40931));
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4803));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6270_9_lut (.I0(GND_net), .I1(n15453[6]), .I2(n597), .I3(n40929), 
            .O(n14693[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6406_4_lut (.I0(GND_net), .I1(n17773[1]), .I2(n244_adj_4696), 
            .I3(n40837), .O(n17293[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[10]), 
            .I3(n40659), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_13_lut (.I0(GND_net), .I1(n17997[10]), .I2(n901), 
            .I3(n41368), .O(n17548[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_13 (.CI(n41368), .I0(n17997[10]), .I1(n901), .CO(n41369));
    SB_LUT4 add_6421_12_lut (.I0(GND_net), .I1(n17997[9]), .I2(n828), 
            .I3(n41367), .O(n17548[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_12 (.CI(n41367), .I0(n17997[9]), .I1(n828), .CO(n41368));
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4802));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6270_9 (.CI(n40929), .I0(n15453[6]), .I1(n597), .CO(n40930));
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4801));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6270_8_lut (.I0(GND_net), .I1(n15453[5]), .I2(n524), .I3(n40928), 
            .O(n14693[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4800));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4799));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4798));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6421_11_lut (.I0(GND_net), .I1(n17997[8]), .I2(n755), 
            .I3(n41366), .O(n17548[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n40659), .I0(GND_net), .I1(n1_adj_4943[10]), 
            .CO(n40660));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[9]), 
            .I3(n40658), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_8 (.CI(n40928), .I0(n15453[5]), .I1(n524), .CO(n40929));
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4796));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n40658), .I0(GND_net), .I1(n1_adj_4943[9]), 
            .CO(n40659));
    SB_CARRY add_6406_4 (.CI(n40837), .I0(n17773[1]), .I1(n244_adj_4696), 
            .CO(n40838));
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n40496), 
            .O(duty_23__N_3772[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6270_7_lut (.I0(GND_net), .I1(n15453[4]), .I2(n451), .I3(n40927), 
            .O(n14693[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_11 (.CI(n41366), .I0(n17997[8]), .I1(n755), .CO(n41367));
    SB_CARRY add_6270_7 (.CI(n40927), .I0(n15453[4]), .I1(n451), .CO(n40928));
    SB_LUT4 add_6421_10_lut (.I0(GND_net), .I1(n17997[7]), .I2(n682), 
            .I3(n41365), .O(n17548[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_10 (.CI(n41365), .I0(n17997[7]), .I1(n682), .CO(n41366));
    SB_LUT4 add_6421_9_lut (.I0(GND_net), .I1(n17997[6]), .I2(n609), .I3(n41364), 
            .O(n17548[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_9 (.CI(n41364), .I0(n17997[6]), .I1(n609), .CO(n41365));
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4795));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35906_2_lut (.I0(n7_adj_4660), .I1(n5_adj_4849), .I2(GND_net), 
            .I3(GND_net), .O(n51388));
    defparam i35906_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4850));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4794));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4793));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26700_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [19]), .I3(\Ki[1] ), 
            .O(n40190));   // verilog/motorControl.v(34[25:36])
    defparam i26700_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_6421_8_lut (.I0(GND_net), .I1(n17997[5]), .I2(n536), .I3(n41363), 
            .O(n17548[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_8 (.CI(n41363), .I0(n17997[5]), .I1(n536), .CO(n41364));
    SB_LUT4 add_6421_7_lut (.I0(GND_net), .I1(n17997[4]), .I2(n463), .I3(n41362), 
            .O(n17548[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_7 (.CI(n41362), .I0(n17997[4]), .I1(n463), .CO(n41363));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[8]), 
            .I3(n40657), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_3 (.CI(n40496), .I0(n106[1]), .I1(n155[1]), .CO(n40497));
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3772[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6270_6_lut (.I0(GND_net), .I1(n15453[3]), .I2(n378), .I3(n40926), 
            .O(n14693[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n40657), .I0(GND_net), .I1(n1_adj_4943[8]), 
            .CO(n40658));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[7]), 
            .I3(n40656), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n40656), .I0(GND_net), .I1(n1_adj_4943[7]), 
            .CO(n40657));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[6]), 
            .I3(n40655), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6421_6_lut (.I0(GND_net), .I1(n17997[3]), .I2(n390), .I3(n41361), 
            .O(n17548[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_6 (.CI(n41361), .I0(n17997[3]), .I1(n390), .CO(n41362));
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4851));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6421_5_lut (.I0(GND_net), .I1(n17997[2]), .I2(n317), .I3(n41360), 
            .O(n17548[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n40496));
    SB_CARRY add_6421_5 (.CI(n41360), .I0(n17997[2]), .I1(n317), .CO(n41361));
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4792));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6421_4_lut (.I0(GND_net), .I1(n17997[1]), .I2(n244), .I3(n41359), 
            .O(n17548[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_4 (.CI(n41359), .I0(n17997[1]), .I1(n244), .CO(n41360));
    SB_LUT4 add_6421_3_lut (.I0(GND_net), .I1(n17997[0]), .I2(n171_adj_4634), 
            .I3(n41358), .O(n17548[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_3 (.CI(n41358), .I0(n17997[0]), .I1(n171_adj_4634), 
            .CO(n41359));
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4852));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4853));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4791));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4790));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6406_3_lut (.I0(GND_net), .I1(n17773[0]), .I2(n171), .I3(n40836), 
            .O(n17293[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_2_lut (.I0(GND_net), .I1(n29_adj_4633), .I2(n98_adj_4632), 
            .I3(GND_net), .O(n17548[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_2 (.CI(GND_net), .I0(n29_adj_4633), .I1(n98_adj_4632), 
            .CO(n41358));
    SB_LUT4 add_6449_15_lut (.I0(GND_net), .I1(n18388[12]), .I2(n1050_adj_4630), 
            .I3(n41357), .O(n17997[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4854));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6449_14_lut (.I0(GND_net), .I1(n18388[11]), .I2(n977_adj_4629), 
            .I3(n41356), .O(n17997[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4787));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4785));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4784));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6449_14 (.CI(n41356), .I0(n18388[11]), .I1(n977_adj_4629), 
            .CO(n41357));
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4783));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6449_13_lut (.I0(GND_net), .I1(n18388[10]), .I2(n904_adj_4622), 
            .I3(n41355), .O(n17997[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4782));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6406_3 (.CI(n40836), .I0(n17773[0]), .I1(n171), .CO(n40837));
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4780));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6449_13 (.CI(n41355), .I0(n18388[10]), .I1(n904_adj_4622), 
            .CO(n41356));
    SB_LUT4 add_6449_12_lut (.I0(GND_net), .I1(n18388[9]), .I2(n831_adj_4619), 
            .I3(n41354), .O(n17997[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_12 (.CI(n41354), .I0(n18388[9]), .I1(n831_adj_4619), 
            .CO(n41355));
    SB_LUT4 add_6449_11_lut (.I0(GND_net), .I1(n18388[8]), .I2(n758_adj_4617), 
            .I3(n41353), .O(n17997[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_11 (.CI(n41353), .I0(n18388[8]), .I1(n758_adj_4617), 
            .CO(n41354));
    SB_LUT4 add_6449_10_lut (.I0(GND_net), .I1(n18388[7]), .I2(n685_adj_4616), 
            .I3(n41352), .O(n17997[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6449_10 (.CI(n41352), .I0(n18388[7]), .I1(n685_adj_4616), 
            .CO(n41353));
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6449_9_lut (.I0(GND_net), .I1(n18388[6]), .I2(n612_adj_4615), 
            .I3(n41351), .O(n17997[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_9 (.CI(n41351), .I0(n18388[6]), .I1(n612_adj_4615), 
            .CO(n41352));
    SB_LUT4 add_6449_8_lut (.I0(GND_net), .I1(n18388[5]), .I2(n539_adj_4614), 
            .I3(n41350), .O(n17997[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_8 (.CI(n41350), .I0(n18388[5]), .I1(n539_adj_4614), 
            .CO(n41351));
    SB_LUT4 add_6449_7_lut (.I0(GND_net), .I1(n18388[4]), .I2(n466_adj_4613), 
            .I3(n41349), .O(n17997[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_7 (.CI(n41349), .I0(n18388[4]), .I1(n466_adj_4613), 
            .CO(n41350));
    SB_LUT4 add_6406_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n17293[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_6 (.CI(n40926), .I0(n15453[3]), .I1(n378), .CO(n40927));
    SB_CARRY unary_minus_16_add_3_8 (.CI(n40655), .I0(GND_net), .I1(n1_adj_4943[6]), 
            .CO(n40656));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[5]), 
            .I3(n40654), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_6_lut (.I0(GND_net), .I1(n18388[3]), .I2(n393_adj_4594), 
            .I3(n41348), .O(n17997[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_6 (.CI(n41348), .I0(n18388[3]), .I1(n393_adj_4594), 
            .CO(n41349));
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4855));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4856));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6449_5_lut (.I0(GND_net), .I1(n18388[2]), .I2(n320_adj_4593), 
            .I3(n41347), .O(n17997[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6270_5_lut (.I0(GND_net), .I1(n15453[2]), .I2(n305), .I3(n40925), 
            .O(n14693[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_5 (.CI(n41347), .I0(n18388[2]), .I1(n320_adj_4593), 
            .CO(n41348));
    SB_LUT4 add_6449_4_lut (.I0(GND_net), .I1(n18388[1]), .I2(n247_adj_4592), 
            .I3(n41346), .O(n17997[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_4 (.CI(n41346), .I0(n18388[1]), .I1(n247_adj_4592), 
            .CO(n41347));
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4857));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6449_3_lut (.I0(GND_net), .I1(n18388[0]), .I2(n174_adj_4591), 
            .I3(n41345), .O(n17997[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4858));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22009_2_lut (.I0(n1[18]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22009_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6449_3 (.CI(n41345), .I0(n18388[0]), .I1(n174_adj_4591), 
            .CO(n41346));
    SB_LUT4 add_6449_2_lut (.I0(GND_net), .I1(n32_adj_4590), .I2(n101_adj_4589), 
            .I3(GND_net), .O(n17997[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_2 (.CI(GND_net), .I0(n32_adj_4590), .I1(n101_adj_4589), 
            .CO(n41345));
    SB_CARRY unary_minus_16_add_3_7 (.CI(n40654), .I0(GND_net), .I1(n1_adj_4943[5]), 
            .CO(n40655));
    SB_CARRY add_6406_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n40836));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[4]), 
            .I3(n40653), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6435_15_lut (.I0(GND_net), .I1(n18193[12]), .I2(n1050), 
            .I3(n40835), .O(n17773[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n40653), .I0(GND_net), .I1(n1_adj_4943[4]), 
            .CO(n40654));
    SB_LUT4 add_6475_14_lut (.I0(GND_net), .I1(n18725[11]), .I2(n980), 
            .I3(n41344), .O(n18388[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6475_13_lut (.I0(GND_net), .I1(n18725[10]), .I2(n907), 
            .I3(n41343), .O(n18388[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_5 (.CI(n40925), .I0(n15453[2]), .I1(n305), .CO(n40926));
    SB_LUT4 add_6435_14_lut (.I0(GND_net), .I1(n18193[11]), .I2(n977), 
            .I3(n40834), .O(n17773[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22013_2_lut (.I0(n1[14]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22013_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6270_4_lut (.I0(GND_net), .I1(n15453[1]), .I2(n232), .I3(n40924), 
            .O(n14693[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_13 (.CI(n41343), .I0(n18725[10]), .I1(n907), .CO(n41344));
    SB_LUT4 add_6475_12_lut (.I0(GND_net), .I1(n18725[9]), .I2(n834), 
            .I3(n41342), .O(n18388[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_12 (.CI(n41342), .I0(n18725[9]), .I1(n834), .CO(n41343));
    SB_LUT4 add_6475_11_lut (.I0(GND_net), .I1(n18725[8]), .I2(n761), 
            .I3(n41341), .O(n18388[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_11 (.CI(n41341), .I0(n18725[8]), .I1(n761), .CO(n41342));
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4859));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6270_4 (.CI(n40924), .I0(n15453[1]), .I1(n232), .CO(n40925));
    SB_CARRY add_6435_14 (.CI(n40834), .I0(n18193[11]), .I1(n977), .CO(n40835));
    SB_LUT4 add_6435_13_lut (.I0(GND_net), .I1(n18193[10]), .I2(n904), 
            .I3(n40833), .O(n17773[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[3]), 
            .I3(n40652), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6475_10_lut (.I0(GND_net), .I1(n18725[7]), .I2(n688), 
            .I3(n41340), .O(n18388[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_10 (.CI(n41340), .I0(n18725[7]), .I1(n688), .CO(n41341));
    SB_LUT4 add_6475_9_lut (.I0(GND_net), .I1(n18725[6]), .I2(n615), .I3(n41339), 
            .O(n18388[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_9 (.CI(n41339), .I0(n18725[6]), .I1(n615), .CO(n41340));
    SB_LUT4 add_6475_8_lut (.I0(GND_net), .I1(n18725[5]), .I2(n542), .I3(n41338), 
            .O(n18388[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_8 (.CI(n41338), .I0(n18725[5]), .I1(n542), .CO(n41339));
    SB_LUT4 add_6475_7_lut (.I0(GND_net), .I1(n18725[4]), .I2(n469), .I3(n41337), 
            .O(n18388[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6270_3_lut (.I0(GND_net), .I1(n15453[0]), .I2(n159), .I3(n40923), 
            .O(n14693[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4777));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6475_7 (.CI(n41337), .I0(n18725[4]), .I1(n469), .CO(n41338));
    SB_CARRY add_6270_3 (.CI(n40923), .I0(n15453[0]), .I1(n159), .CO(n40924));
    SB_LUT4 add_6270_2_lut (.I0(GND_net), .I1(n17_adj_4586), .I2(n86), 
            .I3(GND_net), .O(n14693[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6475_6_lut (.I0(GND_net), .I1(n18725[3]), .I2(n396), .I3(n41336), 
            .O(n18388[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n40652), .I0(GND_net), .I1(n1_adj_4943[3]), 
            .CO(n40653));
    SB_CARRY add_6475_6 (.CI(n41336), .I0(n18725[3]), .I1(n396), .CO(n41337));
    SB_LUT4 add_6475_5_lut (.I0(GND_net), .I1(n18725[2]), .I2(n323), .I3(n41335), 
            .O(n18388[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4860));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6475_5 (.CI(n41335), .I0(n18725[2]), .I1(n323), .CO(n41336));
    SB_LUT4 add_6475_4_lut (.I0(GND_net), .I1(n18725[1]), .I2(n250), .I3(n41334), 
            .O(n18388[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4861));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4862));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6475_4 (.CI(n41334), .I0(n18725[1]), .I1(n250), .CO(n41335));
    SB_LUT4 add_6475_3_lut (.I0(GND_net), .I1(n18725[0]), .I2(n177_adj_4585), 
            .I3(n41333), .O(n18388[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_13 (.CI(n40833), .I0(n18193[10]), .I1(n904), .CO(n40834));
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4863));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22008_2_lut (.I0(n1[19]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22008_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6435_12_lut (.I0(GND_net), .I1(n18193[9]), .I2(n831), 
            .I3(n40832), .O(n17773[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_3 (.CI(n41333), .I0(n18725[0]), .I1(n177_adj_4585), 
            .CO(n41334));
    SB_LUT4 add_6475_2_lut (.I0(GND_net), .I1(n35_adj_4584), .I2(n104_adj_4583), 
            .I3(GND_net), .O(n18388[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_2 (.CI(GND_net), .I0(n35_adj_4584), .I1(n104_adj_4583), 
            .CO(n41333));
    SB_LUT4 add_6499_13_lut (.I0(GND_net), .I1(n19012[10]), .I2(n910_adj_4582), 
            .I3(n41332), .O(n18725[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4864));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22007_2_lut (.I0(n1[20]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22007_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6499_12_lut (.I0(GND_net), .I1(n19012[9]), .I2(n837_adj_4581), 
            .I3(n41331), .O(n18725[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4865));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6499_12 (.CI(n41331), .I0(n19012[9]), .I1(n837_adj_4581), 
            .CO(n41332));
    SB_CARRY add_6435_12 (.CI(n40832), .I0(n18193[9]), .I1(n831), .CO(n40833));
    SB_LUT4 add_6499_11_lut (.I0(GND_net), .I1(n19012[8]), .I2(n764_adj_4580), 
            .I3(n41330), .O(n18725[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4866));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6499_11 (.CI(n41330), .I0(n19012[8]), .I1(n764_adj_4580), 
            .CO(n41331));
    SB_LUT4 add_6435_11_lut (.I0(GND_net), .I1(n18193[8]), .I2(n758), 
            .I3(n40831), .O(n17773[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_11 (.CI(n40831), .I0(n18193[8]), .I1(n758), .CO(n40832));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[2]), 
            .I3(n40651), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_10_lut (.I0(GND_net), .I1(n19012[7]), .I2(n691_adj_4578), 
            .I3(n41329), .O(n18725[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_10 (.CI(n41329), .I0(n19012[7]), .I1(n691_adj_4578), 
            .CO(n41330));
    SB_LUT4 add_6499_9_lut (.I0(GND_net), .I1(n19012[6]), .I2(n618_adj_4577), 
            .I3(n41328), .O(n18725[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n40651), .I0(GND_net), .I1(n1_adj_4943[2]), 
            .CO(n40652));
    SB_CARRY add_6270_2 (.CI(GND_net), .I0(n17_adj_4586), .I1(n86), .CO(n40923));
    SB_CARRY add_6499_9 (.CI(n41328), .I0(n19012[6]), .I1(n618_adj_4577), 
            .CO(n41329));
    SB_LUT4 add_6499_8_lut (.I0(GND_net), .I1(n19012[5]), .I2(n545_adj_4576), 
            .I3(n41327), .O(n18725[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_8 (.CI(n41327), .I0(n19012[5]), .I1(n545_adj_4576), 
            .CO(n41328));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[1]), 
            .I3(n40650), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n40650), .I0(GND_net), .I1(n1_adj_4943[1]), 
            .CO(n40651));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4943[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_7_lut (.I0(GND_net), .I1(n19012[4]), .I2(n472_adj_4573), 
            .I3(n41326), .O(n18725[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_19_lut (.I0(GND_net), .I1(n16137[16]), .I2(GND_net), 
            .I3(n40922), .O(n15453[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4943[0]), 
            .CO(n40650));
    SB_LUT4 add_6435_10_lut (.I0(GND_net), .I1(n18193[7]), .I2(n685), 
            .I3(n40830), .O(n17773[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4942[23]), 
            .I3(n40649), .O(\PID_CONTROLLER.integral_23__N_3723 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_10 (.CI(n40830), .I0(n18193[7]), .I1(n685), .CO(n40831));
    SB_CARRY add_6499_7 (.CI(n41326), .I0(n19012[4]), .I1(n472_adj_4573), 
            .CO(n41327));
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4942[22]), .I3(n40648), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6307_18_lut (.I0(GND_net), .I1(n16137[15]), .I2(GND_net), 
            .I3(n40921), .O(n15453[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6435_9_lut (.I0(GND_net), .I1(n18193[6]), .I2(n612), .I3(n40829), 
            .O(n17773[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_6_lut (.I0(GND_net), .I1(n19012[3]), .I2(n399_adj_4571), 
            .I3(n41325), .O(n18725[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22006_2_lut (.I0(n1[21]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22006_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6435_9 (.CI(n40829), .I0(n18193[6]), .I1(n612), .CO(n40830));
    SB_LUT4 add_6435_8_lut (.I0(GND_net), .I1(n18193[5]), .I2(n539), .I3(n40828), 
            .O(n17773[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4867));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22005_2_lut (.I0(n1[22]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22005_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6307_18 (.CI(n40921), .I0(n16137[15]), .I1(GND_net), 
            .CO(n40922));
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6307_17_lut (.I0(GND_net), .I1(n16137[14]), .I2(GND_net), 
            .I3(n40920), .O(n15453[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_6 (.CI(n41325), .I0(n19012[3]), .I1(n399_adj_4571), 
            .CO(n41326));
    SB_LUT4 add_6499_5_lut (.I0(GND_net), .I1(n19012[2]), .I2(n326_adj_4570), 
            .I3(n41324), .O(n18725[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n40648), .I0(GND_net), .I1(n1_adj_4942[22]), 
            .CO(n40649));
    SB_CARRY add_6499_5 (.CI(n41324), .I0(n19012[2]), .I1(n326_adj_4570), 
            .CO(n41325));
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6499_4_lut (.I0(GND_net), .I1(n19012[1]), .I2(n253_adj_4567), 
            .I3(n41323), .O(n18725[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_4 (.CI(n41323), .I0(n19012[1]), .I1(n253_adj_4567), 
            .CO(n41324));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4942[21]), .I3(n40647), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n40647), .I0(GND_net), .I1(n1_adj_4942[21]), 
            .CO(n40648));
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4869));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22004_2_lut (.I0(n1[23]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22004_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6499_3_lut (.I0(GND_net), .I1(n19012[0]), .I2(n180_adj_4565), 
            .I3(n41322), .O(n18725[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_17 (.CI(n40920), .I0(n16137[14]), .I1(GND_net), 
            .CO(n40921));
    SB_CARRY add_6435_8 (.CI(n40828), .I0(n18193[5]), .I1(n539), .CO(n40829));
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4871));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6499_3 (.CI(n41322), .I0(n19012[0]), .I1(n180_adj_4565), 
            .CO(n41323));
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4872));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4942[20]), .I3(n40646), .O(n41_adj_4665)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6307_16_lut (.I0(GND_net), .I1(n16137[13]), .I2(n1111), 
            .I3(n40919), .O(n15453[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4873));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4874));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6499_2_lut (.I0(GND_net), .I1(n38_adj_4563), .I2(n107_adj_4562), 
            .I3(GND_net), .O(n18725[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4875));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6499_2 (.CI(GND_net), .I0(n38_adj_4563), .I1(n107_adj_4562), 
            .CO(n41322));
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4876));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4878));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4879));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4881));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4882));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n40646), .I0(GND_net), .I1(n1_adj_4942[20]), 
            .CO(n40647));
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4884));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4885));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4886));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4887));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4888));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4890));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6307_16 (.CI(n40919), .I0(n16137[13]), .I1(n1111), .CO(n40920));
    SB_LUT4 add_6307_15_lut (.I0(GND_net), .I1(n16137[12]), .I2(n1038), 
            .I3(n40918), .O(n15453[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4942[19]), .I3(n40645), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6435_7_lut (.I0(GND_net), .I1(n18193[4]), .I2(n466), .I3(n40827), 
            .O(n17773[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_15 (.CI(n40918), .I0(n16137[12]), .I1(n1038), .CO(n40919));
    SB_CARRY add_6435_7 (.CI(n40827), .I0(n18193[4]), .I1(n466), .CO(n40828));
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4891));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4893));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4894));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4896));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n40645), .I0(GND_net), .I1(n1_adj_4942[19]), 
            .CO(n40646));
    SB_LUT4 i22010_2_lut (.I0(n1[17]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22010_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6435_6_lut (.I0(GND_net), .I1(n18193[3]), .I2(n393), .I3(n40826), 
            .O(n17773[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_6 (.CI(n40826), .I0(n18193[3]), .I1(n393), .CO(n40827));
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6307_14_lut (.I0(GND_net), .I1(n16137[11]), .I2(n965), 
            .I3(n40917), .O(n15453[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4899));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4942[18]), .I3(n40644), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6307_14 (.CI(n40917), .I0(n16137[11]), .I1(n965), .CO(n40918));
    SB_LUT4 add_6307_13_lut (.I0(GND_net), .I1(n16137[10]), .I2(n892), 
            .I3(n40916), .O(n15453[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_13 (.CI(n40916), .I0(n16137[10]), .I1(n892), .CO(n40917));
    SB_CARRY unary_minus_5_add_3_20 (.CI(n40644), .I0(GND_net), .I1(n1_adj_4942[18]), 
            .CO(n40645));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4942[17]), .I3(n40643), .O(n35_adj_4611)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6435_5_lut (.I0(GND_net), .I1(n18193[2]), .I2(n320), .I3(n40825), 
            .O(n17773[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_5 (.CI(n40825), .I0(n18193[2]), .I1(n320), .CO(n40826));
    SB_LUT4 add_6307_12_lut (.I0(GND_net), .I1(n16137[9]), .I2(n819), 
            .I3(n40915), .O(n15453[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n40643), .I0(GND_net), .I1(n1_adj_4942[17]), 
            .CO(n40644));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4942[16]), .I3(n40642), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6307_12 (.CI(n40915), .I0(n16137[9]), .I1(n819), .CO(n40916));
    SB_LUT4 add_6307_11_lut (.I0(GND_net), .I1(n16137[8]), .I2(n746), 
            .I3(n40914), .O(n15453[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_11 (.CI(n40914), .I0(n16137[8]), .I1(n746), .CO(n40915));
    SB_LUT4 add_6435_4_lut (.I0(GND_net), .I1(n18193[1]), .I2(n247), .I3(n40824), 
            .O(n17773[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I1(n10300[21]), .I2(GND_net), .I3(n41031), .O(n9793[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6307_10_lut (.I0(GND_net), .I1(n16137[7]), .I2(n673), 
            .I3(n40913), .O(n15453[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_4 (.CI(n40824), .I0(n18193[1]), .I1(n247), .CO(n40825));
    SB_LUT4 add_6435_3_lut (.I0(GND_net), .I1(n18193[0]), .I2(n174), .I3(n40823), 
            .O(n17773[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_3 (.CI(n40823), .I0(n18193[0]), .I1(n174), .CO(n40824));
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22012_2_lut (.I0(n1[15]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22012_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4902));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22011_2_lut (.I0(n1[16]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22011_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4903));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4905));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4906));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n10300[20]), .I2(GND_net), 
            .I3(n41030), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n41030), .I0(n10300[20]), .I1(GND_net), 
            .CO(n41031));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n10300[19]), .I2(GND_net), 
            .I3(n41029), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_10 (.CI(n40913), .I0(n16137[7]), .I1(n673), .CO(n40914));
    SB_LUT4 add_6435_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n17773[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n41029), .I0(n10300[19]), .I1(GND_net), 
            .CO(n41030));
    SB_LUT4 add_6307_9_lut (.I0(GND_net), .I1(n16137[6]), .I2(n600), .I3(n40912), 
            .O(n15453[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n10300[18]), .I2(GND_net), 
            .I3(n41028), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_9 (.CI(n40912), .I0(n16137[6]), .I1(n600), .CO(n40913));
    SB_LUT4 add_6307_8_lut (.I0(GND_net), .I1(n16137[5]), .I2(n527), .I3(n40911), 
            .O(n15453[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_8 (.CI(n40911), .I0(n16137[5]), .I1(n527), .CO(n40912));
    SB_CARRY mult_11_add_1225_21 (.CI(n41028), .I0(n10300[18]), .I1(GND_net), 
            .CO(n41029));
    SB_CARRY unary_minus_5_add_3_18 (.CI(n40642), .I0(GND_net), .I1(n1_adj_4942[16]), 
            .CO(n40643));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4942[15]), .I3(n40641), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n40641), .I0(GND_net), .I1(n1_adj_4942[15]), 
            .CO(n40642));
    SB_LUT4 add_6307_7_lut (.I0(GND_net), .I1(n16137[4]), .I2(n454), .I3(n40910), 
            .O(n15453[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n10300[17]), .I2(GND_net), 
            .I3(n41027), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n40823));
    SB_LUT4 add_6589_8_lut (.I0(GND_net), .I1(n19837[5]), .I2(n560), .I3(n40822), 
            .O(n19740[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4942[14]), .I3(n40640), .O(n29_adj_4606)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4908));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n40640), .I0(GND_net), .I1(n1_adj_4942[14]), 
            .CO(n40641));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4942[13]), .I3(n40639), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n40639), .I0(GND_net), .I1(n1_adj_4942[13]), 
            .CO(n40640));
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4911));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4912));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4913));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4914));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4915));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_11_add_1225_20 (.CI(n41027), .I0(n10300[17]), .I1(GND_net), 
            .CO(n41028));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n10300[16]), .I2(GND_net), 
            .I3(n41026), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4918));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_19 (.CI(n41026), .I0(n10300[16]), .I1(GND_net), 
            .CO(n41027));
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4942[12]), .I3(n40638), .O(n25_adj_4664)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4920));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4921));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4923));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n10300[15]), .I2(GND_net), 
            .I3(n41025), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6589_7_lut (.I0(GND_net), .I1(n19837[4]), .I2(n487_adj_4924), 
            .I3(n40821), .O(n19740[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n41025), .I0(n10300[15]), .I1(GND_net), 
            .CO(n41026));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n10300[14]), .I2(GND_net), 
            .I3(n41024), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6531_11_lut (.I0(GND_net), .I1(n19353[8]), .I2(n770_adj_4925), 
            .I3(n40730), .O(n19133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_7 (.CI(n40910), .I0(n16137[4]), .I1(n454), .CO(n40911));
    SB_LUT4 add_6531_10_lut (.I0(GND_net), .I1(n19353[7]), .I2(n697_adj_4926), 
            .I3(n40729), .O(n19133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4927));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6307_6_lut (.I0(GND_net), .I1(n16137[3]), .I2(n381_adj_4928), 
            .I3(n40909), .O(n15453[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n40638), .I0(GND_net), .I1(n1_adj_4942[12]), 
            .CO(n40639));
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4929));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6589_7 (.CI(n40821), .I0(n19837[4]), .I1(n487_adj_4924), 
            .CO(n40822));
    SB_CARRY add_6307_6 (.CI(n40909), .I0(n16137[3]), .I1(n381_adj_4928), 
            .CO(n40910));
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4930));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4931));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4933));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4942[11]), .I3(n40637), .O(n23_adj_4663)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6589_6_lut (.I0(GND_net), .I1(n19837[3]), .I2(n414_adj_4936), 
            .I3(n40820), .O(n19740[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n40637), .I0(GND_net), .I1(n1_adj_4942[11]), 
            .CO(n40638));
    SB_LUT4 add_6307_5_lut (.I0(GND_net), .I1(n16137[2]), .I2(n308_adj_4937), 
            .I3(n40908), .O(n15453[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4942[10]), .I3(n40636), .O(n21_adj_4662)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6589_6 (.CI(n40820), .I0(n19837[3]), .I1(n414_adj_4936), 
            .CO(n40821));
    SB_CARRY add_6531_10 (.CI(n40729), .I0(n19353[7]), .I1(n697_adj_4926), 
            .CO(n40730));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n40636), .I0(GND_net), .I1(n1_adj_4942[10]), 
            .CO(n40637));
    SB_LUT4 add_6531_9_lut (.I0(GND_net), .I1(n19353[6]), .I2(n624_adj_4933), 
            .I3(n40728), .O(n19133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n41024), .I0(n10300[14]), .I1(GND_net), 
            .CO(n41025));
    SB_CARRY add_6307_5 (.CI(n40908), .I0(n16137[2]), .I1(n308_adj_4937), 
            .CO(n40909));
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4942[9]), .I3(n40635), .O(n19_adj_4550)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n10300[13]), .I2(n1096_adj_4931), 
            .I3(n41023), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_9 (.CI(n40728), .I0(n19353[6]), .I1(n624_adj_4933), 
            .CO(n40729));
    SB_LUT4 add_6589_5_lut (.I0(GND_net), .I1(n19837[2]), .I2(n341_adj_4930), 
            .I3(n40819), .O(n19740[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6589_5 (.CI(n40819), .I0(n19837[2]), .I1(n341_adj_4930), 
            .CO(n40820));
    SB_CARRY mult_11_add_1225_16 (.CI(n41023), .I0(n10300[13]), .I1(n1096_adj_4931), 
            .CO(n41024));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n10300[12]), .I2(n1023_adj_4929), 
            .I3(n41022), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6531_8_lut (.I0(GND_net), .I1(n19353[5]), .I2(n551_adj_4927), 
            .I3(n40727), .O(n19133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_8 (.CI(n40727), .I0(n19353[5]), .I1(n551_adj_4927), 
            .CO(n40728));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n40635), .I0(GND_net), .I1(n1_adj_4942[9]), 
            .CO(n40636));
    SB_LUT4 add_6531_7_lut (.I0(GND_net), .I1(n19353[4]), .I2(n478_adj_4923), 
            .I3(n40726), .O(n19133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4942[8]), .I3(n40634), .O(n17_adj_4556)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6589_4_lut (.I0(GND_net), .I1(n19837[1]), .I2(n268_adj_4921), 
            .I3(n40818), .O(n19740[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n40634), .I0(GND_net), .I1(n1_adj_4942[8]), 
            .CO(n40635));
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4937));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_15 (.CI(n41022), .I0(n10300[12]), .I1(n1023_adj_4929), 
            .CO(n41023));
    SB_CARRY add_6589_4 (.CI(n40818), .I0(n19837[1]), .I1(n268_adj_4921), 
            .CO(n40819));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n10300[11]), .I2(n950_adj_4920), 
            .I3(n41021), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_4_lut (.I0(GND_net), .I1(n16137[1]), .I2(n235_adj_4918), 
            .I3(n40907), .O(n15453[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4936));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4942[7]), .I3(n40633), .O(n15_adj_4608)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n40633), .I0(GND_net), .I1(n1_adj_4942[7]), 
            .CO(n40634));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4942[6]), .I3(n40632), .O(n13_adj_4609)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_11_add_1225_14 (.CI(n41021), .I0(n10300[11]), .I1(n950_adj_4920), 
            .CO(n41022));
    SB_CARRY add_6307_4 (.CI(n40907), .I0(n16137[1]), .I1(n235_adj_4918), 
            .CO(n40908));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n10300[10]), .I2(n877_adj_4915), 
            .I3(n41020), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_3_lut (.I0(GND_net), .I1(n16137[0]), .I2(n162_adj_4914), 
            .I3(n40906), .O(n15453[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6589_3_lut (.I0(GND_net), .I1(n19837[0]), .I2(n195_adj_4913), 
            .I3(n40817), .O(n19740[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_7 (.CI(n40726), .I0(n19353[4]), .I1(n478_adj_4923), 
            .CO(n40727));
    SB_CARRY add_6589_3 (.CI(n40817), .I0(n19837[0]), .I1(n195_adj_4913), 
            .CO(n40818));
    SB_LUT4 add_6589_2_lut (.I0(GND_net), .I1(n53_adj_4912), .I2(n122_adj_4911), 
            .I3(GND_net), .O(n19740[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n41020), .I0(n10300[10]), .I1(n877_adj_4915), 
            .CO(n41021));
    SB_LUT4 add_6531_6_lut (.I0(GND_net), .I1(n19353[3]), .I2(n405_adj_4910), 
            .I3(n40725), .O(n19133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_6 (.CI(n40725), .I0(n19353[3]), .I1(n405_adj_4910), 
            .CO(n40726));
    SB_CARRY unary_minus_5_add_3_8 (.CI(n40632), .I0(GND_net), .I1(n1_adj_4942[6]), 
            .CO(n40633));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4942[5]), .I3(n40631), .O(n11_adj_4938)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6307_3 (.CI(n40906), .I0(n16137[0]), .I1(n162_adj_4914), 
            .CO(n40907));
    SB_LUT4 add_6531_5_lut (.I0(GND_net), .I1(n19353[2]), .I2(n332_adj_4908), 
            .I3(n40724), .O(n19133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_2_lut (.I0(GND_net), .I1(n20_adj_4907), .I2(n89_adj_4906), 
            .I3(GND_net), .O(n15453[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n10300[9]), .I2(n804_adj_4905), 
            .I3(n41019), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6589_2 (.CI(GND_net), .I0(n53_adj_4912), .I1(n122_adj_4911), 
            .CO(n40817));
    SB_CARRY add_6307_2 (.CI(GND_net), .I0(n20_adj_4907), .I1(n89_adj_4906), 
            .CO(n40906));
    SB_CARRY mult_11_add_1225_12 (.CI(n41019), .I0(n10300[9]), .I1(n804_adj_4905), 
            .CO(n41020));
    SB_CARRY unary_minus_5_add_3_7 (.CI(n40631), .I0(GND_net), .I1(n1_adj_4942[5]), 
            .CO(n40632));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n10300[8]), .I2(n731_adj_4904), 
            .I3(n41018), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n41018), .I0(n10300[8]), .I1(n731_adj_4904), 
            .CO(n41019));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n10300[7]), .I2(n658_adj_4903), 
            .I3(n41017), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_5 (.CI(n40724), .I0(n19353[2]), .I1(n332_adj_4908), 
            .CO(n40725));
    SB_LUT4 add_6559_10_lut (.I0(GND_net), .I1(n19613[7]), .I2(n700_adj_4902), 
            .I3(n40905), .O(n19452[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6531_4_lut (.I0(GND_net), .I1(n19353[1]), .I2(n259_adj_4901), 
            .I3(n40723), .O(n19133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n41017), .I0(n10300[7]), .I1(n658_adj_4903), 
            .CO(n41018));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4942[4]), .I3(n40630), .O(n9_adj_4939)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n40630), .I0(GND_net), .I1(n1_adj_4942[4]), 
            .CO(n40631));
    SB_LUT4 add_6559_9_lut (.I0(GND_net), .I1(n19613[6]), .I2(n627_adj_4899), 
            .I3(n40904), .O(n19452[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6462_14_lut (.I0(GND_net), .I1(n18557[11]), .I2(n980_adj_4898), 
            .I3(n40816), .O(n18193[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4942[3]), .I3(n40629), .O(n7_adj_4660)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n10300[6]), .I2(n585_adj_4896), 
            .I3(n41016), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_9 (.CI(n40904), .I0(n19613[6]), .I1(n627_adj_4899), 
            .CO(n40905));
    SB_CARRY mult_11_add_1225_9 (.CI(n41016), .I0(n10300[6]), .I1(n585_adj_4896), 
            .CO(n41017));
    SB_LUT4 add_6462_13_lut (.I0(GND_net), .I1(n18557[10]), .I2(n907_adj_4895), 
            .I3(n40815), .O(n18193[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_13 (.CI(n40815), .I0(n18557[10]), .I1(n907_adj_4895), 
            .CO(n40816));
    SB_LUT4 add_6559_8_lut (.I0(GND_net), .I1(n19613[5]), .I2(n554_adj_4894), 
            .I3(n40903), .O(n19452[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_12_lut (.I0(GND_net), .I1(n19253[9]), .I2(n840_adj_4893), 
            .I3(n41186), .O(n19012[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_11_lut (.I0(GND_net), .I1(n19253[8]), .I2(n767_adj_4892), 
            .I3(n41185), .O(n19012[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n10300[5]), .I2(n512_adj_4891), 
            .I3(n41015), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n41015), .I0(n10300[5]), .I1(n512_adj_4891), 
            .CO(n41016));
    SB_CARRY add_6531_4 (.CI(n40723), .I0(n19353[1]), .I1(n259_adj_4901), 
            .CO(n40724));
    SB_CARRY add_6559_8 (.CI(n40903), .I0(n19613[5]), .I1(n554_adj_4894), 
            .CO(n40904));
    SB_CARRY add_6521_11 (.CI(n41185), .I0(n19253[8]), .I1(n767_adj_4892), 
            .CO(n41186));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n10300[4]), .I2(n439_adj_4890), 
            .I3(n41014), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6531_3_lut (.I0(GND_net), .I1(n19353[0]), .I2(n186_adj_4889), 
            .I3(n40722), .O(n19133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n40629), .I0(GND_net), .I1(n1_adj_4942[3]), 
            .CO(n40630));
    SB_LUT4 add_6521_10_lut (.I0(GND_net), .I1(n19253[7]), .I2(n694_adj_4888), 
            .I3(n41184), .O(n19012[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_10 (.CI(n41184), .I0(n19253[7]), .I1(n694_adj_4888), 
            .CO(n41185));
    SB_LUT4 add_6521_9_lut (.I0(GND_net), .I1(n19253[6]), .I2(n621_adj_4887), 
            .I3(n41183), .O(n19012[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_9 (.CI(n41183), .I0(n19253[6]), .I1(n621_adj_4887), 
            .CO(n41184));
    SB_CARRY add_6531_3 (.CI(n40722), .I0(n19353[0]), .I1(n186_adj_4889), 
            .CO(n40723));
    SB_LUT4 add_6521_8_lut (.I0(GND_net), .I1(n19253[5]), .I2(n548_adj_4886), 
            .I3(n41182), .O(n19012[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6559_7_lut (.I0(GND_net), .I1(n19613[4]), .I2(n481_adj_4885), 
            .I3(n40902), .O(n19452[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_8 (.CI(n41182), .I0(n19253[5]), .I1(n548_adj_4886), 
            .CO(n41183));
    SB_LUT4 add_6462_12_lut (.I0(GND_net), .I1(n18557[9]), .I2(n834_adj_4884), 
            .I3(n40814), .O(n18193[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_7_lut (.I0(GND_net), .I1(n19253[4]), .I2(n475_adj_4883), 
            .I3(n41181), .O(n19012[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_7 (.CI(n41181), .I0(n19253[4]), .I1(n475_adj_4883), 
            .CO(n41182));
    SB_CARRY add_6559_7 (.CI(n40902), .I0(n19613[4]), .I1(n481_adj_4885), 
            .CO(n40903));
    SB_CARRY add_6462_12 (.CI(n40814), .I0(n18557[9]), .I1(n834_adj_4884), 
            .CO(n40815));
    SB_LUT4 add_6531_2_lut (.I0(GND_net), .I1(n44_adj_4882), .I2(n113_adj_4881), 
            .I3(GND_net), .O(n19133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_6_lut (.I0(GND_net), .I1(n19253[3]), .I2(n402_adj_4880), 
            .I3(n41180), .O(n19012[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_2 (.CI(GND_net), .I0(n44_adj_4882), .I1(n113_adj_4881), 
            .CO(n40722));
    SB_CARRY add_6521_6 (.CI(n41180), .I0(n19253[3]), .I1(n402_adj_4880), 
            .CO(n41181));
    SB_LUT4 add_6521_5_lut (.I0(GND_net), .I1(n19253[2]), .I2(n329_adj_4879), 
            .I3(n41179), .O(n19012[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_5 (.CI(n41179), .I0(n19253[2]), .I1(n329_adj_4879), 
            .CO(n41180));
    SB_LUT4 add_6521_4_lut (.I0(GND_net), .I1(n19253[1]), .I2(n256_adj_4878), 
            .I3(n41178), .O(n19012[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4942[2]), .I3(n40628), .O(n5_adj_4849)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6521_4 (.CI(n41178), .I0(n19253[1]), .I1(n256_adj_4878), 
            .CO(n41179));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n40628), .I0(GND_net), .I1(n1_adj_4942[2]), 
            .CO(n40629));
    SB_LUT4 add_6521_3_lut (.I0(GND_net), .I1(n19253[0]), .I2(n183_adj_4876), 
            .I3(n41177), .O(n19012[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6559_6_lut (.I0(GND_net), .I1(n19613[3]), .I2(n408_adj_4875), 
            .I3(n40901), .O(n19452[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_3 (.CI(n41177), .I0(n19253[0]), .I1(n183_adj_4876), 
            .CO(n41178));
    SB_LUT4 add_6521_2_lut (.I0(GND_net), .I1(n41_adj_4874), .I2(n110_adj_4873), 
            .I3(GND_net), .O(n19012[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_6 (.CI(n40901), .I0(n19613[3]), .I1(n408_adj_4875), 
            .CO(n40902));
    SB_CARRY add_6521_2 (.CI(GND_net), .I0(n41_adj_4874), .I1(n110_adj_4873), 
            .CO(n41177));
    SB_LUT4 add_6462_11_lut (.I0(GND_net), .I1(n18557[8]), .I2(n761_adj_4872), 
            .I3(n40813), .O(n18193[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n41014), .I0(n10300[4]), .I1(n439_adj_4890), 
            .CO(n41015));
    SB_LUT4 add_6550_10_lut (.I0(GND_net), .I1(n19533[7]), .I2(n700), 
            .I3(n40721), .O(n19353[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n10300[3]), .I2(n366_adj_4871), 
            .I3(n41013), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4942[1]), .I3(n40627), .O(n3_adj_4604)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_11_add_1225_6 (.CI(n41013), .I0(n10300[3]), .I1(n366_adj_4871), 
            .CO(n41014));
    SB_LUT4 add_904_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n4096[23]), .I3(n40541), .O(\PID_CONTROLLER.integral_23__N_3672 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n10300[2]), .I2(n293_adj_4869), 
            .I3(n41012), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_9_lut (.I0(GND_net), .I1(n19533[6]), .I2(n627), .I3(n40720), 
            .O(n19353[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n40627), .I0(GND_net), .I1(n1_adj_4942[1]), 
            .CO(n40628));
    SB_CARRY mult_11_add_1225_5 (.CI(n41012), .I0(n10300[2]), .I1(n293_adj_4869), 
            .CO(n41013));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4942[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3723 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n4096[22]), .I3(n40540), .O(\PID_CONTROLLER.integral_23__N_3672 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_24 (.CI(n40540), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n4096[22]), .CO(n40541));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n10300[1]), .I2(n220_adj_4867), 
            .I3(n41011), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n4096[21]), .I3(n40539), .O(\PID_CONTROLLER.integral_23__N_3672 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4942[0]), 
            .CO(n40627));
    SB_CARRY mult_11_add_1225_4 (.CI(n41011), .I0(n10300[1]), .I1(n220_adj_4867), 
            .CO(n41012));
    SB_CARRY add_904_23 (.CI(n40539), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n4096[21]), .CO(n40540));
    SB_CARRY add_6462_11 (.CI(n40813), .I0(n18557[8]), .I1(n761_adj_4872), 
            .CO(n40814));
    SB_CARRY add_6550_9 (.CI(n40720), .I0(n19533[6]), .I1(n627), .CO(n40721));
    SB_LUT4 add_6550_8_lut (.I0(GND_net), .I1(n19533[5]), .I2(n554), .I3(n40719), 
            .O(n19353[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_8 (.CI(n40719), .I0(n19533[5]), .I1(n554), .CO(n40720));
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n40626), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n40625), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6462_10_lut (.I0(GND_net), .I1(n18557[7]), .I2(n688_adj_4866), 
            .I3(n40812), .O(n18193[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n10300[0]), .I2(n147_adj_4865), 
            .I3(n41010), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n4096[20]), .I3(n40538), .O(\PID_CONTROLLER.integral_23__N_3672 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6559_5_lut (.I0(GND_net), .I1(n19613[2]), .I2(n335_adj_4864), 
            .I3(n40900), .O(n19452[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_22 (.CI(n40538), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n4096[20]), .CO(n40539));
    SB_CARRY add_6559_5 (.CI(n40900), .I0(n19613[2]), .I1(n335_adj_4864), 
            .CO(n40901));
    SB_LUT4 add_904_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n4096[19]), .I3(n40537), .O(\PID_CONTROLLER.integral_23__N_3672 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_24 (.CI(n40625), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n40626));
    SB_CARRY add_6462_10 (.CI(n40812), .I0(n18557[7]), .I1(n688_adj_4866), 
            .CO(n40813));
    SB_LUT4 add_6559_4_lut (.I0(GND_net), .I1(n19613[1]), .I2(n262_adj_4863), 
            .I3(n40899), .O(n19452[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_4 (.CI(n40899), .I0(n19613[1]), .I1(n262_adj_4863), 
            .CO(n40900));
    SB_CARRY mult_11_add_1225_3 (.CI(n41010), .I0(n10300[0]), .I1(n147_adj_4865), 
            .CO(n41011));
    SB_LUT4 add_6550_7_lut (.I0(GND_net), .I1(n19533[4]), .I2(n481), .I3(n40718), 
            .O(n19353[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4862), .I2(n74_adj_4861), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6559_3_lut (.I0(GND_net), .I1(n19613[0]), .I2(n189_adj_4860), 
            .I3(n40898), .O(n19452[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n40624), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_23 (.CI(n40624), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n40625));
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4862), .I1(n74_adj_4861), 
            .CO(n41010));
    SB_LUT4 add_4572_23_lut (.I0(GND_net), .I1(n11990[20]), .I2(GND_net), 
            .I3(n41009), .O(n10300[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6462_9_lut (.I0(GND_net), .I1(n18557[6]), .I2(n615_adj_4859), 
            .I3(n40811), .O(n18193[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_21 (.CI(n40537), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n4096[19]), .CO(n40538));
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n40623), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_7 (.CI(n40718), .I0(n19533[4]), .I1(n481), .CO(n40719));
    SB_CARRY add_6559_3 (.CI(n40898), .I0(n19613[0]), .I1(n189_adj_4860), 
            .CO(n40899));
    SB_CARRY sub_3_add_2_22 (.CI(n40623), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n40624));
    SB_LUT4 add_4572_22_lut (.I0(GND_net), .I1(n11990[19]), .I2(GND_net), 
            .I3(n41008), .O(n10300[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_22 (.CI(n41008), .I0(n11990[19]), .I1(GND_net), 
            .CO(n41009));
    SB_LUT4 add_904_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4096[18]), .I3(n40536), .O(\PID_CONTROLLER.integral_23__N_3672 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_9 (.CI(n40811), .I0(n18557[6]), .I1(n615_adj_4859), 
            .CO(n40812));
    SB_LUT4 add_6559_2_lut (.I0(GND_net), .I1(n47_adj_4858), .I2(n116_adj_4857), 
            .I3(GND_net), .O(n19452[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35951_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n51433));
    defparam i35951_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 add_4572_21_lut (.I0(GND_net), .I1(n11990[18]), .I2(GND_net), 
            .I3(n41007), .O(n10300[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4572_21 (.CI(n41007), .I0(n11990[18]), .I1(GND_net), 
            .CO(n41008));
    SB_LUT4 add_6550_6_lut (.I0(GND_net), .I1(n19533[3]), .I2(n408), .I3(n40717), 
            .O(n19353[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6462_8_lut (.I0(GND_net), .I1(n18557[5]), .I2(n542_adj_4856), 
            .I3(n40810), .O(n18193[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_8 (.CI(n40810), .I0(n18557[5]), .I1(n542_adj_4856), 
            .CO(n40811));
    SB_CARRY add_6550_6 (.CI(n40717), .I0(n19533[3]), .I1(n408), .CO(n40718));
    SB_LUT4 i35946_3_lut (.I0(n11_adj_4547), .I1(n9_adj_4847), .I2(n51433), 
            .I3(GND_net), .O(n51428));
    defparam i35946_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 add_4572_20_lut (.I0(GND_net), .I1(n11990[17]), .I2(GND_net), 
            .I3(n41006), .O(n10300[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6462_7_lut (.I0(GND_net), .I1(n18557[4]), .I2(n469_adj_4855), 
            .I3(n40809), .O(n18193[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_7 (.CI(n40809), .I0(n18557[4]), .I1(n469_adj_4855), 
            .CO(n40810));
    SB_LUT4 add_6550_5_lut (.I0(GND_net), .I1(n19533[2]), .I2(n335), .I3(n40716), 
            .O(n19353[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n40622), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6462_6_lut (.I0(GND_net), .I1(n18557[3]), .I2(n396_adj_4854), 
            .I3(n40808), .O(n18193[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_6 (.CI(n40808), .I0(n18557[3]), .I1(n396_adj_4854), 
            .CO(n40809));
    SB_CARRY sub_3_add_2_21 (.CI(n40622), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n40623));
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n40621), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_5 (.CI(n40716), .I0(n19533[2]), .I1(n335), .CO(n40717));
    SB_CARRY add_4572_20 (.CI(n41006), .I0(n11990[17]), .I1(GND_net), 
            .CO(n41007));
    SB_CARRY add_904_20 (.CI(n40536), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n4096[18]), .CO(n40537));
    SB_LUT4 add_904_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n4096[17]), .I3(n40535), .O(\PID_CONTROLLER.integral_23__N_3672 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_4_lut (.I0(GND_net), .I1(n19533[1]), .I2(n262_adj_4853), 
            .I3(n40715), .O(n19353[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6462_5_lut (.I0(GND_net), .I1(n18557[2]), .I2(n323_adj_4852), 
            .I3(n40807), .O(n18193[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_4 (.CI(n40715), .I0(n19533[1]), .I1(n262_adj_4853), 
            .CO(n40716));
    SB_CARRY sub_3_add_2_20 (.CI(n40621), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n40622));
    SB_LUT4 add_6550_3_lut (.I0(GND_net), .I1(n19533[0]), .I2(n189_adj_4851), 
            .I3(n40714), .O(n19353[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_2 (.CI(GND_net), .I0(n47_adj_4858), .I1(n116_adj_4857), 
            .CO(n40898));
    SB_CARRY add_6462_5 (.CI(n40807), .I0(n18557[2]), .I1(n323_adj_4852), 
            .CO(n40808));
    SB_LUT4 add_6462_4_lut (.I0(GND_net), .I1(n18557[1]), .I2(n250_adj_4850), 
            .I3(n40806), .O(n18193[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4572_19_lut (.I0(GND_net), .I1(n11990[16]), .I2(GND_net), 
            .I3(n41005), .O(n10300[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4572_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_4 (.CI(n40806), .I0(n18557[1]), .I1(n250_adj_4850), 
            .CO(n40807));
    SB_CARRY add_6550_3 (.CI(n40714), .I0(n19533[0]), .I1(n189_adj_4851), 
            .CO(n40715));
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n40620), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4727));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4720));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4719));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4717));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4716));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4713));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4708));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4705));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4703));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4701));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4695));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4678));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4677));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4676));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4675));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4674));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4672));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4671));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36474_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n53501), 
            .I2(IntegralLimit[7]), .I3(n51428), .O(n51957));
    defparam i36474_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36254_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4848), 
            .I2(IntegralLimit[9]), .I3(n51957), .O(n51736));
    defparam i36254_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4669));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4668));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4659));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4657));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4656));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4655));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4654));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4653));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4652));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4651));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4649));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4648));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4647));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4643));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4642));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4641));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4640));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4639));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4638));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4637));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4636));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4635));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4631));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4628));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4627));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4626));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4625));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4624));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4623));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4621));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36226_4_lut (.I0(n13_adj_4609), .I1(n11_adj_4938), .I2(n9_adj_4939), 
            .I3(n51388), .O(n51708));
    defparam i36226_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_158_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n53484));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_158_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4620));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4599));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4598));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36252_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4848), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4847), .O(n51734));
    defparam i36252_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i26843_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_4940), 
            .I3(n19957[1]), .O(n6_adj_4531));   // verilog/motorControl.v(34[16:22])
    defparam i26843_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n19957[1]), 
            .I3(n4_adj_4940), .O(n19908[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21860_2_lut (.I0(n1[0]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21860_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1519 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n19957[0]), 
            .I3(n40326), .O(n19908[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1519.LUT_INIT = 16'h8778;
    SB_LUT4 i26835_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n40326), 
            .I3(n19957[0]), .O(n4_adj_4940));   // verilog/motorControl.v(34[16:22])
    defparam i26835_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3772[1]), .I1(n257[1]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3747[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3772[2]), .I1(n257[2]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3747[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3747[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3747[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3747[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3747[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3747[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26822_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n19908[0]));   // verilog/motorControl.v(34[16:22])
    defparam i26822_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3747[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3747[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26824_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n40326));   // verilog/motorControl.v(34[16:22])
    defparam i26824_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3747[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3747[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3747[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3747[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3747[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3747[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3747[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3747[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3747[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3747[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3747[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3747[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3747[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3772[23]), .I1(n257[23]), .I2(n256_adj_4839), 
            .I3(GND_net), .O(duty_23__N_3747[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3747[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26781_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n40267), 
            .I3(n20005[0]), .O(n4_adj_4542));   // verilog/motorControl.v(34[16:22])
    defparam i26781_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1520 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n20005[0]), 
            .I3(n40267), .O(n19988[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1520.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1521 (.I0(n62), .I1(n131), .I2(n19988[0]), 
            .I3(n204), .O(n19957[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1521.LUT_INIT = 16'h8778;
    SB_LUT4 i26804_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n19988[0]), 
            .O(n4_adj_4534));   // verilog/motorControl.v(34[16:22])
    defparam i26804_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i26768_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n19988[0]));   // verilog/motorControl.v(34[16:22])
    defparam i26768_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4928));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4926));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26770_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n40267));   // verilog/motorControl.v(34[16:22])
    defparam i26770_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4925));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4924));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26711_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(n40190), .I3(n19973[0]), .O(n4));   // verilog/motorControl.v(34[25:36])
    defparam i26711_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1522 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(n19973[0]), .I3(n40190), .O(n19933[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1522.LUT_INIT = 16'h8778;
    SB_LUT4 i36222_4_lut (.I0(n19_adj_4550), .I1(n17_adj_4556), .I2(n15_adj_4608), 
            .I3(n51708), .O(n51704));
    defparam i36222_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i26673_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n40149), .I3(n19997[0]), .O(n4_adj_4527));   // verilog/motorControl.v(34[25:36])
    defparam i26673_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1523 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n19997[0]), .I3(n40149), .O(n19973[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1523.LUT_INIT = 16'h8778;
    SB_LUT4 i26662_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n40149));   // verilog/motorControl.v(34[25:36])
    defparam i26662_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i26660_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n19973[0]));   // verilog/motorControl.v(34[25:36])
    defparam i26660_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i36694_4_lut (.I0(n25_adj_4664), .I1(n23_adj_4663), .I2(n21_adj_4662), 
            .I3(n51704), .O(n52177));
    defparam i36694_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36250_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n53484), 
            .I2(IntegralLimit[11]), .I3(n51734), .O(n51732));
    defparam i36250_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i36120_2_lut_4_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(duty_23__N_3772[9]), .I3(n257[9]), .O(n51602));
    defparam i36120_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i26750_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n4_adj_4941), .I3(n19933[1]), .O(n6));   // verilog/motorControl.v(34[25:36])
    defparam i26750_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1524 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n19933[1]), .I3(n4_adj_4941), .O(n19873[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1524.LUT_INIT = 16'h8778;
    SB_LUT4 i36208_4_lut (.I0(n27), .I1(n15_adj_4608), .I2(n13_adj_4609), 
            .I3(n11_adj_4938), .O(n51690));
    defparam i36208_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i2_3_lut_4_lut_adj_1525 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n19933[0]), .I3(n40224), .O(n19873[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1525.LUT_INIT = 16'h8778;
    SB_LUT4 i36130_2_lut_4_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(duty_23__N_3772[7]), .I3(n257[7]), .O(n51612));
    defparam i36130_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22026_2_lut (.I0(n1[1]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22026_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22025_2_lut (.I0(n1[2]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22025_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36156_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3772[9]), .O(n51638));
    defparam i36156_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i36166_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3772[7]), .O(n51648));
    defparam i36166_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4603));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i26742_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n40224), .I3(n19933[0]), .O(n4_adj_4941));   // verilog/motorControl.v(34[25:36])
    defparam i26742_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22024_2_lut (.I0(n1[3]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22024_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4561));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36215_4_lut (.I0(n21_adj_4662), .I1(n19_adj_4550), .I2(n17_adj_4556), 
            .I3(n9_adj_4939), .O(n51697));
    defparam i36215_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_4568));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4559));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26791_2_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(\Kp[1] ), 
            .I3(n1[19]), .O(n19957[0]));   // verilog/motorControl.v(34[16:22])
    defparam i26791_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i26729_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n19873[0]));   // verilog/motorControl.v(34[25:36])
    defparam i26729_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i26731_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n40224));   // verilog/motorControl.v(34[25:36])
    defparam i26731_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4942[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000)_U0 
//

module \quadrature_decoder(1,500000)_U0  (\a_new[1] , ENCODER0_B_N_keep, 
            n1653, ENCODER0_A_N_keep, b_prev, direction_N_3907, encoder0_position, 
            GND_net, n29600, n1617, VCC_net) /* synthesis lattice_noprune=1 */ ;
    output \a_new[1] ;
    input ENCODER0_B_N_keep;
    input n1653;
    input ENCODER0_A_N_keep;
    output b_prev;
    output direction_N_3907;
    output [31:0]encoder0_position;
    input GND_net;
    input n29600;
    output n1617;
    input VCC_net;
    
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire a_prev_N_3913, debounce_cnt, n29605, a_prev, n29604;
    wire [31:0]n133;
    
    wire direction_N_3906, direction_N_3910, n41895, n41894, n41893, 
        n41892, n41891, n41890, n41889, n41888, n41887, n41886, 
        n41885, n41884, n41883, n41882, n41881, n41880, n41879, 
        n41878, n41877, n41876, n41875, n41874, n41873, n41872, 
        n41871, n41870, n41869, n41868, n41867, n41866, n41865;
    
    SB_LUT4 i36893_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(57[8:58])
    defparam i36893_4_lut.LUT_INIT = 16'h8421;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1653), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1653), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1653), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1653), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1653), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1653), .D(n29605));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1653), .D(n29604));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2066__i0 (.Q(encoder0_position[0]), .C(n1653), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_DFF direction_57 (.Q(n1617), .C(n1653), .D(n29600));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(\a_new[1] ), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_DFFE position_2066__i1 (.Q(encoder0_position[1]), .C(n1653), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i2 (.Q(encoder0_position[2]), .C(n1653), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i3 (.Q(encoder0_position[3]), .C(n1653), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i4 (.Q(encoder0_position[4]), .C(n1653), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i5 (.Q(encoder0_position[5]), .C(n1653), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i6 (.Q(encoder0_position[6]), .C(n1653), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i7 (.Q(encoder0_position[7]), .C(n1653), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i8 (.Q(encoder0_position[8]), .C(n1653), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i9 (.Q(encoder0_position[9]), .C(n1653), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i10 (.Q(encoder0_position[10]), .C(n1653), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i11 (.Q(encoder0_position[11]), .C(n1653), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i12 (.Q(encoder0_position[12]), .C(n1653), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i13 (.Q(encoder0_position[13]), .C(n1653), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i14 (.Q(encoder0_position[14]), .C(n1653), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i15 (.Q(encoder0_position[15]), .C(n1653), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i16 (.Q(encoder0_position[16]), .C(n1653), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i17 (.Q(encoder0_position[17]), .C(n1653), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i18 (.Q(encoder0_position[18]), .C(n1653), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i19 (.Q(encoder0_position[19]), .C(n1653), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i20 (.Q(encoder0_position[20]), .C(n1653), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i21 (.Q(encoder0_position[21]), .C(n1653), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i22 (.Q(encoder0_position[22]), .C(n1653), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i23 (.Q(encoder0_position[23]), .C(n1653), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i24 (.Q(encoder0_position[24]), .C(n1653), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i25 (.Q(encoder0_position[25]), .C(n1653), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i26 (.Q(encoder0_position[26]), .C(n1653), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i27 (.Q(encoder0_position[27]), .C(n1653), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i28 (.Q(encoder0_position[28]), .C(n1653), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i29 (.Q(encoder0_position[29]), .C(n1653), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i30 (.Q(encoder0_position[30]), .C(n1653), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i31 (.Q(encoder0_position[31]), .C(n1653), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 i16083_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n29605));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16083_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16082_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n29604));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16082_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 position_2066_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[31]), .I3(n41895), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2066_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[30]), .I3(n41894), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_32 (.CI(n41894), .I0(direction_N_3906), 
            .I1(encoder0_position[30]), .CO(n41895));
    SB_LUT4 position_2066_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[29]), .I3(n41893), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_31 (.CI(n41893), .I0(direction_N_3906), 
            .I1(encoder0_position[29]), .CO(n41894));
    SB_LUT4 position_2066_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[28]), .I3(n41892), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_30 (.CI(n41892), .I0(direction_N_3906), 
            .I1(encoder0_position[28]), .CO(n41893));
    SB_LUT4 position_2066_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[27]), .I3(n41891), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_29 (.CI(n41891), .I0(direction_N_3906), 
            .I1(encoder0_position[27]), .CO(n41892));
    SB_LUT4 position_2066_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[26]), .I3(n41890), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_28 (.CI(n41890), .I0(direction_N_3906), 
            .I1(encoder0_position[26]), .CO(n41891));
    SB_LUT4 position_2066_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[25]), .I3(n41889), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_27 (.CI(n41889), .I0(direction_N_3906), 
            .I1(encoder0_position[25]), .CO(n41890));
    SB_LUT4 position_2066_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[24]), .I3(n41888), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_26 (.CI(n41888), .I0(direction_N_3906), 
            .I1(encoder0_position[24]), .CO(n41889));
    SB_LUT4 position_2066_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[23]), .I3(n41887), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_25 (.CI(n41887), .I0(direction_N_3906), 
            .I1(encoder0_position[23]), .CO(n41888));
    SB_LUT4 position_2066_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[22]), .I3(n41886), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_24 (.CI(n41886), .I0(direction_N_3906), 
            .I1(encoder0_position[22]), .CO(n41887));
    SB_LUT4 position_2066_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[21]), .I3(n41885), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_23 (.CI(n41885), .I0(direction_N_3906), 
            .I1(encoder0_position[21]), .CO(n41886));
    SB_LUT4 position_2066_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[20]), .I3(n41884), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_22 (.CI(n41884), .I0(direction_N_3906), 
            .I1(encoder0_position[20]), .CO(n41885));
    SB_LUT4 position_2066_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[19]), .I3(n41883), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_21 (.CI(n41883), .I0(direction_N_3906), 
            .I1(encoder0_position[19]), .CO(n41884));
    SB_LUT4 position_2066_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[18]), .I3(n41882), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_20 (.CI(n41882), .I0(direction_N_3906), 
            .I1(encoder0_position[18]), .CO(n41883));
    SB_LUT4 position_2066_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[17]), .I3(n41881), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_19 (.CI(n41881), .I0(direction_N_3906), 
            .I1(encoder0_position[17]), .CO(n41882));
    SB_LUT4 position_2066_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[16]), .I3(n41880), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_18 (.CI(n41880), .I0(direction_N_3906), 
            .I1(encoder0_position[16]), .CO(n41881));
    SB_LUT4 position_2066_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[15]), .I3(n41879), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_17 (.CI(n41879), .I0(direction_N_3906), 
            .I1(encoder0_position[15]), .CO(n41880));
    SB_LUT4 position_2066_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[14]), .I3(n41878), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_16 (.CI(n41878), .I0(direction_N_3906), 
            .I1(encoder0_position[14]), .CO(n41879));
    SB_LUT4 position_2066_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[13]), .I3(n41877), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_15 (.CI(n41877), .I0(direction_N_3906), 
            .I1(encoder0_position[13]), .CO(n41878));
    SB_LUT4 position_2066_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[12]), .I3(n41876), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_14 (.CI(n41876), .I0(direction_N_3906), 
            .I1(encoder0_position[12]), .CO(n41877));
    SB_LUT4 position_2066_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[11]), .I3(n41875), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_13 (.CI(n41875), .I0(direction_N_3906), 
            .I1(encoder0_position[11]), .CO(n41876));
    SB_LUT4 position_2066_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[10]), .I3(n41874), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_12 (.CI(n41874), .I0(direction_N_3906), 
            .I1(encoder0_position[10]), .CO(n41875));
    SB_LUT4 position_2066_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[9]), .I3(n41873), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_11 (.CI(n41873), .I0(direction_N_3906), 
            .I1(encoder0_position[9]), .CO(n41874));
    SB_LUT4 position_2066_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[8]), .I3(n41872), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_10 (.CI(n41872), .I0(direction_N_3906), 
            .I1(encoder0_position[8]), .CO(n41873));
    SB_LUT4 position_2066_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[7]), .I3(n41871), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_9 (.CI(n41871), .I0(direction_N_3906), 
            .I1(encoder0_position[7]), .CO(n41872));
    SB_LUT4 position_2066_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[6]), .I3(n41870), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_8 (.CI(n41870), .I0(direction_N_3906), 
            .I1(encoder0_position[6]), .CO(n41871));
    SB_LUT4 position_2066_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[5]), .I3(n41869), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_7 (.CI(n41869), .I0(direction_N_3906), 
            .I1(encoder0_position[5]), .CO(n41870));
    SB_LUT4 position_2066_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[4]), .I3(n41868), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_6 (.CI(n41868), .I0(direction_N_3906), 
            .I1(encoder0_position[4]), .CO(n41869));
    SB_LUT4 position_2066_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[3]), .I3(n41867), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_5 (.CI(n41867), .I0(direction_N_3906), 
            .I1(encoder0_position[3]), .CO(n41868));
    SB_LUT4 position_2066_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[2]), .I3(n41866), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_4 (.CI(n41866), .I0(direction_N_3906), 
            .I1(encoder0_position[2]), .CO(n41867));
    SB_LUT4 position_2066_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[1]), .I3(n41865), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_3 (.CI(n41865), .I0(direction_N_3906), 
            .I1(encoder0_position[1]), .CO(n41866));
    SB_LUT4 position_2066_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n41865));
    
endmodule
//
// Verilog Description of module \grp_debouncer(3,1000) 
//

module \grp_debouncer(3,1000)  (reg_B, CLK_c, GND_net, VCC_net, n29608, 
            data_o, n29606, data_i, n48513, n29540);
    output [2:0]reg_B;
    input CLK_c;
    input GND_net;
    input VCC_net;
    input n29608;
    output [2:0]data_o;
    input n29606;
    input [2:0]data_i;
    output n48513;
    input n29540;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [9:0]n45;
    wire [9:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n41818, n41817, n41816, n41815, n41814, n41813, n41812, 
        n41811, n41810, cnt_next_9__N_812, n6, n16, n17;
    
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(CLK_c), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_2060_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[9]), 
            .I3(n41818), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_2060_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[8]), 
            .I3(n41817), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_10 (.CI(n41817), .I0(GND_net), .I1(cnt_reg[8]), 
            .CO(n41818));
    SB_LUT4 cnt_reg_2060_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[7]), 
            .I3(n41816), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_9 (.CI(n41816), .I0(GND_net), .I1(cnt_reg[7]), 
            .CO(n41817));
    SB_LUT4 cnt_reg_2060_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n41815), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_8 (.CI(n41815), .I0(GND_net), .I1(cnt_reg[6]), 
            .CO(n41816));
    SB_LUT4 cnt_reg_2060_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n41814), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_7 (.CI(n41814), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n41815));
    SB_LUT4 cnt_reg_2060_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n41813), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_6 (.CI(n41813), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n41814));
    SB_LUT4 cnt_reg_2060_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n41812), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_5 (.CI(n41812), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n41813));
    SB_LUT4 cnt_reg_2060_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n41811), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_4 (.CI(n41811), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n41812));
    SB_LUT4 cnt_reg_2060_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n41810), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_3 (.CI(n41810), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n41811));
    SB_LUT4 cnt_reg_2060_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n41810));
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(CLK_c), .D(n29608));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i2 (.Q(data_o[2]), .C(CLK_c), .D(n29606));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_2060__i0 (.Q(cnt_reg[0]), .C(CLK_c), .D(n45[0]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i2 (.Q(reg_B[2]), .C(CLK_c), .D(reg_A[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(CLK_c), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(CLK_c), .D(data_i[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(CLK_c), .D(data_i[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i2_4_lut (.I0(reg_B[2]), .I1(reg_B[1]), .I2(reg_A[2]), .I3(reg_A[1]), 
            .O(n6));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut (.I0(reg_B[0]), .I1(n6), .I2(n48513), .I3(reg_A[0]), 
            .O(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i3_4_lut.LUT_INIT = 16'hdfef;
    SB_DFFSR cnt_reg_2060__i1 (.Q(cnt_reg[1]), .C(CLK_c), .D(n45[1]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i2 (.Q(cnt_reg[2]), .C(CLK_c), .D(n45[2]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i3 (.Q(cnt_reg[3]), .C(CLK_c), .D(n45[3]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i4 (.Q(cnt_reg[4]), .C(CLK_c), .D(n45[4]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i5 (.Q(cnt_reg[5]), .C(CLK_c), .D(n45[5]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i6 (.Q(cnt_reg[6]), .C(CLK_c), .D(n45[6]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i7 (.Q(cnt_reg[7]), .C(CLK_c), .D(n45[7]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i8 (.Q(cnt_reg[8]), .C(CLK_c), .D(n45[8]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i9 (.Q(cnt_reg[9]), .C(CLK_c), .D(n45[9]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(CLK_c), .D(n29540));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i2 (.Q(reg_A[2]), .C(CLK_c), .D(data_i[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i6_4_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[7]), 
            .I3(cnt_reg[2]), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut (.I0(cnt_reg[4]), .I1(cnt_reg[9]), .I2(cnt_reg[8]), 
            .I3(cnt_reg[5]), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(cnt_reg[6]), .I2(n16), .I3(cnt_reg[3]), 
            .O(n48513));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    
endmodule
//
// Verilog Description of module coms
//

module coms (CLK_c, n122, GND_net, n63, n3684, n8, n3303, \FRAME_MATCHER.state_31__N_2788[2] , 
            \FRAME_MATCHER.i_31__N_2626 , n4452, n7, \data_out_frame[20] , 
            \data_out_frame[24] , \data_in[1] , \data_in[0] , \data_in[3] , 
            \data_in[2] , n771, n29106, n29671, control_mode, \FRAME_MATCHER.state[0] , 
            n63_adj_10, \data_out_frame[25] , n48070, n29670, n29669, 
            n29668, \data_out_frame[14] , \data_out_frame[15] , \data_out_frame[12] , 
            \data_out_frame[13] , n29667, n25095, n29666, n29665, 
            n29664, PWMLimit, n29663, rx_data_ready, setpoint, n29662, 
            n29661, n29660, n29659, n29658, n29657, n29656, n29655, 
            \data_out_frame[8] , \data_out_frame[9] , \data_out_frame[10] , 
            \data_out_frame[11] , n29654, n29653, n29652, n29651, 
            n29650, n29649, n29648, n29647, n29646, n29645, n29644, 
            n29643, n29642, n53344, n53345, DE_c, LED_c, \data_out_frame[6] , 
            \data_out_frame[7] , \data_out_frame[4] , \data_out_frame[5] , 
            \data_out_frame[23] , rx_data, \data_in_frame[1] , \data_in_frame[2] , 
            \data_in_frame[3] , \data_in_frame[4] , tx_active, \data_in_frame[5] , 
            \data_in_frame[6] , \state[2] , \state[3] , n10, \data_out_frame[19] , 
            \data_out_frame[17] , \data_out_frame[18] , \data_out_frame[16] , 
            \data_in_frame[8] , \data_in_frame[9] , \data_in_frame[11] , 
            \data_in_frame[13] , \data_in_frame[12] , \data_in_frame[10] , 
            n30122, IntegralLimit, n30121, n30120, n30119, n30118, 
            n30117, n30116, n30115, n30114, n30113, n30112, n30111, 
            n30110, n30109, n30108, n30107, n30106, n30105, n30104, 
            n30103, n30102, n30101, n30100, n30099, n30098, n30097, 
            n30096, n30095, n30094, n30093, n30092, n30091, n30090, 
            n30089, n30088, n30087, n30086, n30085, n30084, n30083, 
            n30082, n30081, n30080, n30079, n30078, n30077, n30076, 
            n30075, n30074, n30073, n30072, n30071, n30070, n30069, 
            n30068, \Kp[1] , n30067, \Kp[2] , n30066, \Kp[3] , n30065, 
            \Kp[4] , n30064, \Kp[5] , n30063, \Kp[6] , n30062, \Kp[7] , 
            n30061, \Kp[8] , n30060, \Kp[9] , n30059, \Kp[10] , 
            n30058, \Kp[11] , n30057, \Kp[12] , n30056, \Kp[13] , 
            n30055, \Kp[14] , n30054, \Kp[15] , n30053, \Ki[1] , 
            n30052, \Ki[2] , n30051, \Ki[3] , n30050, \Ki[4] , n30049, 
            \Ki[5] , n30048, \Ki[6] , n30047, \Ki[7] , n30046, \Ki[8] , 
            n30045, \Ki[9] , n30044, \Ki[10] , n30043, \Ki[11] , 
            n30042, \Ki[12] , n30041, \Ki[13] , n30040, \Ki[14] , 
            n30039, \Ki[15] , n30038, n30037, n30036, n30035, n30034, 
            n30033, n30032, n30031, n30030, n30029, n30028, n30027, 
            n30026, n30025, n30024, n30023, n30022, n30021, n30020, 
            n30019, n30018, n30017, n30016, n30015, n30014, n30013, 
            n30012, n30011, n30010, n30009, n30008, n30007, n30006, 
            n30005, n30004, n30003, n30002, n30001, n30000, n29999, 
            n29998, n29997, n29996, n29995, n29994, n29993, n29991, 
            n29990, n29989, n29988, n29987, n29986, n29985, n29984, 
            n29983, n29982, n29981, n29980, n29979, n29978, n29977, 
            n29976, n29975, n29974, n29973, n29972, n29971, n29970, 
            n29969, n29968, n29967, n29966, n29965, n29964, n29963, 
            n29962, n29961, n29960, n29959, n29958, n29957, n29956, 
            n29955, n29954, n29953, n29952, n29951, n29950, n29949, 
            n29948, n29947, n29946, n29945, n29944, n29943, n29942, 
            n29941, n29940, n29939, n29938, n29937, n29936, n29935, 
            n29934, n29933, n29932, n29931, n29930, n29929, n29928, 
            n29927, n29926, n29925, n29924, n29923, n29922, n29921, 
            n29920, n29919, n29918, n29917, n29916, n29915, n29914, 
            n29913, n29912, n29911, n29910, n29909, n29908, n29907, 
            n29906, n29905, n29904, n29903, n29902, n29901, n29900, 
            n29899, n29898, n29897, n29896, n29895, n29894, n29893, 
            n29892, n29891, n29890, n29889, n29888, n29887, n29886, 
            n29885, n29884, n29883, n29882, n29881, n29880, n29879, 
            n29878, n29877, neopxl_color, n29876, n29875, n29874, 
            n29873, n29872, n29871, n29870, n29869, n29868, n29867, 
            n29866, n29865, n29864, n29863, n29862, n29861, n29860, 
            n29859, n29858, n29857, n29856, n29855, n44955, n29570, 
            n29569, n29566, n29565, \Ki[0] , n29564, \Kp[0] , n29542, 
            n29541, n25059, n123, ID, n48426, n45588, n113, n114, 
            \state[0] , n6935, n29165, tx_o, r_SM_Main, \r_SM_Main_2__N_3613[1] , 
            \r_Bit_Index[0] , n45528, n29578, n29579, n53403, VCC_net, 
            n20247, n4, tx_enable, n29175, r_SM_Main_adj_18, r_Rx_Data, 
            RX_N_10, \r_SM_Main_2__N_3542[2] , \r_Bit_Index[0]_adj_14 , 
            n27903, n4_adj_15, n45526, n29587, n29582, n45179, n29561, 
            n29560, n29559, n29558, n29557, n29556, n29555, n45591, 
            n4_adj_16, n4_adj_17, n27898, n35507) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    output n122;
    input GND_net;
    output n63;
    output n3684;
    output n8;
    output n3303;
    output \FRAME_MATCHER.state_31__N_2788[2] ;
    output \FRAME_MATCHER.i_31__N_2626 ;
    output n4452;
    output n7;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[24] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[2] ;
    output n771;
    output n29106;
    input n29671;
    output [7:0]control_mode;
    output \FRAME_MATCHER.state[0] ;
    output n63_adj_10;
    output [7:0]\data_out_frame[25] ;
    output n48070;
    input n29670;
    input n29669;
    input n29668;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[13] ;
    input n29667;
    output n25095;
    input n29666;
    input n29665;
    input n29664;
    output [23:0]PWMLimit;
    input n29663;
    output rx_data_ready;
    output [23:0]setpoint;
    input n29662;
    input n29661;
    input n29660;
    input n29659;
    input n29658;
    input n29657;
    input n29656;
    input n29655;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[11] ;
    input n29654;
    input n29653;
    input n29652;
    input n29651;
    input n29650;
    input n29649;
    input n29648;
    input n29647;
    input n29646;
    input n29645;
    input n29644;
    input n29643;
    input n29642;
    input n53344;
    input n53345;
    output DE_c;
    output LED_c;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_in_frame[4] ;
    output tx_active;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[6] ;
    input \state[2] ;
    input \state[3] ;
    output n10;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[10] ;
    input n30122;
    output [23:0]IntegralLimit;
    input n30121;
    input n30120;
    input n30119;
    input n30118;
    input n30117;
    input n30116;
    input n30115;
    input n30114;
    input n30113;
    input n30112;
    input n30111;
    input n30110;
    input n30109;
    input n30108;
    input n30107;
    input n30106;
    input n30105;
    input n30104;
    input n30103;
    input n30102;
    input n30101;
    input n30100;
    input n30099;
    input n30098;
    input n30097;
    input n30096;
    input n30095;
    input n30094;
    input n30093;
    input n30092;
    input n30091;
    input n30090;
    input n30089;
    input n30088;
    input n30087;
    input n30086;
    input n30085;
    input n30084;
    input n30083;
    input n30082;
    input n30081;
    input n30080;
    input n30079;
    input n30078;
    input n30077;
    input n30076;
    input n30075;
    input n30074;
    input n30073;
    input n30072;
    input n30071;
    input n30070;
    input n30069;
    input n30068;
    output \Kp[1] ;
    input n30067;
    output \Kp[2] ;
    input n30066;
    output \Kp[3] ;
    input n30065;
    output \Kp[4] ;
    input n30064;
    output \Kp[5] ;
    input n30063;
    output \Kp[6] ;
    input n30062;
    output \Kp[7] ;
    input n30061;
    output \Kp[8] ;
    input n30060;
    output \Kp[9] ;
    input n30059;
    output \Kp[10] ;
    input n30058;
    output \Kp[11] ;
    input n30057;
    output \Kp[12] ;
    input n30056;
    output \Kp[13] ;
    input n30055;
    output \Kp[14] ;
    input n30054;
    output \Kp[15] ;
    input n30053;
    output \Ki[1] ;
    input n30052;
    output \Ki[2] ;
    input n30051;
    output \Ki[3] ;
    input n30050;
    output \Ki[4] ;
    input n30049;
    output \Ki[5] ;
    input n30048;
    output \Ki[6] ;
    input n30047;
    output \Ki[7] ;
    input n30046;
    output \Ki[8] ;
    input n30045;
    output \Ki[9] ;
    input n30044;
    output \Ki[10] ;
    input n30043;
    output \Ki[11] ;
    input n30042;
    output \Ki[12] ;
    input n30041;
    output \Ki[13] ;
    input n30040;
    output \Ki[14] ;
    input n30039;
    output \Ki[15] ;
    input n30038;
    input n30037;
    input n30036;
    input n30035;
    input n30034;
    input n30033;
    input n30032;
    input n30031;
    input n30030;
    input n30029;
    input n30028;
    input n30027;
    input n30026;
    input n30025;
    input n30024;
    input n30023;
    input n30022;
    input n30021;
    input n30020;
    input n30019;
    input n30018;
    input n30017;
    input n30016;
    input n30015;
    input n30014;
    input n30013;
    input n30012;
    input n30011;
    input n30010;
    input n30009;
    input n30008;
    input n30007;
    input n30006;
    input n30005;
    input n30004;
    input n30003;
    input n30002;
    input n30001;
    input n30000;
    input n29999;
    input n29998;
    input n29997;
    input n29996;
    input n29995;
    input n29994;
    input n29993;
    input n29991;
    input n29990;
    input n29989;
    input n29988;
    input n29987;
    input n29986;
    input n29985;
    input n29984;
    input n29983;
    input n29982;
    input n29981;
    input n29980;
    input n29979;
    input n29978;
    input n29977;
    input n29976;
    input n29975;
    input n29974;
    input n29973;
    input n29972;
    input n29971;
    input n29970;
    input n29969;
    input n29968;
    input n29967;
    input n29966;
    input n29965;
    input n29964;
    input n29963;
    input n29962;
    input n29961;
    input n29960;
    input n29959;
    input n29958;
    input n29957;
    input n29956;
    input n29955;
    input n29954;
    input n29953;
    input n29952;
    input n29951;
    input n29950;
    input n29949;
    input n29948;
    input n29947;
    input n29946;
    input n29945;
    input n29944;
    input n29943;
    input n29942;
    input n29941;
    input n29940;
    input n29939;
    input n29938;
    input n29937;
    input n29936;
    input n29935;
    input n29934;
    input n29933;
    input n29932;
    input n29931;
    input n29930;
    input n29929;
    input n29928;
    input n29927;
    input n29926;
    input n29925;
    input n29924;
    input n29923;
    input n29922;
    input n29921;
    input n29920;
    input n29919;
    input n29918;
    input n29917;
    input n29916;
    input n29915;
    input n29914;
    input n29913;
    input n29912;
    input n29911;
    input n29910;
    input n29909;
    input n29908;
    input n29907;
    input n29906;
    input n29905;
    input n29904;
    input n29903;
    input n29902;
    input n29901;
    input n29900;
    input n29899;
    input n29898;
    input n29897;
    input n29896;
    input n29895;
    input n29894;
    input n29893;
    input n29892;
    input n29891;
    input n29890;
    input n29889;
    input n29888;
    input n29887;
    input n29886;
    input n29885;
    input n29884;
    input n29883;
    input n29882;
    input n29881;
    input n29880;
    input n29879;
    input n29878;
    input n29877;
    output [23:0]neopxl_color;
    input n29876;
    input n29875;
    input n29874;
    input n29873;
    input n29872;
    input n29871;
    input n29870;
    input n29869;
    input n29868;
    input n29867;
    input n29866;
    input n29865;
    input n29864;
    input n29863;
    input n29862;
    input n29861;
    input n29860;
    input n29859;
    input n29858;
    input n29857;
    input n29856;
    input n29855;
    input n44955;
    input n29570;
    input n29569;
    input n29566;
    input n29565;
    output \Ki[0] ;
    input n29564;
    output \Kp[0] ;
    input n29542;
    input n29541;
    output n25059;
    output n123;
    input [7:0]ID;
    output n48426;
    output n45588;
    output n113;
    output n114;
    input \state[0] ;
    output n6935;
    output n29165;
    output tx_o;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3613[1] ;
    output \r_Bit_Index[0] ;
    output n45528;
    input n29578;
    input n29579;
    input n53403;
    input VCC_net;
    output n20247;
    output n4;
    output tx_enable;
    output n29175;
    output [2:0]r_SM_Main_adj_18;
    output r_Rx_Data;
    input RX_N_10;
    output \r_SM_Main_2__N_3542[2] ;
    output \r_Bit_Index[0]_adj_14 ;
    output n27903;
    output n4_adj_15;
    output n45526;
    input n29587;
    input n29582;
    input n45179;
    input n29561;
    input n29560;
    input n29559;
    input n29558;
    input n29557;
    input n29556;
    input n29555;
    input n45591;
    output n4_adj_16;
    output n4_adj_17;
    output n27898;
    output n35507;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n29678;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    
    wire n29677, n29676, n29675, n29674, n29673;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n63_c, n63_adj_4213, n43235, n42795, n45985, n28342, n46348, 
        n45947, n45854, n46144, n16, n17, n27895, n27792, n16_adj_4215, 
        n17_adj_4216, n27959, n27965, n18, n20, n15, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3, n8_adj_4217, n27770, n29672, n27908, n43868, n5, 
        n123_c, n35344, n126, n39684, n33, n44, n42, n43, n41, 
        n40, n39, n50, n45, n8_adj_4218, n39679, n48572, n5_adj_4219, 
        n27974, n10_c, n2_adj_4221, n40467, n2987, n50168, n15_adj_4222, 
        n40468, n42807, n42887, n28364, n10_adj_4223, n14, n20_adj_4224, 
        n19, n50170, n46231, n43927, n47712, n6, n46207;
    wire [7:0]n8825;
    
    wire n29149;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n39687, n43866, n45862, n47334, n43883, n19_adj_4225, n43923, 
        n46210, n46194, n46190, n2_adj_4226, n40466, n43936, n46335, 
        n50452, n50451;
    wire [31:0]\FRAME_MATCHER.state_31__N_2724 ;
    
    wire n36612, n10_adj_4227;
    wire [0:0]n5426;
    wire [2:0]r_SM_Main_2__N_3616;
    
    wire n5389, \FRAME_MATCHER.rx_data_ready_prev , n6560, n29116, n2_adj_4228, 
        n40465, n50360, n50358, n7_adj_4229, n50354, n50352, n7_adj_4230, 
        n2_adj_4231, n40464, n50345, n50343, n7_adj_4232, n50339, 
        n50337, n7_adj_4233, n50321, n50319, n7_adj_4234, n50327, 
        n50325, n7_adj_4235, n50333, n50331, n7_adj_4236, n50318, 
        n50316, n7_adj_4237, n2_adj_4238, n40463, n50436, n50437, 
        n50368, n50367, n50370, n50371, n50374, n50373, n2_adj_4239, 
        n40462, n2_adj_4240, n40461, n2_adj_4241, n40460, n50442, 
        n50443, n50416, n50415, n50376, n2_adj_4242, n40459, n50377, 
        n50386, n50385, n50379, n50380, n50347, n50346, n39690, 
        n27917, n48518, n29367, n45554, n48025, n50382, n50383, 
        n50311, n50310, n50406, n50407, n50413, n50412, n2_adj_4243, 
        n40458, n161, n6583, n6582, n6581, n6580, n6579, n6578, 
        n6577, n6576, n6575, n6574, n6573, n6572, n6571, n6570, 
        n6569, n6568, n6567, n6566, n6565, n6564, n6563, n6562, 
        n6561, n53266, n51354, n50308, n53152, n52005, n53272, 
        n51357, n50305, n53140, n52007, n50344, n45620;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n29568, n4_c, n29840, n29841, n29842, n29843, n53278, 
        n51360, n29844, n50302, n53134, n52009, n29846, n29847, 
        n10_adj_4244, n50338, n53284, n51363, n50296, n53128, n52011, 
        n10_adj_4245, n53302, n51372, n50287, n53104, n52013, n45097, 
        n45011, n45606, n29832, n7_adj_4246, n8_adj_4247, n29833, 
        n29834, n35325, n35323, n45093, n45013, n45089, n45015, 
        n35321, n44947, n35319, n44925, n7_adj_4248, n8_adj_4249, 
        n45085, n44973, n7_adj_4250, n8_adj_4251, n7_adj_4252, n8_adj_4253, 
        n7_adj_4254, n8_adj_4255, n7_adj_4256, n8_adj_4257, n35317, 
        n36148, n35315, n36146, n7_adj_4258, n8_adj_4259, n45081, 
        n44979, n7_adj_4260, n8_adj_4261, n7_adj_4262, n8_adj_4263, 
        n35313, n36144, n45077, n45017, n35311, n36142, n50326, 
        n45073, n44977, n7_adj_4264, n8_adj_4265, n29835, n45069, 
        n44975, n45065, n45019, n45061, n44965, n35309, n44963, 
        n44957, n44983, n45811, n45667, n43663, n46244, n10_adj_4266, 
        n3_adj_4267, n45726, n45661, n13, n11, n42840, Kp_23__N_1237;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n16_adj_4268, n45638, n45610, n5_adj_4269, n28657, n45923, 
        n46014, n17_adj_4270, n29836, n28259, n28264, n48543, n28544, 
        n28226, n28232, n12, n28368, n4_adj_4271, n28537, n31, 
        n25302, n31_adj_4272, n24851, n10_adj_4273, n36131, n9, 
        n36340, n53296, n51369, n50290, n53116, n52015, n29837, 
        n50317, n29838, n29839, n53308, n51336, n8_adj_4274, n29824, 
        n29825, n29826, n29827, n29828, n29829, n45957, n29243;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n47924, n45843, n47539, n47585, n45841, n47083;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n47535, n48369, n47676, n47312, n48140, n47307, n29830, 
        n29831, n51867, n51366, n53311, n53200;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n53305, n53299, n53293, n53287, n53290, n53281, n53275, 
        n2_adj_4275, n3_adj_4276, n8_adj_4277, n2_adj_4278, n3_adj_4279, 
        n2_adj_4280, n3_adj_4281, n2_adj_4282, n3_adj_4283, n2_adj_4284, 
        n3_adj_4285, n2_adj_4286, n3_adj_4287, n2_adj_4288, n3_adj_4289, 
        n2_adj_4290, n3_adj_4291, n2_adj_4292, n3_adj_4293, n2_adj_4294, 
        n3_adj_4295, n2_adj_4296, n3_adj_4297, n2_adj_4298, n3_adj_4299, 
        n2_adj_4300, n3_adj_4301, n2_adj_4302, n3_adj_4303, n2_adj_4304, 
        n3_adj_4305, n2_adj_4306, n3_adj_4307, n2_adj_4308, n3_adj_4309, 
        n2_adj_4310, n3_adj_4311, n2_adj_4312, n3_adj_4313, n2_adj_4314, 
        n3_adj_4315, n2_adj_4316, n3_adj_4317, n3_adj_4318, n3_adj_4319, 
        n3_adj_4320, n3_adj_4321, n3_adj_4322, n3_adj_4323, n3_adj_4324, 
        n3_adj_4325, n3_adj_4326, n3_adj_4327, n8_adj_4328, n45628, 
        n29679;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n36614, n39678, n4_adj_4329, n6_adj_4330, tx_transmit_N_3513, 
        n29816, n29817, n29818, n29819, n8_adj_4331, n29820, n29821, 
        n29822, n29823, n53269, n53263, n53146, n53257, n53176, 
        n53251, n53218, n53245, n53158, n53239, n53194, n53233, 
        n53188, n53227, n53182, n8_adj_4332, n29808, n29809, n29810, 
        n29811, n29812, n40495, n40494, n40493, n29813, n29814, 
        n29815, n40492, n53221, n27968, n39685, n40491, n35330, 
        n39686, n6_adj_4333, n29800, n29801, n29802, n50332, n29803, 
        n29804, n40490, n29805, n50293, n53122, n29806, n29807, 
        n40489, n28111, n45860, n45848, n6_adj_4334, n46362, n15_adj_4335, 
        n8_adj_4336, n29792, n29793, n45959, n14_adj_4337, n29794, 
        n46141, n45884, n43805, n45979, n46222, n29795, n29796, 
        n43876, n42781, n6_adj_4338, n40488, n40487, n29797, n28526, 
        n45697, n6_adj_4339, n14_adj_4341, n46316, n43593, n43920, 
        n15_adj_4342, n27992, n29798, n46213, n45840, n53164, n53215, 
        n53197, n28418, n45674, n29799, n36193, n29784, n29785, 
        n42913, n29786, n53191, n43437, n42923, n29787, n43850, 
        n29, n46228, n28114, n20_adj_4343, n42875, n28149, n28, 
        n42909, n26, n32, n29788, n53185, n53179, n40486, n6_adj_4344, 
        n29789, n46250, n45930, n28331, n12_adj_4345, n29790, n42822, 
        n46178, n42897, n42958, n27578, n53173, n53161, n29791, 
        n28077, n45916, n6_adj_4346, n45612, n29776, n40485, n6_adj_4347, 
        n29777;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n29778, n43846, n40484, n40483, n29779, n45744, n46082, 
        n47119, n29780, n29781, n28584, n45749, n29782, n29783, 
        n28155, n45859, n29768, n43943, n29769, n45707, n46056, 
        n28193, n1699, n28353, n10_adj_4348, n46300, n46371, n10_adj_4349, 
        n46203, n42820, n26026, n24, n45942, n1513, n1516, n22, 
        n27502, n18_adj_4350, n1510, n26_adj_4351, n1241, n1519, 
        n45664, n28466, n28014, n46216, n10_adj_4352, n45867, n45872, 
        n12_adj_4353, n28006, n46150, n29770, n28074, n45688, n46353, 
        n6_adj_4354, n46263;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n46046, n46024, n46294, n8_adj_4355, n17_adj_4356, n46345, 
        n21, n28022, n4_adj_4357, n20_adj_4358, n45818, n29001, 
        n24_adj_4359, n29771, n28645, n28912, n28129, n42915, n46225, 
        n45896;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n46277, n43591, n46260, n43819, n45950;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n45893, n42581, n28279, n45764, n46166, n46156, n46285, 
        n28_adj_4360, n45890, n32_adj_4361, n28447, n46187, n45779, 
        n30, n29772, n31_adj_4362, n29773, n29774, n46099, n28439, 
        n29_adj_4363, n11_adj_4364, n46116, n16_adj_4365, n46257, 
        n17_adj_4366, n48172, n46288, n45881, n12_adj_4367, n45801, 
        n45997, n8_adj_4368, n28275, n45953, n27538, n46380, n24_adj_4369, 
        n36137, n34, n11_adj_4370, n48381, n45836, n38, n28035, 
        n28456, n28_adj_4371, n29775, n28068, n26_adj_4372, n43839, 
        n46122, n46282, n27, n46304, n46103, n25, n40482, n46159, 
        n45815, Kp_23__N_981, n36, n40481, n22_adj_4373, n37, n46092, 
        n46356, n35, n45684, n43009, n46039, n46254, n45878, n14_adj_4374, 
        n46331, n28689, n10_adj_4375, n28486, n46269, n6_adj_4376, 
        n45736, n46272, Kp_23__N_1195, n7_adj_4377, n46077, n45910, 
        n45741, n45825, n12_adj_4378, n46128, n28902, n46377, n28046, 
        n46365, n12_adj_4379, n45982, n28084, n53155, n45644, n45648, 
        n12_adj_4380, n46089, n46237, n46328, n46374, n6_adj_4381, 
        n46181, n46072, n45851, n46386, n66, n6_adj_4382, n28881, 
        n45716, n74, n45993, n28146, n46383, n72, n46006, n29760, 
        n12_adj_4383, n46086, n26083, n46200, n18_adj_4384, n73, 
        n45899, n46350, n20_adj_4385, n42817, n71, n28676, n70, 
        n46313, n16_adj_4386, n46000, n43916, n68, n29761, n45640, 
        n45936, n1191, n12_adj_4387, n29762, n46111, n46042, n69, 
        n29763, n27527, n46307, n46175, n46368, n67, n46172, n46322, 
        n76, n82, n75, n83, n46009, n28651, n46075, n48418, 
        n6_adj_4388, n24_adj_4389, n17_adj_4390, n22_adj_4391, n26_adj_4392, 
        n40480, n45913, n46197, n29764, n50365, n50364, n29765, 
        n10_adj_4393, Kp_23__N_1217, n53149, n51337, n51338, n53143, 
        n17_adj_4394, n16_adj_4395, n29766, n29767, n29752, n6_adj_4396, 
        n27529, n45972, n10_adj_4397, n29753, n29759, n29758, n29757, 
        n29756, n29755, n29754, n29751, n29750, n29749, n29748, 
        n29747, n29746, n29745, n29744, n29743, n29742, n29741, 
        n29740, n29739, n29738, n29737, n29736, n29735, n29734, 
        n29733, n29732, n29731, n29730, n27975, n8_adj_4398, n29729, 
        n29728, n29727, n29726, n29725, n29724, n2076, n29723, 
        n29722, n29721, n29720, n29719, n29718, n29717, n29716, 
        n29715, n29714, n29713, n29712, n29711, n29710, n29709, 
        n29708, n29707, n29706, n29705, n29704, n29703, n29702, 
        n29701, n29700, n29699, n29698, n29697, n29696, n29695, 
        n29694, n29693, n29692, n29691, n29690, n29689, n29688, 
        n29687;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n29686, n29685, n29684, n29683, n29682, n29681, n29680, 
        n28533, n45704, n40479, n6_adj_4399, n28581, n45738, n45758, 
        n45821, n12_adj_4400, n46125, n46133, n8_adj_4401, n45804, 
        n6_adj_4402, n40478, n45797, n45785, n6_adj_4403, n40477, 
        n6_adj_4404, n45788, n12_adj_4405, n46163, n28800, n46234, 
        n40476, n7_adj_4406, n28771, n8_adj_4407, n45902, n10_adj_4408, 
        n7_adj_4409, n9_adj_4410, n45887, n12_adj_4411, n29014, n28213, 
        n14_adj_4412, n46053, n60, n40475, n58, n45990, n42_adj_4413, 
        n68_adj_4414, n66_adj_4415, n67_adj_4416, n45939, n45710, 
        n65, n24_adj_4417, n46003, n62, n64, n63_adj_4418, n40474, 
        n74_adj_4419, n45773, n45_adj_4420, n69_adj_4421, n22_adj_4422, 
        n28992, n18_adj_4423, n26_adj_4424, n48223, n46291, n45791, 
        Kp_23__N_1020, n46119, n28857, n28_adj_4425, n32_adj_4426, 
        n28120, n46067, n46297, n45794, n30_adj_4427, n29005, n45679, 
        n46027, n29_adj_4428, n31_adj_4429, n40473, n53137, n6_adj_4430, 
        n40472, n49, n2_adj_4432, n40471, n45782, n40470, n45926, 
        n46059, n10_adj_4433, n28299, n8_adj_4434, n4_adj_4435, n45969, 
        n28219, n45971, n46342, Kp_23__N_1183, n10_adj_4436, n40469, 
        n16_adj_4437, Kp_23__N_1214, n9_adj_4438, n46049, n46266, 
        n17_adj_4439, n42805, n45807, n28176, n6_adj_4440, n45719, 
        n46095, n12_adj_4441, n45713, n45652, n6_adj_4442, n46359, 
        n46310, n12_adj_4443, n45845, n28287, n28414, n26983, n45905, 
        n10_adj_4444, n6_adj_4445, n12_adj_4446, n45933, n14_adj_4447, 
        n10_adj_4448, n45722, n28540, n42799, n46136, n10_adj_4449, 
        n45833, n10_adj_4450, Kp_23__N_979, n45956, Kp_23__N_988, 
        n45694, n6_adj_4451, n28937, n6_adj_4452, n28673, n6_adj_4453, 
        n45656, n53131, Kp_23__N_977, n14_adj_4454, n10_adj_4455, 
        n12_adj_4456, n46036, n45729, n45671, n6_adj_4457, n12_adj_4458, 
        n45975, n47441, n34776, n8_adj_4459, n46247, n10_adj_4460, 
        n6_adj_4461, n16_adj_4462, n46219, n8_adj_4463, n8_adj_4464, 
        n47492, n46319, n14_adj_4465, n14_adj_4466, n13_adj_4467, 
        n46338, n13_adj_4468, n14_adj_4469, n42881, n15_adj_4470, 
        n10_adj_4471, n48007, n28140, n8_adj_4472, n6_adj_4473, n47431, 
        n18_adj_4474, n14_adj_4475, n17_adj_4476, n13_adj_4477, n12_adj_4478, 
        n11_adj_4479, n24_adj_4480, n53125, n48304, n46153, n8_adj_4481, 
        n14_adj_4482, n7_adj_4483, n13_adj_4484, n6_adj_4485, n47374, 
        n20_adj_4486, n18_adj_4487, n19_adj_4488, n17_adj_4489, n50031, 
        n28_adj_4490, n21_adj_4491, n29_adj_4492, n12_adj_4493, n10_adj_4494, 
        n11_adj_4495, n9_adj_4496, n10_adj_4497, n45517, n20_adj_4498, 
        n19_adj_4499, n21_adj_4500, n6_adj_4501, n25249, n25262, n34_adj_4502, 
        n45_adj_4503, n27916, n1, n5_adj_4504, n46585, n50049, n45770, 
        n35859, n19_adj_4505, n10_adj_4506, n28108, n22_adj_4507, 
        n4_adj_4508, n28_adj_4509, n53119, n53113, n50051, n30_adj_4510, 
        n23, n31_adj_4511, n6_adj_4512, n53101;
    
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(CLK_c), 
           .D(n29678));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(CLK_c), 
           .D(n29677));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(CLK_c), 
           .D(n29676));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(CLK_c), 
           .D(n29675));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(CLK_c), 
           .D(n29674));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(CLK_c), 
           .D(n29673));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_c), .I2(n63_adj_4213), 
            .I3(GND_net), .O(n122));   // verilog/coms.v(112[11:16])
    defparam i1_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_650_Select_2_i8_3_lut (.I0(n63), .I1(n3684), .I2(n122), 
            .I3(GND_net), .O(n8));
    defparam select_650_Select_2_i8_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i21895_3_lut (.I0(n63), .I1(n3303), .I2(n122), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2788[2] ));   // verilog/coms.v(227[6] 229[9])
    defparam i21895_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 select_650_Select_2_i7_4_lut (.I0(n63), .I1(\FRAME_MATCHER.i_31__N_2626 ), 
            .I2(n4452), .I3(n122), .O(n7));
    defparam select_650_Select_2_i7_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i1_2_lut_4_lut (.I0(n43235), .I1(n42795), .I2(\data_out_frame[20] [5]), 
            .I3(\data_out_frame[24] [7]), .O(n45985));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut (.I0(n28342), .I1(n46348), .I2(n45947), .I3(n45854), 
            .O(n46144));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), .I2(\data_in[3] [2]), 
            .I3(\data_in[0] [5]), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [2]), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_in[1] [6]), .I2(n16), .I3(\data_in[3] [7]), 
            .O(n27895));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_871 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n27792), .O(n16_adj_4215));
    defparam i6_4_lut_adj_871.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_872 (.I0(n27895), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_4216));
    defparam i7_4_lut_adj_872.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_873 (.I0(n17_adj_4216), .I1(\data_in[3] [5]), .I2(n16_adj_4215), 
            .I3(\data_in[3] [3]), .O(n63_adj_4213));
    defparam i9_4_lut_adj_873.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_874 (.I0(\data_in[2] [4]), .I1(n27959), .I2(n27965), 
            .I3(\data_in[2] [2]), .O(n18));
    defparam i7_4_lut_adj_874.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_875 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n27895), .O(n20));
    defparam i9_4_lut_adj_875.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [5]), .I1(\data_in[1] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n15));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n15), .I1(n20), .I2(\data_in[0] [3]), .I3(\data_in[1] [4]), 
            .O(n63_c));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i22062_4_lut (.I0(n8_adj_4217), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27770), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i22062_4_lut.LUT_INIT = 16'h3230;
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(CLK_c), 
           .D(n29672));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n27908), .I2(GND_net), 
            .I3(GND_net), .O(n27770));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut (.I0(n28342), .I1(n46348), .I2(\data_out_frame[20] [4]), 
            .I3(GND_net), .O(n43868));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i22061_4_lut (.I0(n5), .I1(\FRAME_MATCHER.i [31]), .I2(\FRAME_MATCHER.i [2]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i22061_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i3_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n123_c), .I2(n35344), 
            .I3(n126), .O(n29106));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_adj_876 (.I0(\FRAME_MATCHER.state [2]), .I1(n39684), 
            .I2(GND_net), .I3(GND_net), .O(n33));
    defparam i1_2_lut_adj_876.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(CLK_c), .D(n29671));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40), .O(n27908));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22064_4_lut (.I0(n8_adj_4218), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27908), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i22064_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n123_c), .I3(n39679), .O(n48572));
    defparam i2_4_lut.LUT_INIT = 16'hffcd;
    SB_LUT4 i3_4_lut_adj_877 (.I0(n5_adj_4219), .I1(n63_adj_10), .I2(n27974), 
            .I3(n48572), .O(n3684));
    defparam i3_4_lut_adj_877.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 add_43_12_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n40467), .O(n2_adj_4221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_3_lut (.I0(\data_in[2] [7]), .I1(n10_c), .I2(\data_in[3] [4]), 
            .I3(GND_net), .O(n27959));
    defparam i5_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i34795_3_lut (.I0(\data_in[3] [0]), .I1(\data_in[2] [2]), .I2(\data_in[1] [5]), 
            .I3(GND_net), .O(n50168));
    defparam i34795_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6_4_lut_adj_878 (.I0(\data_in[1] [0]), .I1(\data_in[0] [6]), 
            .I2(\data_in[2] [4]), .I3(\data_in[0] [3]), .O(n15_adj_4222));
    defparam i6_4_lut_adj_878.LUT_INIT = 16'hfdff;
    SB_CARRY add_43_12 (.CI(n40467), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n40468));
    SB_LUT4 i1_2_lut_3_lut_adj_879 (.I0(\data_out_frame[25] [1]), .I1(n42807), 
            .I2(n42887), .I3(GND_net), .O(n28364));
    defparam i1_2_lut_3_lut_adj_879.LUT_INIT = 16'h6969;
    SB_LUT4 i8_4_lut (.I0(n15_adj_4222), .I1(\data_in[1] [4]), .I2(n50168), 
            .I3(n27959), .O(n27792));
    defparam i8_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4223));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_880 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14));
    defparam i6_4_lut_adj_880.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_881 (.I0(\data_in[3] [6]), .I1(n14), .I2(n10_adj_4223), 
            .I3(\data_in[2] [1]), .O(n27965));
    defparam i7_4_lut_adj_881.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_882 (.I0(n27965), .I1(\data_in[1] [3]), .I2(n27792), 
            .I3(\data_in[2] [0]), .O(n20_adj_4224));
    defparam i8_4_lut_adj_882.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_883 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19));
    defparam i7_4_lut_adj_883.LUT_INIT = 16'hfeff;
    SB_LUT4 i34797_4_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [5]), .I2(\data_in[0] [5]), 
            .I3(\data_in[3] [2]), .O(n50170));
    defparam i34797_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n50170), .I1(n19), .I2(n20_adj_4224), .I3(GND_net), 
            .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[25] [1]), .I1(n42807), .I2(n46231), 
            .I3(n43927), .O(n47712));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_adj_884 (.I0(n33), .I1(n63), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n771), .O(n48070));
    defparam i2_4_lut_adj_884.LUT_INIT = 16'hfafe;
    SB_LUT4 i1_2_lut_3_lut_adj_885 (.I0(\data_out_frame[20] [3]), .I1(n45947), 
            .I2(n45985), .I3(GND_net), .O(n6));
    defparam i1_2_lut_3_lut_adj_885.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_886 (.I0(\data_out_frame[20] [3]), .I1(n45947), 
            .I2(\data_out_frame[24] [5]), .I3(GND_net), .O(n46207));
    defparam i1_2_lut_3_lut_adj_886.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
            .E(n29149), .D(n8825[1]), .R(n39687));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(CLK_c), 
            .E(n29149), .D(n8825[2]), .R(n39687));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(CLK_c), 
            .E(n29149), .D(n8825[3]), .R(n39687));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(CLK_c), 
            .E(n29149), .D(n8825[4]), .R(n39687));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
            .E(n29149), .D(n8825[5]), .R(n39687));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
            .E(n29149), .D(n8825[6]), .R(n39687));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
            .E(n29149), .D(n8825[7]), .R(n39687));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(CLK_c), .D(n29670));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_887 (.I0(n43866), .I1(\data_out_frame[24] [4]), 
            .I2(n43927), .I3(n45862), .O(n47334));
    defparam i2_3_lut_4_lut_adj_887.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut (.I0(n43866), .I1(\data_out_frame[24] [4]), .I2(n43883), 
            .I3(GND_net), .O(n19_adj_4225));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_888 (.I0(n43923), .I1(n46210), .I2(n46194), 
            .I3(n46190), .O(n43883));
    defparam i2_3_lut_4_lut_adj_888.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_11_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n40466), .O(n2_adj_4226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_889 (.I0(n43923), .I1(n46210), .I2(n43936), 
            .I3(n46335), .O(n43866));
    defparam i2_3_lut_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(CLK_c), .D(n29669));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(CLK_c), .D(n29668));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i34970_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50452));
    defparam i34970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34969_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50451));
    defparam i34969_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(CLK_c), .D(n29667));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_890 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state_31__N_2724 [3]), 
            .I2(n36612), .I3(\FRAME_MATCHER.state [3]), .O(n10_adj_4227));
    defparam i4_4_lut_adj_890.LUT_INIT = 16'h0008;
    SB_LUT4 i5_3_lut_adj_891 (.I0(\FRAME_MATCHER.state[0] ), .I1(n10_adj_4227), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n25095));
    defparam i5_3_lut_adj_891.LUT_INIT = 16'h0404;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(CLK_c), .D(n29666));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(CLK_c), .D(n29665));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(CLK_c), .D(n29664));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(CLK_c), .D(n29663));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_11 (.CI(n40466), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n40467));
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3616[0]), .C(CLK_c), .D(n5426[0]), 
            .R(n5389));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(CLK_c), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(CLK_c), .E(n29116), .D(n6560));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
            .E(n29149), .D(n8825[0]), .R(n39687));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_10_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n40465), .O(n2_adj_4228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(CLK_c), .D(n29662));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(CLK_c), .D(n29661));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(CLK_c), .D(n29660));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_10 (.CI(n40465), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n40466));
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(CLK_c), .D(n29659));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(CLK_c), .D(n29658));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50360), .I3(n50358), .O(n7_adj_4229));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(CLK_c), .D(n29657));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(CLK_c), .D(n29656));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50354), .I3(n50352), .O(n7_adj_4230));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 add_43_9_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n40464), .O(n2_adj_4231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50345), .I3(n50343), .O(n7_adj_4232));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50339), .I3(n50337), .O(n7_adj_4233));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50321), .I3(n50319), .O(n7_adj_4234));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50327), .I3(n50325), .O(n7_adj_4235));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(CLK_c), .D(n29655));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_9 (.CI(n40464), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n40465));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50333), .I3(n50331), .O(n7_adj_4236));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50318), .I3(n50316), .O(n7_adj_4237));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 add_43_8_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n40463), .O(n2_adj_4238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i34954_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50436));
    defparam i34954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34955_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50437));
    defparam i34955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34886_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50368));
    defparam i34886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34885_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50367));
    defparam i34885_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(CLK_c), .D(n29654));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i34888_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50370));
    defparam i34888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34889_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50371));
    defparam i34889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34892_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50374));
    defparam i34892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34891_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50373));
    defparam i34891_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_8 (.CI(n40463), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n40464));
    SB_LUT4 add_43_7_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n40462), .O(n2_adj_4239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_7 (.CI(n40462), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n40463));
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(CLK_c), .D(n29653));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(CLK_c), .D(n29652));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(CLK_c), .D(n29651));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(CLK_c), .D(n29650));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(CLK_c), .D(n29649));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(CLK_c), .D(n29648));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(CLK_c), .D(n29647));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(CLK_c), .D(n29646));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(CLK_c), .D(n29645));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(CLK_c), .D(n29644));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(CLK_c), .D(n29643));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_6_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n40461), .O(n2_adj_4240)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(CLK_c), .D(n29642));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_6 (.CI(n40461), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n40462));
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(CLK_c), 
           .D(n53344));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(CLK_c), 
           .D(n53345));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_5_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n40460), .O(n2_adj_4241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_5 (.CI(n40460), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n40461));
    SB_LUT4 i34960_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50442));
    defparam i34960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34961_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50443));
    defparam i34961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34934_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50416));
    defparam i34934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34933_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50415));
    defparam i34933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34894_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50376));
    defparam i34894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n40459), .O(n2_adj_4242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i34895_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50377));
    defparam i34895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34904_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50386));
    defparam i34904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34903_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50385));
    defparam i34903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34897_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50379));
    defparam i34897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34898_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50380));
    defparam i34898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34865_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50347));
    defparam i34865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34864_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50346));
    defparam i34864_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_4 (.CI(n40459), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n40460));
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(CLK_c), .E(n27917), .D(n39690), 
            .R(n48518));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR LED_3874 (.Q(LED_c), .C(CLK_c), .E(n45554), .D(n29367), 
            .R(n48025));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i34900_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50382));
    defparam i34900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34901_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50383));
    defparam i34901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34829_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50311));
    defparam i34829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34828_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50310));
    defparam i34828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34924_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50406));
    defparam i34924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34925_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50407));
    defparam i34925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34931_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50413));
    defparam i34931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34930_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50412));
    defparam i34930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34878_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n50360));
    defparam i34878_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i34876_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50358));
    defparam i34876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_3_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n40458), .O(n2_adj_4243)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_3 (.CI(n40458), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n40459));
    SB_LUT4 add_43_2_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(CLK_c), .E(n29116), .D(n6583));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(CLK_c), .E(n29116), .D(n6582));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(CLK_c), .E(n29116), .D(n6581));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(CLK_c), .E(n29116), .D(n6580));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(CLK_c), .E(n29116), .D(n6579));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(CLK_c), .E(n29116), .D(n6578));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(CLK_c), .E(n29116), .D(n6577));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(CLK_c), .E(n29116), .D(n6576));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(CLK_c), .E(n29116), .D(n6575));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(CLK_c), .E(n29116), .D(n6574));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(CLK_c), .E(n29116), .D(n6573));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(CLK_c), .E(n29116), .D(n6572));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(CLK_c), .E(n29116), .D(n6571));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(CLK_c), .E(n29116), .D(n6570));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(CLK_c), .E(n29116), .D(n6569));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(CLK_c), .E(n29116), .D(n6568));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(CLK_c), .E(n29116), .D(n6567));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(CLK_c), .E(n29116), .D(n6566));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(CLK_c), .E(n29116), .D(n6565));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(CLK_c), .E(n29116), .D(n6564));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(CLK_c), .E(n29116), .D(n6563));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(CLK_c), .E(n29116), .D(n6562));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(CLK_c), .E(n29116), .D(n6561));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n40458));
    SB_LUT4 i36056_2_lut (.I0(n53266), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51354));
    defparam i36056_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34826_4_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n50308));
    defparam i34826_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i36522_3_lut (.I0(n53152), .I1(n50308), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n52005));
    defparam i36522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34872_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n50354));
    defparam i34872_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i34870_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50352));
    defparam i34870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36072_2_lut (.I0(n53272), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51357));
    defparam i36072_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34823_4_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n50305));
    defparam i34823_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i36524_3_lut (.I0(n53140), .I1(n50305), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n52007));
    defparam i36524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34862_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50344));
    defparam i34862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16046_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45620), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n29568));
    defparam i16046_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i36887_3_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(n39690), 
            .I2(n4_c), .I3(n36612), .O(n5389));   // verilog/coms.v(127[12] 300[6])
    defparam i36887_3_lut_4_lut.LUT_INIT = 16'hff0b;
    SB_LUT4 i34863_4_lut (.I0(n50344), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n50345));
    defparam i34863_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i34861_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50343));
    defparam i34861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16318_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45620), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n29840));
    defparam i16318_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16319_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45620), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n29841));
    defparam i16319_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16320_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45620), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n29842));
    defparam i16320_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16321_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45620), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n29843));
    defparam i16321_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i36068_2_lut (.I0(n53278), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51360));
    defparam i36068_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16322_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45620), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n29844));
    defparam i16322_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34820_4_lut (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[23] [5]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n50302));
    defparam i34820_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i36526_3_lut (.I0(n53134), .I1(n50302), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n52009));
    defparam i36526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16324_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45620), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n29846));
    defparam i16324_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16325_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45620), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n29847));
    defparam i16325_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_290_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4244));   // verilog/coms.v(154[7:23])
    defparam equal_290_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i34856_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50338));
    defparam i34856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34857_4_lut (.I0(n50338), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n50339));
    defparam i34857_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i34855_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50337));
    defparam i34855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36065_2_lut (.I0(n53284), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51363));
    defparam i36065_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34814_4_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n50296));
    defparam i34814_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i36528_3_lut (.I0(n53128), .I1(n50296), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n52011));
    defparam i36528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_298_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4245));   // verilog/coms.v(154[7:23])
    defparam equal_298_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i34839_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n50321));
    defparam i34839_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i34837_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50319));
    defparam i34837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36054_2_lut (.I0(n53302), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51372));
    defparam i36054_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34805_4_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n50287));
    defparam i34805_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i36530_3_lut (.I0(n53104), .I1(n50287), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n52013));
    defparam i36530_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(CLK_c), 
            .D(n45097), .S(n45011));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16310_3_lut_4_lut (.I0(n10_adj_4245), .I1(n45606), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29832));
    defparam i16310_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(CLK_c), 
            .D(n7_adj_4246), .S(n8_adj_4247));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16311_3_lut_4_lut (.I0(n10_adj_4245), .I1(n45606), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n29833));
    defparam i16311_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16312_3_lut_4_lut (.I0(n10_adj_4245), .I1(n45606), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29834));
    defparam i16312_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(CLK_c), 
            .D(n35325), .S(n35323));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(CLK_c), 
            .D(n45093), .S(n45013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(CLK_c), 
            .D(n45089), .S(n45015));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(CLK_c), 
            .D(n35321), .S(n44947));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(CLK_c), 
            .D(n35319), .S(n44925));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(CLK_c), 
            .D(n7_adj_4248), .S(n8_adj_4249));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(CLK_c), 
            .D(n45085), .S(n44973));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(CLK_c), 
            .D(n7_adj_4250), .S(n8_adj_4251));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(CLK_c), 
            .D(n7_adj_4252), .S(n8_adj_4253));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(CLK_c), 
            .D(n7_adj_4254), .S(n8_adj_4255));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(CLK_c), 
            .D(n7_adj_4256), .S(n8_adj_4257));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(CLK_c), 
            .D(n35317), .S(n36148));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(CLK_c), 
            .D(n35315), .S(n36146));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(CLK_c), 
            .D(n7_adj_4258), .S(n8_adj_4259));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(CLK_c), 
            .D(n45081), .S(n44979));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(CLK_c), 
            .D(n7_adj_4260), .S(n8_adj_4261));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(CLK_c), 
            .D(n7_adj_4262), .S(n8_adj_4263));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(CLK_c), 
            .D(n35313), .S(n36144));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(CLK_c), 
            .D(n45077), .S(n45017));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(CLK_c), 
            .D(n35311), .S(n36142));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i34844_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50326));
    defparam i34844_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(CLK_c), 
            .D(n45073), .S(n44977));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(CLK_c), 
            .D(n7_adj_4264), .S(n8_adj_4265));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16313_3_lut_4_lut (.I0(n10_adj_4245), .I1(n45606), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29835));
    defparam i16313_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(CLK_c), 
            .D(n45069), .S(n44975));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(CLK_c), 
            .D(n45065), .S(n45019));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(CLK_c), 
            .D(n45061), .S(n44965));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(CLK_c), 
            .D(n35309), .S(n44963));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(CLK_c), 
            .D(n44957), .S(n44983));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i34845_4_lut (.I0(n50326), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n50327));
    defparam i34845_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i34843_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50325));
    defparam i34843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_892 (.I0(n45811), .I1(n45667), .I2(n43663), .I3(n46244), 
            .O(n10_adj_4266));
    defparam i4_4_lut_adj_892.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_893 (.I0(n3_adj_4267), .I1(n45726), .I2(n10_adj_4266), 
            .I3(n45661), .O(n13));
    defparam i3_4_lut_adj_893.LUT_INIT = 16'hebbe;
    SB_LUT4 i6_4_lut_adj_894 (.I0(n11), .I1(n42840), .I2(Kp_23__N_1237), 
            .I3(\data_in_frame[7] [2]), .O(n16_adj_4268));
    defparam i6_4_lut_adj_894.LUT_INIT = 16'hbffb;
    SB_LUT4 i1_2_lut_3_lut_adj_895 (.I0(n45638), .I1(n45610), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(GND_net), .O(n5_adj_4269));
    defparam i1_2_lut_3_lut_adj_895.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_896 (.I0(n13), .I1(n28657), .I2(n45923), .I3(n46014), 
            .O(n17_adj_4270));
    defparam i7_4_lut_adj_896.LUT_INIT = 16'hfeef;
    SB_LUT4 i16314_3_lut_4_lut (.I0(n10_adj_4245), .I1(n45606), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n29836));
    defparam i16314_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_897 (.I0(n17_adj_4270), .I1(n28259), .I2(n16_adj_4268), 
            .I3(n28264), .O(n48543));
    defparam i9_4_lut_adj_897.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_4_lut (.I0(n48543), .I1(n28544), .I2(n28226), .I3(n28232), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_898 (.I0(n28368), .I1(n12), .I2(n4_adj_4271), 
            .I3(n28537), .O(n31));
    defparam i6_4_lut_adj_898.LUT_INIT = 16'hfffe;
    SB_LUT4 i21833_2_lut (.I0(n31), .I1(n25302), .I2(GND_net), .I3(GND_net), 
            .O(n35344));
    defparam i21833_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i8336_3_lut (.I0(n31_adj_4272), .I1(n31), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n24851));   // verilog/coms.v(145[4] 299[11])
    defparam i8336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut (.I0(n24851), .I1(\FRAME_MATCHER.state [3]), .I2(\FRAME_MATCHER.state [2]), 
            .I3(GND_net), .O(n10_adj_4273));
    defparam i3_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_2_lut_adj_899 (.I0(n25302), .I1(n36131), .I2(GND_net), 
            .I3(GND_net), .O(n9));
    defparam i2_2_lut_adj_899.LUT_INIT = 16'heeee;
    SB_LUT4 i36863_4_lut (.I0(n36340), .I1(n9), .I2(n5_adj_4269), .I3(n10_adj_4273), 
            .O(n29116));
    defparam i36863_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_3_lut_4_lut_adj_900 (.I0(n45638), .I1(n45610), .I2(n36131), 
            .I3(n36340), .O(n36612));
    defparam i2_3_lut_4_lut_adj_900.LUT_INIT = 16'hfffe;
    SB_LUT4 i36059_2_lut (.I0(n53296), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51369));
    defparam i36059_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34808_4_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n50290));
    defparam i34808_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i36532_3_lut (.I0(n53116), .I1(n50290), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n52015));
    defparam i36532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16315_3_lut_4_lut (.I0(n10_adj_4245), .I1(n45606), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n29837));
    defparam i16315_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34835_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50317));
    defparam i34835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34836_4_lut (.I0(n50317), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n50318));
    defparam i34836_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i34834_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50316));
    defparam i34834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16316_3_lut_4_lut (.I0(n10_adj_4245), .I1(n45606), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n29838));
    defparam i16316_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16317_3_lut_4_lut (.I0(n10_adj_4245), .I1(n45606), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n29839));
    defparam i16317_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i35980_2_lut (.I0(n53308), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51336));
    defparam i35980_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16302_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45620), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29824));
    defparam i16302_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16303_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45620), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n29825));
    defparam i16303_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16304_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45620), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n29826));
    defparam i16304_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16305_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45620), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n29827));
    defparam i16305_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16306_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45620), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n29828));
    defparam i16306_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16307_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45620), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n29829));
    defparam i16307_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(CLK_c), 
            .E(n29243), .D(n45957));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(CLK_c), 
            .E(n29243), .D(n47924));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(CLK_c), 
            .E(n29243), .D(n45843));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(CLK_c), 
            .E(n29243), .D(n47539));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(CLK_c), 
            .E(n29243), .D(n28364));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(CLK_c), 
            .E(n29243), .D(n47712));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(CLK_c), 
            .E(n29243), .D(n47585));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(CLK_c), 
            .E(n29243), .D(n45841));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(CLK_c), 
            .E(n29243), .D(n47083));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(CLK_c), 
            .E(n29243), .D(n47535));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(CLK_c), 
            .E(n29243), .D(n47334));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(CLK_c), 
            .E(n29243), .D(n48369));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(CLK_c), 
            .E(n29243), .D(n47676));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(CLK_c), 
            .E(n29243), .D(n47312));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(CLK_c), 
            .E(n29243), .D(n48140));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(CLK_c), 
            .E(n29243), .D(n47307));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16308_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45620), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n29830));
    defparam i16308_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16309_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45620), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29831));
    defparam i16309_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n51867), .I2(n51366), .I3(byte_transmit_counter[4]), .O(n53311));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n53311_bdd_4_lut (.I0(n53311), .I1(n53200), .I2(n7_adj_4236), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n53311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n53305));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n53305_bdd_4_lut (.I0(n53305), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n53308));
    defparam n53305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37786 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n53299));
    defparam byte_transmit_counter_0__bdd_4_lut_37786.LUT_INIT = 16'he4aa;
    SB_LUT4 n53299_bdd_4_lut (.I0(n53299), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n53302));
    defparam n53299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37781 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n53293));
    defparam byte_transmit_counter_0__bdd_4_lut_37781.LUT_INIT = 16'he4aa;
    SB_LUT4 n53293_bdd_4_lut (.I0(n53293), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n53296));
    defparam n53293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 equal_287_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4274));   // verilog/coms.v(154[7:23])
    defparam equal_287_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37776 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n53287));
    defparam byte_transmit_counter_0__bdd_4_lut_37776.LUT_INIT = 16'he4aa;
    SB_LUT4 n53287_bdd_4_lut (.I0(n53287), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n53290));
    defparam n53287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37771 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n53281));
    defparam byte_transmit_counter_0__bdd_4_lut_37771.LUT_INIT = 16'he4aa;
    SB_LUT4 n53281_bdd_4_lut (.I0(n53281), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n53284));
    defparam n53281_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37766 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n53275));
    defparam byte_transmit_counter_0__bdd_4_lut_37766.LUT_INIT = 16'he4aa;
    SB_LUT4 n53275_bdd_4_lut (.I0(n53275), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n53278));
    defparam n53275_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(CLK_c), 
            .D(n2_adj_4275), .S(n3_adj_4276));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_278_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4277));   // verilog/coms.v(154[7:23])
    defparam equal_278_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_4278), .S(n3_adj_4279));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_4280), .S(n3_adj_4281));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_4282), .S(n3_adj_4283));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n2_adj_4284), .S(n3_adj_4285));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n2_adj_4286), .S(n3_adj_4287));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n2_adj_4288), .S(n3_adj_4289));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n2_adj_4290), .S(n3_adj_4291));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n2_adj_4292), .S(n3_adj_4293));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n2_adj_4294), .S(n3_adj_4295));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n2_adj_4296), .S(n3_adj_4297));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n2_adj_4298), .S(n3_adj_4299));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n2_adj_4300), .S(n3_adj_4301));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n2_adj_4302), .S(n3_adj_4303));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n2_adj_4304), .S(n3_adj_4305));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n2_adj_4306), .S(n3_adj_4307));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n2_adj_4308), .S(n3_adj_4309));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n2_adj_4310), .S(n3_adj_4311));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n2_adj_4312), .S(n3_adj_4313));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n2_adj_4314), .S(n3_adj_4315));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n2_adj_4316), .S(n3_adj_4317));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n2_adj_4221), .S(n3_adj_4318));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n2_adj_4226), .S(n3_adj_4319));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n2_adj_4228), .S(n3_adj_4320));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_4231), .S(n3_adj_4321));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_4238), .S(n3_adj_4322));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_4239), .S(n3_adj_4323));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_4240), .S(n3_adj_4324));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2_adj_4241), .S(n3_adj_4325));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_4242), .S(n3_adj_4326));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_4243), .S(n3_adj_4327));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16157_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45628), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n29679));
    defparam i16157_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16150_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45628), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n29672));
    defparam i16150_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16151_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45628), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n29673));
    defparam i16151_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16152_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45628), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n29674));
    defparam i16152_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16153_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45628), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n29675));
    defparam i16153_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16154_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45628), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n29676));
    defparam i16154_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i36931_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n39690));   // verilog/coms.v(127[12] 300[6])
    defparam i36931_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i16155_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45628), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n29677));
    defparam i16155_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[19] [1]), .O(n6561));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_901 (.I0(\FRAME_MATCHER.state [3]), .I1(n36614), 
            .I2(GND_net), .I3(GND_net), .O(n39678));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_901.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[2]), 
            .I2(byte_transmit_counter[0]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_4329));   // verilog/coms.v(102[12:33])
    defparam i1_4_lut.LUT_INIT = 16'ha888;
    SB_LUT4 i2_2_lut_adj_902 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4330));   // verilog/coms.v(102[12:33])
    defparam i2_2_lut_adj_902.LUT_INIT = 16'heeee;
    SB_LUT4 i36989_4_lut (.I0(byte_transmit_counter[3]), .I1(n6_adj_4330), 
            .I2(byte_transmit_counter[5]), .I3(n4_adj_4329), .O(tx_transmit_N_3513));
    defparam i36989_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 i1_4_lut_adj_903 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n4_c));
    defparam i1_4_lut_adj_903.LUT_INIT = 16'h5554;
    SB_LUT4 i16156_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45628), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n29678));
    defparam i16156_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[19] [2]), .O(n6562));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1817_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[19] [3]), .O(n6563));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16294_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45620), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n29816));
    defparam i16294_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16295_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45620), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n29817));
    defparam i16295_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16296_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45620), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n29818));
    defparam i16296_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16297_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45620), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n29819));
    defparam i16297_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_904 (.I0(tx_transmit_N_3513), .I1(n39678), .I2(n8_adj_4331), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n5426[0]));
    defparam i1_4_lut_adj_904.LUT_INIT = 16'heccc;
    SB_LUT4 i16298_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45620), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n29820));
    defparam i16298_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16299_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45620), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n29821));
    defparam i16299_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16300_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45620), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n29822));
    defparam i16300_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16301_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45620), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n29823));
    defparam i16301_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37761 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n53269));
    defparam byte_transmit_counter_0__bdd_4_lut_37761.LUT_INIT = 16'he4aa;
    SB_LUT4 n53269_bdd_4_lut (.I0(n53269), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n53272));
    defparam n53269_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37756 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n53263));
    defparam byte_transmit_counter_0__bdd_4_lut_37756.LUT_INIT = 16'he4aa;
    SB_LUT4 n53263_bdd_4_lut (.I0(n53263), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n53266));
    defparam n53263_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37791 (.I0(byte_transmit_counter[3]), 
            .I1(n53146), .I2(n51336), .I3(byte_transmit_counter[4]), .O(n53257));
    defparam byte_transmit_counter_3__bdd_4_lut_37791.LUT_INIT = 16'he4aa;
    SB_LUT4 n53257_bdd_4_lut (.I0(n53257), .I1(n53176), .I2(n7_adj_4237), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n53257_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37746 (.I0(byte_transmit_counter[3]), 
            .I1(n52015), .I2(n51369), .I3(byte_transmit_counter[4]), .O(n53251));
    defparam byte_transmit_counter_3__bdd_4_lut_37746.LUT_INIT = 16'he4aa;
    SB_LUT4 n53251_bdd_4_lut (.I0(n53251), .I1(n53218), .I2(n7_adj_4235), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n53251_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37741 (.I0(byte_transmit_counter[3]), 
            .I1(n52013), .I2(n51372), .I3(byte_transmit_counter[4]), .O(n53245));
    defparam byte_transmit_counter_3__bdd_4_lut_37741.LUT_INIT = 16'he4aa;
    SB_LUT4 n53245_bdd_4_lut (.I0(n53245), .I1(n53158), .I2(n7_adj_4234), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n53245_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37736 (.I0(byte_transmit_counter[3]), 
            .I1(n52011), .I2(n51363), .I3(byte_transmit_counter[4]), .O(n53239));
    defparam byte_transmit_counter_3__bdd_4_lut_37736.LUT_INIT = 16'he4aa;
    SB_LUT4 n53239_bdd_4_lut (.I0(n53239), .I1(n53194), .I2(n7_adj_4233), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n53239_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37731 (.I0(byte_transmit_counter[3]), 
            .I1(n52009), .I2(n51360), .I3(byte_transmit_counter[4]), .O(n53233));
    defparam byte_transmit_counter_3__bdd_4_lut_37731.LUT_INIT = 16'he4aa;
    SB_LUT4 n53233_bdd_4_lut (.I0(n53233), .I1(n53188), .I2(n7_adj_4232), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n53233_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37726 (.I0(byte_transmit_counter[3]), 
            .I1(n52007), .I2(n51357), .I3(byte_transmit_counter[4]), .O(n53227));
    defparam byte_transmit_counter_3__bdd_4_lut_37726.LUT_INIT = 16'he4aa;
    SB_LUT4 n53227_bdd_4_lut (.I0(n53227), .I1(n53182), .I2(n7_adj_4230), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n53227_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16286_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45620), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n29808));
    defparam i16286_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16287_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45620), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n29809));
    defparam i16287_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16288_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45620), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n29810));
    defparam i16288_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[19] [4]), .O(n6564));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16289_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45620), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n29811));
    defparam i16289_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16290_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45620), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n29812));
    defparam i16290_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n40495), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n40494), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_8 (.CI(n40494), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n40495));
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n40493), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_7 (.CI(n40493), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n40494));
    SB_LUT4 i16291_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45620), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n29813));
    defparam i16291_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16292_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45620), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n29814));
    defparam i16292_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16293_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45620), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n29815));
    defparam i16293_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_292_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4328));   // verilog/coms.v(154[7:23])
    defparam equal_292_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 mux_1817_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[19] [5]), .O(n6565));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 equal_293_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4332));   // verilog/coms.v(154[7:23])
    defparam equal_293_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n40492), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37721 (.I0(byte_transmit_counter[3]), 
            .I1(n52005), .I2(n51354), .I3(byte_transmit_counter[4]), .O(n53221));
    defparam byte_transmit_counter_3__bdd_4_lut_37721.LUT_INIT = 16'he4aa;
    SB_CARRY add_3971_6 (.CI(n40492), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n40493));
    SB_LUT4 i1_2_lut_adj_905 (.I0(\FRAME_MATCHER.state [3]), .I1(n27968), 
            .I2(GND_net), .I3(GND_net), .O(n63_adj_10));   // verilog/coms.v(201[5:24])
    defparam i1_2_lut_adj_905.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_906 (.I0(\FRAME_MATCHER.state [2]), .I1(n39684), 
            .I2(GND_net), .I3(GND_net), .O(n39685));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_906.LUT_INIT = 16'hdddd;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n40491), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21819_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3616[0]), .I2(GND_net), 
            .I3(GND_net), .O(n35330));
    defparam i21819_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_3971_5 (.CI(n40491), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n40492));
    SB_LUT4 i1_2_lut_adj_907 (.I0(n29149), .I1(n39686), .I2(GND_net), 
            .I3(GND_net), .O(n39687));
    defparam i1_2_lut_adj_907.LUT_INIT = 16'h8888;
    SB_LUT4 i36866_4_lut (.I0(n39684), .I1(n63_adj_10), .I2(n6_adj_4333), 
            .I3(\FRAME_MATCHER.state [1]), .O(n29149));
    defparam i36866_4_lut.LUT_INIT = 16'h3733;
    SB_LUT4 i16278_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45620), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n29800));
    defparam i16278_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16279_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45620), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n29801));
    defparam i16279_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16280_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45620), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n29802));
    defparam i16280_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34850_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50332));
    defparam i34850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34851_4_lut (.I0(n50332), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n50333));
    defparam i34851_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i34849_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50331));
    defparam i34849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16281_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45620), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n29803));
    defparam i16281_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16282_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45620), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n29804));
    defparam i16282_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n40490), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36062_2_lut (.I0(n53290), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51366));
    defparam i36062_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_3971_4 (.CI(n40490), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n40491));
    SB_LUT4 i16283_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45620), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n29805));
    defparam i16283_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34811_4_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n50293));
    defparam i34811_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i36384_3_lut (.I0(n53122), .I1(n50293), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n51867));
    defparam i36384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16284_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45620), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n29806));
    defparam i16284_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16285_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45620), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n29807));
    defparam i16285_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n40489), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_3 (.CI(n40489), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n40490));
    SB_LUT4 i4_4_lut_adj_908 (.I0(n28111), .I1(n45860), .I2(n45848), .I3(n6_adj_4334), 
            .O(n47307));
    defparam i4_4_lut_adj_908.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_909 (.I0(n46362), .I1(n43866), .I2(n43923), .I3(n46335), 
            .O(n15_adj_4335));
    defparam i6_4_lut_adj_909.LUT_INIT = 16'h9669;
    SB_LUT4 i16270_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45620), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n29792));
    defparam i16270_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16271_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45620), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n29793));
    defparam i16271_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_910 (.I0(n15_adj_4335), .I1(n45959), .I2(n14_adj_4337), 
            .I3(\data_out_frame[23] [7]), .O(n48140));
    defparam i8_4_lut_adj_910.LUT_INIT = 16'h9669;
    SB_LUT4 i16272_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45620), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n29794));
    defparam i16272_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_911 (.I0(\data_out_frame[24] [1]), .I1(n46141), 
            .I2(n45884), .I3(n43805), .O(n47312));
    defparam i3_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(n45979), .I1(n46222), .I2(n43866), .I3(GND_net), 
            .O(n47676));
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i16273_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45620), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n29795));
    defparam i16273_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16274_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45620), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n29796));
    defparam i16274_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3513), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3513), 
            .CO(n40489));
    SB_LUT4 i1_2_lut_adj_912 (.I0(n43876), .I1(n42781), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4338));
    defparam i1_2_lut_adj_912.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_33_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n40488), .O(n2_adj_4275)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_913 (.I0(n45862), .I1(n45884), .I2(\data_out_frame[24] [2]), 
            .I3(n6_adj_4338), .O(n48369));
    defparam i4_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_32_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n40487), .O(n2_adj_4278)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16275_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45620), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n29797));
    defparam i16275_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_914 (.I0(\data_out_frame[20] [0]), .I1(n28526), 
            .I2(n45697), .I3(n6_adj_4339), .O(n42781));
    defparam i4_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_915 (.I0(\data_out_frame[24] [4]), .I1(n46207), 
            .I2(n45959), .I3(n42781), .O(n47535));
    defparam i3_4_lut_adj_915.LUT_INIT = 16'h9669;
    SB_LUT4 i21934_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i21934_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_3_lut_adj_916 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[24] [0]), 
            .I2(\data_out_frame[25] [2]), .I3(GND_net), .O(n14_adj_4341));
    defparam i5_3_lut_adj_916.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_917 (.I0(n46316), .I1(n43593), .I2(n43920), .I3(n46207), 
            .O(n15_adj_4342));
    defparam i6_4_lut_adj_917.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_918 (.I0(n15_adj_4342), .I1(n27992), .I2(n14_adj_4341), 
            .I3(\data_out_frame[25] [0]), .O(n47083));
    defparam i8_4_lut_adj_918.LUT_INIT = 16'h6996;
    SB_CARRY add_43_32 (.CI(n40487), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n40488));
    SB_LUT4 i16276_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45620), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n29798));
    defparam i16276_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_919 (.I0(n46213), .I1(n45840), .I2(n46231), .I3(n43920), 
            .O(n45841));
    defparam i1_4_lut_adj_919.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1817_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[19] [6]), .O(n6566));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_920 (.I0(\data_out_frame[20] [1]), .I1(n43883), 
            .I2(GND_net), .I3(GND_net), .O(n43920));
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_921 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(\data_out_frame[23] [7]), .I3(GND_net), .O(n46222));
    defparam i2_3_lut_adj_921.LUT_INIT = 16'h9696;
    SB_LUT4 n53221_bdd_4_lut (.I0(n53221), .I1(n53164), .I2(n7_adj_4229), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n53221_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n50412), .I2(n50413), .I3(byte_transmit_counter[2]), .O(n53215));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n53215_bdd_4_lut (.I0(n53215), .I1(n50407), .I2(n50406), .I3(byte_transmit_counter[2]), 
            .O(n53218));
    defparam n53215_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37712 (.I0(byte_transmit_counter[1]), 
            .I1(n50310), .I2(n50311), .I3(byte_transmit_counter[2]), .O(n53197));
    defparam byte_transmit_counter_1__bdd_4_lut_37712.LUT_INIT = 16'he4aa;
    SB_LUT4 n53197_bdd_4_lut (.I0(n53197), .I1(n50383), .I2(n50382), .I3(byte_transmit_counter[2]), 
            .O(n53200));
    defparam n53197_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_922 (.I0(n28418), .I1(n45674), .I2(\data_out_frame[19] [7]), 
            .I3(\data_out_frame[17] [5]), .O(n46210));
    defparam i3_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_LUT4 i16277_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45620), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n29799));
    defparam i16277_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16262_3_lut_4_lut (.I0(n36193), .I1(n45620), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n29784));
    defparam i16262_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16263_3_lut_4_lut (.I0(n36193), .I1(n45620), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n29785));
    defparam i16263_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_923 (.I0(n42913), .I1(\data_out_frame[24] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43805));
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h6666;
    SB_LUT4 i16264_3_lut_4_lut (.I0(n36193), .I1(n45620), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n29786));
    defparam i16264_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37698 (.I0(byte_transmit_counter[1]), 
            .I1(n50346), .I2(n50347), .I3(byte_transmit_counter[2]), .O(n53191));
    defparam byte_transmit_counter_1__bdd_4_lut_37698.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_924 (.I0(n43437), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43936));
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_925 (.I0(n43805), .I1(\data_out_frame[23] [5]), 
            .I2(n42923), .I3(n45959), .O(n46362));
    defparam i3_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_LUT4 i16265_3_lut_4_lut (.I0(n36193), .I1(n45620), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n29787));
    defparam i16265_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12_4_lut (.I0(n46144), .I1(n43850), .I2(\data_out_frame[24] [6]), 
            .I3(n43936), .O(n29));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_926 (.I0(n46228), .I1(n28114), .I2(\data_out_frame[20] [1]), 
            .I3(\data_out_frame[20] [2]), .O(n20_adj_4343));
    defparam i3_4_lut_adj_926.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(n42875), .I1(\data_out_frame[24] [5]), .I2(n28149), 
            .I3(n46222), .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_927 (.I0(n29), .I1(n42909), .I2(n26), .I3(\data_out_frame[23] [6]), 
            .O(n32));
    defparam i15_4_lut_adj_927.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_928 (.I0(n19_adj_4225), .I1(n32), .I2(n28), 
            .I3(n20_adj_4343), .O(n43593));
    defparam i16_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i16266_3_lut_4_lut (.I0(n36193), .I1(n45620), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n29788));
    defparam i16266_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_929 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[25] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n28111));
    defparam i1_2_lut_adj_929.LUT_INIT = 16'h6666;
    SB_LUT4 n53191_bdd_4_lut (.I0(n53191), .I1(n50380), .I2(n50379), .I3(byte_transmit_counter[2]), 
            .O(n53194));
    defparam n53191_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37693 (.I0(byte_transmit_counter[1]), 
            .I1(n50385), .I2(n50386), .I3(byte_transmit_counter[2]), .O(n53185));
    defparam byte_transmit_counter_1__bdd_4_lut_37693.LUT_INIT = 16'he4aa;
    SB_LUT4 n53185_bdd_4_lut (.I0(n53185), .I1(n50377), .I2(n50376), .I3(byte_transmit_counter[2]), 
            .O(n53188));
    defparam n53185_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37688 (.I0(byte_transmit_counter[1]), 
            .I1(n50415), .I2(n50416), .I3(byte_transmit_counter[2]), .O(n53179));
    defparam byte_transmit_counter_1__bdd_4_lut_37688.LUT_INIT = 16'he4aa;
    SB_LUT4 n53179_bdd_4_lut (.I0(n53179), .I1(n50443), .I2(n50442), .I3(byte_transmit_counter[2]), 
            .O(n53182));
    defparam n53179_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_43_31_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n40486), .O(n2_adj_4280)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_930 (.I0(n42807), .I1(n45843), .I2(n6_adj_4344), 
            .I3(n42887), .O(n45840));
    defparam i1_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i16267_3_lut_4_lut (.I0(n36193), .I1(n45620), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n29789));
    defparam i16267_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_931 (.I0(n43593), .I1(n46362), .I2(GND_net), 
            .I3(GND_net), .O(n46213));
    defparam i1_2_lut_adj_931.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_932 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46194));
    defparam i1_2_lut_adj_932.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_933 (.I0(\data_out_frame[17] [6]), .I1(n28526), 
            .I2(GND_net), .I3(GND_net), .O(n46250));
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_934 (.I0(\data_out_frame[18] [1]), .I1(n46250), 
            .I2(n46194), .I3(n45930), .O(n43850));
    defparam i3_4_lut_adj_934.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_935 (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[25] [0]), 
            .I2(n43868), .I3(n6), .O(n46231));
    defparam i4_4_lut_adj_935.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_936 (.I0(\data_out_frame[20] [2]), .I1(n43850), 
            .I2(GND_net), .I3(GND_net), .O(n43927));
    defparam i1_2_lut_adj_936.LUT_INIT = 16'h6666;
    SB_CARRY add_43_31 (.CI(n40486), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n40487));
    SB_LUT4 i5_4_lut_adj_937 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [5]), 
            .I2(n28331), .I3(\data_out_frame[15] [4]), .O(n12_adj_4345));
    defparam i5_4_lut_adj_937.LUT_INIT = 16'h6996;
    SB_LUT4 i16268_3_lut_4_lut (.I0(n36193), .I1(n45620), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n29790));
    defparam i16268_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_938 (.I0(\data_out_frame[16] [0]), .I1(n12_adj_4345), 
            .I2(n42822), .I3(\data_out_frame[13] [6]), .O(n45930));
    defparam i6_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_939 (.I0(n45930), .I1(n46190), .I2(\data_out_frame[18] [1]), 
            .I3(n28342), .O(n45947));
    defparam i3_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28114));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_941 (.I0(n46178), .I1(n42897), .I2(n45985), .I3(n42958), 
            .O(n46228));
    defparam i3_4_lut_adj_941.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_942 (.I0(n27578), .I1(n46228), .I2(n28114), .I3(n46144), 
            .O(n42807));
    defparam i2_4_lut_adj_942.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37683 (.I0(byte_transmit_counter[1]), 
            .I1(n50373), .I2(n50374), .I3(byte_transmit_counter[2]), .O(n53173));
    defparam byte_transmit_counter_1__bdd_4_lut_37683.LUT_INIT = 16'he4aa;
    SB_LUT4 n53173_bdd_4_lut (.I0(n53173), .I1(n50371), .I2(n50370), .I3(byte_transmit_counter[2]), 
            .O(n53176));
    defparam n53173_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37678 (.I0(byte_transmit_counter[1]), 
            .I1(n50367), .I2(n50368), .I3(byte_transmit_counter[2]), .O(n53161));
    defparam byte_transmit_counter_1__bdd_4_lut_37678.LUT_INIT = 16'he4aa;
    SB_LUT4 n53161_bdd_4_lut (.I0(n53161), .I1(n50437), .I2(n50436), .I3(byte_transmit_counter[2]), 
            .O(n53164));
    defparam n53161_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16269_3_lut_4_lut (.I0(n36193), .I1(n45620), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n29791));
    defparam i16269_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_943 (.I0(n42897), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n45854));
    defparam i1_2_lut_adj_943.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1817_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[19] [7]), .O(n6567));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_944 (.I0(n28077), .I1(\data_out_frame[13] [6]), 
            .I2(n45916), .I3(n6_adj_4346), .O(n28342));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_LUT4 i16254_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45612), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n29776));
    defparam i16254_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_30_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n40485), .O(n2_adj_4282)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_945 (.I0(\data_out_frame[25] [2]), .I1(n27578), 
            .I2(n45854), .I3(n6_adj_4347), .O(n42887));
    defparam i4_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_CARRY add_43_30 (.CI(n40485), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n40486));
    SB_LUT4 i16255_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45612), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n29777));
    defparam i16255_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[18] [0]), .O(n6568));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16256_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45612), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n29778));
    defparam i16256_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i22668_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n36193));
    defparam i22668_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 equal_283_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4336));
    defparam equal_283_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i2_3_lut_adj_946 (.I0(\data_out_frame[25] [3]), .I1(n43846), 
            .I2(n42887), .I3(GND_net), .O(n47539));
    defparam i2_3_lut_adj_946.LUT_INIT = 16'h6969;
    SB_LUT4 add_43_29_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n40484), .O(n2_adj_4284)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_29 (.CI(n40484), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n40485));
    SB_LUT4 add_43_28_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n40483), .O(n2_adj_4286)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_28 (.CI(n40483), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n40484));
    SB_LUT4 i16257_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45612), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n29779));
    defparam i16257_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_947 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27992));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_947.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1817_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[18] [1]), .O(n6569));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_948 (.I0(\data_out_frame[23] [2]), .I1(n45744), 
            .I2(n46082), .I3(n42958), .O(n43846));
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_949 (.I0(n43846), .I1(n47119), .I2(n27992), .I3(GND_net), 
            .O(n45843));
    defparam i2_3_lut_adj_949.LUT_INIT = 16'h9696;
    SB_LUT4 i16258_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45612), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n29780));
    defparam i16258_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16259_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45612), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n29781));
    defparam i16259_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_950 (.I0(\data_out_frame[20] [6]), .I1(n28584), 
            .I2(n45749), .I3(\data_out_frame[18] [5]), .O(n45744));
    defparam i3_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i16260_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45612), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n29782));
    defparam i16260_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[18] [2]), .O(n6570));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16261_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45612), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n29783));
    defparam i16261_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\data_out_frame[23] [3]), .I1(\data_out_frame[23] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28155));
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_952 (.I0(n42897), .I1(n45859), .I2(n28155), .I3(n27578), 
            .O(n47119));
    defparam i3_4_lut_adj_952.LUT_INIT = 16'h6996;
    SB_LUT4 i16246_3_lut_4_lut (.I0(n10_adj_4244), .I1(n45606), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n29768));
    defparam i16246_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[18] [3]), .O(n6571));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_953 (.I0(\data_out_frame[25] [5]), .I1(n43943), 
            .I2(\data_out_frame[25] [4]), .I3(n47119), .O(n47924));
    defparam i3_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i16247_3_lut_4_lut (.I0(n10_adj_4244), .I1(n45606), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n29769));
    defparam i16247_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_954 (.I0(n45707), .I1(n46056), .I2(GND_net), 
            .I3(GND_net), .O(n28193));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_955 (.I0(\data_out_frame[18] [4]), .I1(n28331), 
            .I2(n1699), .I3(n28353), .O(n10_adj_4348));
    defparam i4_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_956 (.I0(n46300), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[18] [3]), .I3(n46371), .O(n10_adj_4349));
    defparam i4_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_957 (.I0(n46203), .I1(n10_adj_4349), .I2(n42820), 
            .I3(GND_net), .O(n46348));
    defparam i5_3_lut_adj_957.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_958 (.I0(n46348), .I1(n45749), .I2(GND_net), 
            .I3(GND_net), .O(n43235));
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_959 (.I0(\data_out_frame[13] [7]), .I1(n28193), 
            .I2(\data_out_frame[16] [1]), .I3(\data_out_frame[18] [2]), 
            .O(n45916));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_960 (.I0(n42822), .I1(\data_out_frame[10] [5]), 
            .I2(n26026), .I3(\data_out_frame[8] [3]), .O(n24));
    defparam i10_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_961 (.I0(n45942), .I1(n1513), .I2(n1516), .I3(\data_out_frame[12] [0]), 
            .O(n22));
    defparam i8_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_962 (.I0(n27502), .I1(n24), .I2(n18_adj_4350), 
            .I3(n1510), .O(n26_adj_4351));
    defparam i12_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n1241), .I1(n26_adj_4351), .I2(n22), .I3(\data_out_frame[8] [4]), 
            .O(n46203));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_963 (.I0(\data_out_frame[13] [7]), .I1(n46203), 
            .I2(GND_net), .I3(GND_net), .O(n28353));
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_964 (.I0(n1519), .I1(n45664), .I2(GND_net), .I3(GND_net), 
            .O(n28466));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_965 (.I0(n28014), .I1(\data_out_frame[15] [1]), 
            .I2(n46216), .I3(\data_out_frame[17] [1]), .O(n10_adj_4352));
    defparam i4_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_966 (.I0(\data_out_frame[16] [7]), .I1(n10_adj_4352), 
            .I2(\data_out_frame[14] [5]), .I3(GND_net), .O(n45867));
    defparam i5_3_lut_adj_966.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_967 (.I0(n45674), .I1(n45872), .I2(\data_out_frame[13] [1]), 
            .I3(n28466), .O(n12_adj_4353));
    defparam i5_4_lut_adj_967.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_968 (.I0(n28006), .I1(n12_adj_4353), .I2(n46150), 
            .I3(\data_out_frame[14] [7]), .O(n43437));
    defparam i6_4_lut_adj_968.LUT_INIT = 16'h6996;
    SB_LUT4 i16248_3_lut_4_lut (.I0(n10_adj_4244), .I1(n45606), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n29770));
    defparam i16248_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_969 (.I0(n28074), .I1(n45688), .I2(n46353), .I3(n6_adj_4354), 
            .O(n46263));
    defparam i4_4_lut_adj_969.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_970 (.I0(\data_in_frame[15] [7]), .I1(n46263), 
            .I2(\data_in_frame[16] [1]), .I3(GND_net), .O(n46046));
    defparam i2_3_lut_adj_970.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_971 (.I0(n46024), .I1(n46294), .I2(n8_adj_4355), 
            .I3(\data_in_frame[3] [7]), .O(n17_adj_4356));
    defparam i4_4_lut_adj_971.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_972 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[5] [0]), 
            .I2(n46345), .I3(\data_in_frame[11] [5]), .O(n21));
    defparam i8_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_973 (.I0(n28022), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(n45872), .O(n45697));
    defparam i3_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(\data_in_frame[5] [2]), .I1(n4_adj_4357), .I2(\data_in_frame[13] [7]), 
            .I3(GND_net), .O(n20_adj_4358));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_974 (.I0(n21), .I1(n17_adj_4356), .I2(n45818), 
            .I3(n29001), .O(n24_adj_4359));
    defparam i11_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i16249_3_lut_4_lut (.I0(n10_adj_4244), .I1(n45606), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n29771));
    defparam i16249_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_975 (.I0(\data_out_frame[19] [5]), .I1(n43437), 
            .I2(\data_out_frame[19] [3]), .I3(n45867), .O(n45979));
    defparam i3_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_976 (.I0(n28645), .I1(n24_adj_4359), .I2(n20_adj_4358), 
            .I3(\data_in_frame[2] [1]), .O(n28912));
    defparam i12_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_977 (.I0(n28912), .I1(n28129), .I2(n42915), .I3(GND_net), 
            .O(n46225));
    defparam i2_3_lut_adj_977.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_978 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n45896));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_978.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_979 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46277));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_980 (.I0(\data_in_frame[18] [1]), .I1(n43591), 
            .I2(\data_in_frame[18] [2]), .I3(GND_net), .O(n46260));
    defparam i2_3_lut_adj_980.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_981 (.I0(n43819), .I1(\data_in_frame[16] [5]), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n45950));
    defparam i2_3_lut_adj_981.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_982 (.I0(\data_in_frame[14] [4]), .I1(n45893), 
            .I2(n42581), .I3(\data_in_frame[12] [2]), .O(n28279));
    defparam i3_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(71[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_983 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(n45764), .I3(\data_out_frame[6] [4]), .O(n46166));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_983.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_984 (.I0(\data_in_frame[18] [6]), .I1(n28279), 
            .I2(n45950), .I3(GND_net), .O(n46156));
    defparam i1_3_lut_adj_984.LUT_INIT = 16'h6969;
    SB_LUT4 i10_4_lut_adj_985 (.I0(\data_out_frame[9] [7]), .I1(n46285), 
            .I2(\data_out_frame[9] [5]), .I3(\data_out_frame[7] [4]), .O(n28_adj_4360));
    defparam i10_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_986 (.I0(\data_in_frame[9] [6]), .I1(n28264), .I2(GND_net), 
            .I3(GND_net), .O(n45890));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h6666;
    SB_LUT4 i14_3_lut (.I0(\data_out_frame[5] [3]), .I1(n28_adj_4360), .I2(\data_out_frame[5] [4]), 
            .I3(GND_net), .O(n32_adj_4361));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_987 (.I0(n28447), .I1(n46187), .I2(\data_out_frame[8] [4]), 
            .I3(n45779), .O(n30));
    defparam i12_4_lut_adj_987.LUT_INIT = 16'h6996;
    SB_LUT4 i16250_3_lut_4_lut (.I0(n10_adj_4244), .I1(n45606), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n29772));
    defparam i16250_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_988 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[4] [7]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[4] [0]), .O(n31_adj_4362));
    defparam i13_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 i16251_3_lut_4_lut (.I0(n10_adj_4244), .I1(n45606), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n29773));
    defparam i16251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16252_3_lut_4_lut (.I0(n10_adj_4244), .I1(n45606), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n29774));
    defparam i16252_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_989 (.I0(\data_out_frame[8] [2]), .I1(n46099), 
            .I2(\data_out_frame[7] [1]), .I3(n28439), .O(n29_adj_4363));
    defparam i11_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut (.I0(n11_adj_4364), .I1(n42581), .I2(n46116), .I3(GND_net), 
            .O(n16_adj_4365));   // verilog/coms.v(85[17:63])
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_990 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[8] [3]), .I3(n46257), .O(n17_adj_4366));   // verilog/coms.v(85[17:63])
    defparam i7_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_991 (.I0(n29_adj_4363), .I1(n31_adj_4362), .I2(n30), 
            .I3(n32_adj_4361), .O(n48172));
    defparam i17_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_992 (.I0(n48172), .I1(n46288), .I2(n45881), .I3(n46166), 
            .O(n12_adj_4367));
    defparam i5_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_993 (.I0(n17_adj_4366), .I1(n45801), .I2(n16_adj_4365), 
            .I3(n28368), .O(n45997));   // verilog/coms.v(85[17:63])
    defparam i9_4_lut_adj_993.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_994 (.I0(\data_out_frame[11] [0]), .I1(n1241), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n8_adj_4368));
    defparam i3_3_lut_adj_994.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_995 (.I0(\data_in_frame[18] [4]), .I1(n28275), 
            .I2(\data_in_frame[18] [5]), .I3(GND_net), .O(n45953));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_995.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut (.I0(n27538), .I1(n46380), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4369));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n36137), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(n10_adj_4244), .O(n45612));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i13_4_lut_adj_996 (.I0(n45997), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[10] [0]), .O(n34));
    defparam i13_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_997 (.I0(n11_adj_4370), .I1(n8_adj_4368), .I2(\data_out_frame[10] [0]), 
            .I3(n12_adj_4367), .O(n48381));
    defparam i4_4_lut_adj_997.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_998 (.I0(\data_in_frame[11] [7]), .I1(n34), .I2(n24_adj_4369), 
            .I3(n45836), .O(n38));
    defparam i17_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_999 (.I0(n28035), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[11] [6]), .I3(n28456), .O(n28_adj_4371));
    defparam i12_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 i16253_3_lut_4_lut (.I0(n10_adj_4244), .I1(n45606), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n29775));
    defparam i16253_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1000 (.I0(\data_out_frame[11] [5]), .I1(n28068), 
            .I2(n46166), .I3(\data_out_frame[11] [7]), .O(n26_adj_4372));
    defparam i10_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1001 (.I0(n43839), .I1(n46122), .I2(n46282), 
            .I3(n46099), .O(n27));
    defparam i11_4_lut_adj_1001.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1002 (.I0(n48381), .I1(n46304), .I2(n46103), 
            .I3(\data_out_frame[10] [1]), .O(n25));
    defparam i9_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1003 (.I0(n25), .I1(n27), .I2(n26_adj_4372), 
            .I3(n28_adj_4371), .O(n26026));
    defparam i15_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(n26026), .I1(\data_out_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n45942));
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_27_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n40482), .O(n2_adj_4288)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46159));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut_adj_1006 (.I0(n45815), .I1(\data_in_frame[11] [6]), 
            .I2(Kp_23__N_981), .I3(n29001), .O(n36));
    defparam i15_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(CLK_c), .D(n30122));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(CLK_c), .D(n30121));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(CLK_c), .D(n30120));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(CLK_c), .D(n30119));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(CLK_c), .D(n30118));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(CLK_c), .D(n30117));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(CLK_c), .D(n30116));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(CLK_c), .D(n30115));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(CLK_c), .D(n30114));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(CLK_c), .D(n30113));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(CLK_c), .D(n30112));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(CLK_c), .D(n30111));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(CLK_c), .D(n30110));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(CLK_c), .D(n30109));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(CLK_c), .D(n30108));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(CLK_c), .D(n30107));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(CLK_c), .D(n30106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(CLK_c), .D(n30105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(CLK_c), .D(n30104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(CLK_c), .D(n30103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(CLK_c), .D(n30102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(CLK_c), .D(n30101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(CLK_c), .D(n30100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(CLK_c), .D(n30099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(CLK_c), .D(n30098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(CLK_c), .D(n30097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(CLK_c), .D(n30096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(CLK_c), .D(n30095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(CLK_c), .D(n30094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n30093));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(CLK_c), .D(n30092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n30091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n30090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(CLK_c), .D(n30089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(CLK_c), .D(n30088));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(CLK_c), .D(n30087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(CLK_c), .D(n30086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(CLK_c), .D(n30085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(CLK_c), .D(n30084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(CLK_c), .D(n30083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n30082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(CLK_c), .D(n30081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n30080));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(CLK_c), .D(n30079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(CLK_c), .D(n30078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(CLK_c), .D(n30077));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n30076));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(CLK_c), .D(n30075));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(CLK_c), .D(n30074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(CLK_c), .D(n30073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n30072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(CLK_c), .D(n30071));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(CLK_c), .D(n30070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(CLK_c), .D(n30069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(CLK_c), .D(n30068));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(CLK_c), .D(n30067));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(CLK_c), .D(n30066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(CLK_c), .D(n30065));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(CLK_c), .D(n30064));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(CLK_c), .D(n30063));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(CLK_c), .D(n30062));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(CLK_c), .D(n30061));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(CLK_c), .D(n30060));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(CLK_c), .D(n30059));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(CLK_c), .D(n30058));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(CLK_c), .D(n30057));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(CLK_c), .D(n30056));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(CLK_c), .D(n30055));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(CLK_c), .D(n30054));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(CLK_c), .D(n30053));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(CLK_c), .D(n30052));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(CLK_c), .D(n30051));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(CLK_c), .D(n30050));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(CLK_c), .D(n30049));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(CLK_c), .D(n30048));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(CLK_c), .D(n30047));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(CLK_c), .D(n30046));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(CLK_c), .D(n30045));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(CLK_c), .D(n30044));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(CLK_c), .D(n30043));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(CLK_c), .D(n30042));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(CLK_c), .D(n30041));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(CLK_c), .D(n30040));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(CLK_c), .D(n30039));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(CLK_c), 
           .D(n30038));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(CLK_c), 
           .D(n30037));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(CLK_c), 
           .D(n30036));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(CLK_c), 
           .D(n30035));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(CLK_c), 
           .D(n30034));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(CLK_c), 
           .D(n30033));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(CLK_c), 
           .D(n30032));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(CLK_c), 
           .D(n30031));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(CLK_c), 
           .D(n30030));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(CLK_c), 
           .D(n30029));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_27 (.CI(n40482), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n40483));
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(CLK_c), 
           .D(n30028));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(CLK_c), 
           .D(n30027));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_26_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n40481), .O(n2_adj_4290)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16_4_lut_adj_1007 (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[7] [0]), .I3(n22_adj_4373), .O(n37));
    defparam i16_4_lut_adj_1007.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1008 (.I0(\data_in_frame[12] [0]), .I1(n46092), 
            .I2(n46356), .I3(n45890), .O(n35));
    defparam i14_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n37), .I2(n36), .I3(n38), .O(n43819));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1009 (.I0(\data_in_frame[9] [3]), .I1(n45684), 
            .I2(n43009), .I3(\data_in_frame[18] [0]), .O(n46039));
    defparam i3_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1010 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[15] [5]), 
            .I2(\data_in_frame[13] [5]), .I3(GND_net), .O(n46254));
    defparam i2_3_lut_adj_1010.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1011 (.I0(n45878), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[8] [7]), .I3(\data_out_frame[4] [4]), .O(n14_adj_4374));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_1011.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(\data_in_frame[14] [2]), .I1(n46331), 
            .I2(GND_net), .I3(GND_net), .O(n46380));
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28689));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1014 (.I0(n46304), .I1(n14_adj_4374), .I2(n10_adj_4375), 
            .I3(\data_out_frame[6] [6]), .O(n28526));   // verilog/coms.v(76[16:27])
    defparam i7_4_lut_adj_1014.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_out_frame[13] [0]), .I1(n28526), 
            .I2(GND_net), .I3(GND_net), .O(n28486));
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1016 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46353));
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1017 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[14] [0]), 
            .I2(n46269), .I3(n6_adj_4376), .O(n45707));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\data_in_frame[13] [0]), .I1(n45736), 
            .I2(GND_net), .I3(GND_net), .O(n46272));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(\data_in_frame[8] [6]), .I1(Kp_23__N_1195), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4377));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1020 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[14] [7]), 
            .I2(n46272), .I3(n46077), .O(n45910));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1021 (.I0(n45741), .I1(n45825), .I2(\data_in_frame[13] [1]), 
            .I3(\data_in_frame[13] [0]), .O(n12_adj_4378));   // verilog/coms.v(76[16:43])
    defparam i5_4_lut_adj_1021.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1022 (.I0(\data_in_frame[15] [2]), .I1(n12_adj_4378), 
            .I2(n46128), .I3(n7_adj_4377), .O(n28902));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46377));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1024 (.I0(n28046), .I1(n46365), .I2(Kp_23__N_1237), 
            .I3(\data_in_frame[13] [4]), .O(n12_adj_4379));
    defparam i5_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1025 (.I0(\data_in_frame[16] [2]), .I1(n12_adj_4379), 
            .I2(n46377), .I3(\data_in_frame[15] [6]), .O(n45982));
    defparam i6_4_lut_adj_1025.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28006));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n46282));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1028 (.I0(n28902), .I1(n45910), .I2(\data_in_frame[17] [3]), 
            .I3(GND_net), .O(n28084));
    defparam i2_3_lut_adj_1028.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37668 (.I0(byte_transmit_counter[1]), 
            .I1(n50451), .I2(n50452), .I3(byte_transmit_counter[2]), .O(n53155));
    defparam byte_transmit_counter_1__bdd_4_lut_37668.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1029 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n28439));
    defparam i2_3_lut_adj_1029.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1030 (.I0(\data_in_frame[12] [0]), .I1(n45644), 
            .I2(\data_in_frame[9] [6]), .I3(GND_net), .O(n46294));
    defparam i2_3_lut_adj_1030.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(CLK_c), 
           .D(n30026));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(CLK_c), 
           .D(n30025));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(CLK_c), 
           .D(n30024));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(CLK_c), 
           .D(n30023));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(CLK_c), 
           .D(n30022));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(CLK_c), 
           .D(n30021));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(CLK_c), 
           .D(n30020));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(CLK_c), 
           .D(n30019));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(CLK_c), 
           .D(n30018));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(CLK_c), 
           .D(n30017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(CLK_c), 
           .D(n30016));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(CLK_c), 
           .D(n30015));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(CLK_c), 
           .D(n30014));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(CLK_c), 
           .D(n30013));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(CLK_c), 
           .D(n30012));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(CLK_c), 
           .D(n30011));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(CLK_c), 
           .D(n30010));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(CLK_c), 
           .D(n30009));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(CLK_c), 
           .D(n30008));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(CLK_c), 
           .D(n30007));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(CLK_c), 
           .D(n30006));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(CLK_c), 
           .D(n30005));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(CLK_c), 
           .D(n30004));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(CLK_c), 
           .D(n30003));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(CLK_c), 
           .D(n30002));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(CLK_c), 
           .D(n30001));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(CLK_c), 
           .D(n30000));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(CLK_c), 
           .D(n29999));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(CLK_c), 
           .D(n29998));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(CLK_c), 
           .D(n29997));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(CLK_c), 
           .D(n29996));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1031 (.I0(n45648), .I1(n46014), .I2(\data_in_frame[7] [7]), 
            .I3(\data_in_frame[7] [6]), .O(n12_adj_4380));
    defparam i5_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n46089));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1033 (.I0(\data_in_frame[10] [2]), .I1(n12_adj_4380), 
            .I2(n46237), .I3(\data_in_frame[8] [1]), .O(n46328));
    defparam i6_4_lut_adj_1033.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1034 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n46374));
    defparam i1_2_lut_adj_1034.LUT_INIT = 16'h6666;
    SB_CARRY add_43_26 (.CI(n40481), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n40482));
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(CLK_c), 
           .D(n29995));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(CLK_c), 
           .D(n29994));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(CLK_c), 
           .D(n29993));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(CLK_c), 
           .D(n29991));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(CLK_c), 
           .D(n29990));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(CLK_c), 
           .D(n29989));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(CLK_c), 
           .D(n29988));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(CLK_c), 
           .D(n29987));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(CLK_c), 
           .D(n29986));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1035 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[4] [1]), .I3(n6_adj_4381), .O(n1519));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(CLK_c), 
           .D(n29985));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1036 (.I0(n46181), .I1(n46277), .I2(\data_in_frame[16] [6]), 
            .I3(GND_net), .O(n46072));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1036.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(CLK_c), 
           .D(n29984));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i23_4_lut (.I0(n45851), .I1(n46072), .I2(n46386), .I3(n28259), 
            .O(n66));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1037 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4382));
    defparam i1_2_lut_adj_1037.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(CLK_c), 
           .D(n29983));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31_4_lut (.I0(n46374), .I1(n28881), .I2(n46328), .I3(n45716), 
            .O(n74));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(CLK_c), 
           .D(n29982));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i29_4_lut (.I0(n45993), .I1(n28146), .I2(n46353), .I3(n46383), 
            .O(n72));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(CLK_c), 
           .D(n29981));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1038 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[14] [5]), 
            .I2(\data_out_frame[14] [3]), .I3(n6_adj_4382), .O(n46006));
    defparam i4_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(CLK_c), 
           .D(n29980));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(CLK_c), 
           .D(n29979));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(CLK_c), 
           .D(n29978));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(CLK_c), 
           .D(n29977));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(CLK_c), 
           .D(n29976));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(CLK_c), 
           .D(n29975));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(CLK_c), 
           .D(n29974));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(CLK_c), 
           .D(n29973));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(CLK_c), 
           .D(n29972));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(CLK_c), 
           .D(n29971));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(CLK_c), 
           .D(n29970));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(CLK_c), 
           .D(n29969));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(CLK_c), 
           .D(n29968));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(CLK_c), 
           .D(n29967));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(CLK_c), 
           .D(n29966));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(CLK_c), 
           .D(n29965));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(CLK_c), 
           .D(n29964));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(CLK_c), 
           .D(n29963));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(CLK_c), 
           .D(n29962));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(CLK_c), 
           .D(n29961));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16238_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45612), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n29760));
    defparam i16238_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(CLK_c), 
           .D(n29960));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1039 (.I0(\data_out_frame[14] [4]), .I1(n46006), 
            .I2(n1519), .I3(\data_out_frame[12] [5]), .O(n12_adj_4383));
    defparam i5_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(CLK_c), 
           .D(n29959));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1040 (.I0(\data_out_frame[18] [7]), .I1(n12_adj_4383), 
            .I2(n46086), .I3(\data_out_frame[17] [0]), .O(n26083));
    defparam i6_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1041 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(n46200), .I3(n28014), .O(n18_adj_4384));
    defparam i7_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(CLK_c), 
           .D(n29958));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(CLK_c), 
           .D(n29957));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30_4_lut (.I0(n46294), .I1(\data_in_frame[12] [2]), .I2(\data_in_frame[9] [5]), 
            .I3(\data_in_frame[12] [7]), .O(n73));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1042 (.I0(\data_out_frame[5] [7]), .I1(n18_adj_4384), 
            .I2(n45899), .I3(n46350), .O(n20_adj_4385));
    defparam i9_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(CLK_c), 
           .D(n29956));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(CLK_c), 
           .D(n29955));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(CLK_c), 
           .D(n29954));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(CLK_c), 
           .D(n29953));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(CLK_c), 
           .D(n29952));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(CLK_c), 
           .D(n29951));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(CLK_c), 
           .D(n29950));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(CLK_c), 
           .D(n29949));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(CLK_c), 
           .D(n29948));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(CLK_c), 
           .D(n29947));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(CLK_c), 
           .D(n29946));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(CLK_c), 
           .D(n29945));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(CLK_c), 
           .D(n29944));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(CLK_c), 
           .D(n29943));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(CLK_c), 
           .D(n29942));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(CLK_c), 
           .D(n29941));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(CLK_c), 
           .D(n29940));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(CLK_c), 
           .D(n29939));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(CLK_c), 
           .D(n29938));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(CLK_c), 
           .D(n29937));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28_4_lut (.I0(n28264), .I1(n42817), .I2(\data_in_frame[14] [6]), 
            .I3(\data_in_frame[12] [5]), .O(n71));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(CLK_c), 
           .D(n29936));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i27_4_lut (.I0(n45893), .I1(n28676), .I2(\data_in_frame[17] [6]), 
            .I3(\data_in_frame[15] [2]), .O(n70));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(CLK_c), 
           .D(n29935));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i10_4_lut_adj_1043 (.I0(n46313), .I1(n20_adj_4385), .I2(n16_adj_4386), 
            .I3(n46000), .O(n43916));
    defparam i10_4_lut_adj_1043.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n45899));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(CLK_c), 
           .D(n29934));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1045 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n46200));
    defparam i2_3_lut_adj_1045.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(CLK_c), 
           .D(n29933));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i25_4_lut_adj_1046 (.I0(n28537), .I1(n28689), .I2(\data_in_frame[16] [1]), 
            .I3(n46380), .O(n68));
    defparam i25_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(CLK_c), 
           .D(n29932));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(CLK_c), 
           .D(n29931));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(CLK_c), 
           .D(n29930));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(CLK_c), 
           .D(n29929));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(CLK_c), 
           .D(n29928));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(CLK_c), 
           .D(n29927));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(CLK_c), 
           .D(n29926));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(CLK_c), 
           .D(n29925));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(CLK_c), 
           .D(n29924));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(CLK_c), 
           .D(n29923));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(CLK_c), 
           .D(n29922));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(CLK_c), 
           .D(n29921));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(CLK_c), 
           .D(n29920));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(CLK_c), 
           .D(n29919));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(CLK_c), 
           .D(n29918));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(CLK_c), 
           .D(n29917));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(CLK_c), 
           .D(n29916));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(CLK_c), 
           .D(n29915));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(CLK_c), 
           .D(n29914));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(CLK_c), 
           .D(n29913));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(CLK_c), 
           .D(n29912));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(CLK_c), 
           .D(n29911));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(CLK_c), 
           .D(n29910));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(CLK_c), 
           .D(n29909));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(CLK_c), 
           .D(n29908));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(CLK_c), 
           .D(n29907));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(CLK_c), 
           .D(n29906));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(CLK_c), 
           .D(n29905));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(CLK_c), 
           .D(n29904));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(CLK_c), 
           .D(n29903));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(CLK_c), 
           .D(n29902));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(CLK_c), 
           .D(n29901));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(CLK_c), 
           .D(n29900));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(CLK_c), 
           .D(n29899));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(CLK_c), 
           .D(n29898));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(CLK_c), 
           .D(n29897));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(CLK_c), 
           .D(n29896));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(CLK_c), 
           .D(n29895));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16239_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45612), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n29761));
    defparam i16239_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1047 (.I0(n45640), .I1(n45936), .I2(n1191), .I3(\data_out_frame[8] [3]), 
            .O(n12_adj_4387));
    defparam i5_4_lut_adj_1047.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(CLK_c), 
           .D(n29894));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(CLK_c), 
           .D(n29893));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(CLK_c), 
           .D(n29892));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(CLK_c), 
           .D(n29891));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16240_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45612), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n29762));
    defparam i16240_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[18] [4]), .O(n6572));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(CLK_c), 
           .D(n29890));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(CLK_c), 
           .D(n29889));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i26_4_lut (.I0(n46345), .I1(n46111), .I2(n46254), .I3(n46042), 
            .O(n69));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16241_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45612), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n29763));
    defparam i16241_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(CLK_c), 
           .D(n29888));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_1817_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[18] [5]), .O(n6573));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(CLK_c), 
           .D(n29887));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(CLK_c), 
           .D(n29886));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(CLK_c), 
           .D(n29885));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(CLK_c), 
           .D(n29884));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(CLK_c), 
           .D(n29883));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(CLK_c), 
           .D(n29882));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(CLK_c), 
           .D(n29881));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(CLK_c), 
           .D(n29880));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(CLK_c), 
           .D(n29879));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(CLK_c), 
           .D(n29878));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(CLK_c), .D(n29877));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(CLK_c), .D(n29876));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(CLK_c), .D(n29875));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(CLK_c), .D(n29874));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(CLK_c), .D(n29873));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(CLK_c), .D(n29872));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(CLK_c), .D(n29871));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(CLK_c), .D(n29870));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(CLK_c), .D(n29869));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(CLK_c), .D(n29868));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(CLK_c), .D(n29867));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(CLK_c), .D(n29866));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(CLK_c), .D(n29865));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(CLK_c), .D(n29864));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(CLK_c), .D(n29863));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(CLK_c), .D(n29862));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(CLK_c), .D(n29861));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(CLK_c), .D(n29860));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(CLK_c), .D(n29859));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(CLK_c), .D(n29858));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(CLK_c), .D(n29857));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(CLK_c), .D(n29856));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(CLK_c), .D(n29855));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1048 (.I0(n28456), .I1(n12_adj_4387), .I2(n46200), 
            .I3(\data_out_frame[12] [6]), .O(n27527));
    defparam i6_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n29847));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1049 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46307));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n29846));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n29844));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i24_4_lut_adj_1050 (.I0(n28084), .I1(n46175), .I2(n46368), 
            .I3(n45982), .O(n67));
    defparam i24_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n29843));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1051 (.I0(n46172), .I1(n46307), .I2(\data_out_frame[8] [4]), 
            .I3(GND_net), .O(n45878));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1051.LUT_INIT = 16'h9696;
    SB_LUT4 i33_4_lut (.I0(\data_in_frame[14] [5]), .I1(n66), .I2(n46322), 
            .I3(\data_in_frame[17] [5]), .O(n76));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n29842));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n29841));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1052 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n45640));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'h6666;
    SB_LUT4 i39_4_lut (.I0(n67), .I1(n69), .I2(n68), .I3(n70), .O(n82));
    defparam i39_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n29840));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i32_4_lut (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[11] [3]), .I3(\data_in_frame[12] [4]), .O(n75));
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n29839));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n29838));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i40_4_lut (.I0(n71), .I1(n73), .I2(n72), .I3(n74), .O(n83));
    defparam i40_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n46009));
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n29837));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1054 (.I0(n28651), .I1(\data_in_frame[17] [5]), 
            .I2(n46075), .I3(GND_net), .O(n43009));
    defparam i1_2_lut_3_lut_adj_1054.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1055 (.I0(n27527), .I1(\data_out_frame[14] [6]), 
            .I2(\data_out_frame[14] [7]), .I3(GND_net), .O(n46000));
    defparam i2_3_lut_adj_1055.LUT_INIT = 16'h9696;
    SB_LUT4 i42_4_lut (.I0(n83), .I1(n75), .I2(n82), .I3(n76), .O(n48418));
    defparam i42_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n29836));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1056 (.I0(n45664), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[13] [0]), .I3(n6_adj_4388), .O(n46216));
    defparam i4_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n29835));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n29834));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n29833));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n29832));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n29831));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n29830));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i10_4_lut_adj_1057 (.I0(n46039), .I1(\data_in_frame[18] [7]), 
            .I2(\data_in_frame[16] [4]), .I3(\data_in_frame[19] [1]), .O(n24_adj_4389));
    defparam i10_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1058 (.I0(n43819), .I1(n45953), .I2(\data_in_frame[18] [3]), 
            .I3(GND_net), .O(n17_adj_4390));
    defparam i3_3_lut_adj_1058.LUT_INIT = 16'h6969;
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n29829));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n29828));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i8_4_lut_adj_1059 (.I0(n42915), .I1(n46009), .I2(\data_in_frame[19] [7]), 
            .I3(n46156), .O(n22_adj_4391));
    defparam i8_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n29827));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_4_lut_adj_1060 (.I0(n17_adj_4390), .I1(n24_adj_4389), .I2(n48418), 
            .I3(n46260), .O(n26_adj_4392));
    defparam i12_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n29826));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_25_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n40480), .O(n2_adj_4292)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13_4_lut_adj_1061 (.I0(n45913), .I1(n26_adj_4392), .I2(n22_adj_4391), 
            .I3(\data_in_frame[19] [2]), .O(n46197));
    defparam i13_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n29825));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16242_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45612), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n29764));
    defparam i16242_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n53155_bdd_4_lut (.I0(n53155), .I1(n50365), .I2(n50364), .I3(byte_transmit_counter[2]), 
            .O(n53158));
    defparam n53155_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46383));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1817_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[18] [6]), .O(n6574));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16243_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45612), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n29765));
    defparam i16243_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n46111));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1064 (.I0(n46089), .I1(\data_out_frame[10] [5]), 
            .I2(n28439), .I3(n46282), .O(n10_adj_4393));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\data_in_frame[7] [0]), .I1(Kp_23__N_1217), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4271));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37751 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n53149));
    defparam byte_transmit_counter_0__bdd_4_lut_37751.LUT_INIT = 16'he4aa;
    SB_LUT4 n53149_bdd_4_lut (.I0(n53149), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n53152));
    defparam n53149_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37663 (.I0(byte_transmit_counter[1]), 
            .I1(n51337), .I2(n51338), .I3(byte_transmit_counter[2]), .O(n53143));
    defparam byte_transmit_counter_1__bdd_4_lut_37663.LUT_INIT = 16'he4aa;
    SB_LUT4 n53143_bdd_4_lut (.I0(n53143), .I1(n17_adj_4394), .I2(n16_adj_4395), 
            .I3(byte_transmit_counter[2]), .O(n53146));
    defparam n53143_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16244_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45612), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n29766));
    defparam i16244_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(CLK_c), 
           .D(n44955));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16245_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45612), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n29767));
    defparam i16245_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(CLK_c), .D(n29570));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(CLK_c), .D(n29569));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n29568));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(CLK_c), .D(n29566));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(CLK_c), .D(n29565));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(CLK_c), .D(n29564));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n29824));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), .D(n29823));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), .D(n29822));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), .D(n29821));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), .D(n29820));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), .D(n29819));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), .D(n29818));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), .D(n29817));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), .D(n29816));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(CLK_c), .D(n29815));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(CLK_c), .D(n29814));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(CLK_c), .D(n29813));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(CLK_c), .D(n29812));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(CLK_c), .D(n29811));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(CLK_c), .D(n29810));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(CLK_c), .D(n29809));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(CLK_c), .D(n29808));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), .D(n29807));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), .D(n29806));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), .D(n29805));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), .D(n29804));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), .D(n29803));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), .D(n29802));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), .D(n29801));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), .D(n29800));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n29799));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n29798));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n29797));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n29796));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n29795));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n29794));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16230_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45612), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n29752));
    defparam i16230_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(\data_in_frame[10] [6]), .I1(n28226), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4396));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1067 (.I0(n45878), .I1(n10_adj_4393), .I2(\data_out_frame[12] [7]), 
            .I3(GND_net), .O(n27529));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_adj_1067.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1068 (.I0(n45972), .I1(n27529), .I2(\data_out_frame[17] [3]), 
            .I3(n46216), .O(n10_adj_4397));
    defparam i4_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1069 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[15] [2]), 
            .I2(n10_adj_4397), .I3(\data_out_frame[13] [1]), .O(n43876));
    defparam i1_4_lut_adj_1069.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1070 (.I0(\data_out_frame[19] [2]), .I1(n43916), 
            .I2(\data_out_frame[19] [1]), .I3(n26083), .O(n42923));
    defparam i3_4_lut_adj_1070.LUT_INIT = 16'h9669;
    SB_LUT4 i16231_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45612), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n29753));
    defparam i16231_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n29793));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n29792));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(CLK_c), .D(n29791));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), .D(n29790));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), .D(n29789));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), .D(n29788));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), .D(n29787));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), .D(n29786));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), .D(n29785));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), .D(n29784));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(CLK_c), .D(n29783));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(CLK_c), .D(n29782));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(CLK_c), .D(n29781));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(CLK_c), .D(n29780));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(CLK_c), .D(n29779));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(CLK_c), .D(n29778));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(CLK_c), .D(n29777));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(CLK_c), .D(n29776));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), .D(n29775));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), .D(n29774));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), .D(n29773));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), .D(n29772));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), .D(n29771));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), .D(n29770));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(CLK_c), .D(n29769));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), .D(n29768));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n29767));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n29766));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n29765));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n29764));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n29763));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n29762));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(CLK_c), 
           .D(n29761));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n29760));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(CLK_c), 
           .D(n29759));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(CLK_c), 
           .D(n29758));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(CLK_c), 
           .D(n29757));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(CLK_c), 
           .D(n29756));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(CLK_c), 
           .D(n29755));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(CLK_c), 
           .D(n29754));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(CLK_c), 
           .D(n29753));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(CLK_c), 
           .D(n29752));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(CLK_c), 
           .D(n29751));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(CLK_c), 
           .D(n29750));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(CLK_c), 
           .D(n29749));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(CLK_c), 
           .D(n29748));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(CLK_c), 
           .D(n29747));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(CLK_c), 
           .D(n29746));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(CLK_c), 
           .D(n29745));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(CLK_c), 
           .D(n29744));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(CLK_c), 
           .D(n29743));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(CLK_c), 
           .D(n29742));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(CLK_c), 
           .D(n29741));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(CLK_c), 
           .D(n29740));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(CLK_c), 
           .D(n29739));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(CLK_c), 
           .D(n29738));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(CLK_c), 
           .D(n29737));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(CLK_c), 
           .D(n29736));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(CLK_c), 
           .D(n29735));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(CLK_c), 
           .D(n29734));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(CLK_c), 
           .D(n29733));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(CLK_c), 
           .D(n29732));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(CLK_c), 
           .D(n29731));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(CLK_c), 
           .D(n29730));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16232_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45612), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n29754));
    defparam i16232_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(n27975), .I1(\data_out_frame[11] [5]), 
            .I2(n8_adj_4398), .I3(\data_out_frame[7] [1]), .O(n42822));
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(CLK_c), 
           .D(n29729));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(CLK_c), 
           .D(n29728));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(CLK_c), 
           .D(n29727));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(CLK_c), 
           .D(n29726));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(CLK_c), 
           .D(n29725));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(CLK_c), 
           .D(n29724));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1072 (.I0(n42822), .I1(\data_out_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n46300));
    defparam i1_2_lut_adj_1072.LUT_INIT = 16'h6666;
    SB_LUT4 i1288_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2076));   // verilog/coms.v(85[17:28])
    defparam i1288_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(CLK_c), .D(n29542));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(CLK_c), .D(n29541));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(CLK_c), 
           .D(n29723));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(CLK_c), 
           .D(n29722));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(CLK_c), 
           .D(n29721));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(CLK_c), 
           .D(n29720));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(CLK_c), 
           .D(n29719));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(CLK_c), 
           .D(n29718));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(CLK_c), 
           .D(n29717));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(CLK_c), 
           .D(n29716));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n45764));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 i16233_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45612), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n29755));
    defparam i16233_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16234_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45612), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n29756));
    defparam i16234_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(CLK_c), 
           .D(n29715));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(CLK_c), 
           .D(n29714));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(CLK_c), 
           .D(n29713));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(CLK_c), 
           .D(n29712));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(CLK_c), 
           .D(n29711));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(CLK_c), 
           .D(n29710));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(CLK_c), 
           .D(n29709));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(CLK_c), 
           .D(n29708));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(CLK_c), 
           .D(n29707));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(CLK_c), 
           .D(n29706));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(CLK_c), 
           .D(n29705));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(CLK_c), 
           .D(n29704));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(CLK_c), 
           .D(n29703));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(CLK_c), 
           .D(n29702));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(CLK_c), 
           .D(n29701));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(CLK_c), 
           .D(n29700));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(CLK_c), 
           .D(n29699));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(CLK_c), 
           .D(n29698));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(CLK_c), 
           .D(n29697));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(CLK_c), 
           .D(n29696));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(CLK_c), 
           .D(n29695));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(CLK_c), 
           .D(n29694));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(CLK_c), 
           .D(n29693));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(CLK_c), 
           .D(n29692));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(CLK_c), 
           .D(n29691));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(CLK_c), 
           .D(n29690));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(CLK_c), 
           .D(n29689));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(CLK_c), 
           .D(n29688));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(CLK_c), 
           .D(n29687));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(CLK_c), 
           .D(n29686));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(CLK_c), 
           .D(n29685));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(CLK_c), 
           .D(n29684));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(CLK_c), 
           .D(n29683));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(CLK_c), 
           .D(n29682));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(CLK_c), 
           .D(n29681));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(CLK_c), 
           .D(n29680));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_25 (.CI(n40480), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n40481));
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\data_out_frame[13] [1]), .I1(n28533), 
            .I2(GND_net), .I3(GND_net), .O(n28418));
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n45704));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_24_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n40479), .O(n2_adj_4294)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_24 (.CI(n40479), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n40480));
    SB_LUT4 i4_4_lut_adj_1076 (.I0(\data_in_frame[12] [7]), .I1(n28232), 
            .I2(\data_in_frame[10] [5]), .I3(n6_adj_4396), .O(n45736));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(\data_in_frame[13] [1]), .I1(n45736), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4399));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h6666;
    SB_LUT4 i16235_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45612), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n29757));
    defparam i16235_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16236_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45612), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n29758));
    defparam i16236_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16237_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45612), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n29759));
    defparam i16237_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1078 (.I0(n28581), .I1(\data_in_frame[15] [3]), 
            .I2(\data_in_frame[13] [2]), .I3(n6_adj_4399), .O(n46075));
    defparam i4_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\data_in_frame[17] [5]), .I1(n46075), 
            .I2(GND_net), .I3(GND_net), .O(n45738));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1080 (.I0(n45758), .I1(n45821), .I2(\data_out_frame[7] [0]), 
            .I3(\data_out_frame[5] [1]), .O(n12_adj_4400));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1081 (.I0(\data_out_frame[9] [2]), .I1(n12_adj_4400), 
            .I2(n46125), .I3(\data_out_frame[4] [4]), .O(n28331));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i16222_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45612), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n29744));
    defparam i16222_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(n28331), .I1(n42820), .I2(GND_net), 
            .I3(GND_net), .O(n46133));
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1083 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28077));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1084 (.I0(\data_out_frame[17] [7]), .I1(n43839), 
            .I2(n8_adj_4401), .I3(\data_out_frame[15] [4]), .O(n46190));
    defparam i1_4_lut_adj_1084.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1085 (.I0(n28657), .I1(\data_in_frame[13] [2]), 
            .I2(n45804), .I3(n6_adj_4402), .O(n28651));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i16223_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45612), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n29745));
    defparam i16223_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28022));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n46150));
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_23_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n40478), .O(n2_adj_4296)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(71[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1088 (.I0(n1191), .I1(n45797), .I2(\data_out_frame[5] [3]), 
            .I3(GND_net), .O(n27975));
    defparam i2_3_lut_adj_1088.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1089 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(n27975), .O(n45785));   // verilog/coms.v(71[16:62])
    defparam i3_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46099));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1091 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n46122));
    defparam i2_3_lut_adj_1091.LUT_INIT = 16'h9696;
    SB_CARRY add_43_23 (.CI(n40478), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n40479));
    SB_LUT4 i16224_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45612), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n29746));
    defparam i16224_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_in_frame[9] [2]), .I1(n28544), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4403));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 i16225_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45612), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n29747));
    defparam i16225_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16226_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45612), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n29748));
    defparam i16226_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16227_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45612), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n29749));
    defparam i16227_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1093 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n45821));
    defparam i1_2_lut_adj_1093.LUT_INIT = 16'h6666;
    SB_LUT4 i16228_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45612), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n29750));
    defparam i16228_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n46103));
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1095 (.I0(\data_in_frame[11] [3]), .I1(n28537), 
            .I2(\data_in_frame[9] [1]), .I3(n6_adj_4403), .O(n28129));   // verilog/coms.v(72[16:41])
    defparam i4_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_22_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n40477), .O(n2_adj_4298)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16229_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45612), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n29751));
    defparam i16229_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1096 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n45881));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1096.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4404));
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1098 (.I0(n45788), .I1(\data_out_frame[4] [3]), 
            .I2(n46103), .I3(n6_adj_4404), .O(n42820));
    defparam i4_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1099 (.I0(\data_out_frame[4] [2]), .I1(n45881), 
            .I2(\data_out_frame[4] [5]), .I3(\data_out_frame[8] [6]), .O(n12_adj_4405));   // verilog/coms.v(76[16:27])
    defparam i5_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_CARRY add_43_22 (.CI(n40477), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n40478));
    SB_LUT4 mux_1817_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[18] [7]), .O(n6575));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1100 (.I0(\data_out_frame[6] [5]), .I1(n12_adj_4405), 
            .I2(n46163), .I3(n28447), .O(n28800));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1101 (.I0(n28232), .I1(n46234), .I2(n28544), 
            .I3(n42840), .O(n27538));
    defparam i3_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_21_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n40476), .O(n2_adj_4300)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28046));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1103 (.I0(n28800), .I1(n42820), .I2(GND_net), 
            .I3(GND_net), .O(n43839));
    defparam i1_2_lut_adj_1103.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1104 (.I0(\data_in_frame[9] [1]), .I1(n27538), 
            .I2(GND_net), .I3(GND_net), .O(n46042));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1105 (.I0(n28232), .I1(n46042), .I2(n45688), 
            .I3(\data_in_frame[9] [0]), .O(n46257));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n46175));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_CARRY add_43_21 (.CI(n40476), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n40477));
    SB_LUT4 i5_4_lut_adj_1107 (.I0(n7_adj_4406), .I1(n28771), .I2(n8_adj_4407), 
            .I3(\data_in_frame[7] [4]), .O(n28259));
    defparam i5_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n45902));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1109 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[8] [2]), 
            .I2(\data_in_frame[8] [6]), .I3(\data_in_frame[8] [1]), .O(n29001));
    defparam i3_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46172));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1111 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4408));   // verilog/coms.v(78[16:27])
    defparam i2_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1112 (.I0(\data_out_frame[4] [1]), .I1(n46172), 
            .I2(n45902), .I3(\data_out_frame[8] [7]), .O(n45779));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1113 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [5]), .O(n44965));
    defparam i1_2_lut_4_lut_adj_1113.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n46125));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1115 (.I0(n45779), .I1(n45887), .I2(\data_out_frame[13] [3]), 
            .I3(\data_out_frame[11] [1]), .O(n12_adj_4411));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1116 (.I0(n29014), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[4] [4]), .I3(n28213), .O(n14_adj_4412));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1117 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [6]), .O(n45019));
    defparam i1_2_lut_4_lut_adj_1117.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1118 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [7]), .O(n44975));
    defparam i1_2_lut_4_lut_adj_1118.LUT_INIT = 16'hba00;
    SB_LUT4 i6_4_lut_adj_1119 (.I0(\data_out_frame[10] [7]), .I1(n12_adj_4411), 
            .I2(n46163), .I3(\data_out_frame[9] [1]), .O(n28533));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1817_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[17] [0]), .O(n6576));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_out_frame[17] [6]), .I1(n43923), 
            .I2(GND_net), .I3(GND_net), .O(n46053));
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1121 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46313));
    defparam i1_2_lut_adj_1121.LUT_INIT = 16'h6666;
    SB_LUT4 i22_4_lut (.I0(n46053), .I1(\data_out_frame[17] [5]), .I2(n28533), 
            .I3(n46125), .O(n60));   // verilog/coms.v(85[17:28])
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1122 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [9]), .O(n44977));
    defparam i1_2_lut_4_lut_adj_1122.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_3_lut_adj_1123 (.I0(n63_c), .I1(n63_adj_4213), .I2(n63), 
            .I3(GND_net), .O(n25059));   // verilog/coms.v(139[7:80])
    defparam i1_2_lut_3_lut_adj_1123.LUT_INIT = 16'h8080;
    SB_LUT4 add_43_20_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n40475), .O(n2_adj_4302)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n40475), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n40476));
    SB_LUT4 i1_2_lut_4_lut_adj_1124 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [11]), .O(n45017));
    defparam i1_2_lut_4_lut_adj_1124.LUT_INIT = 16'hba00;
    SB_LUT4 i20_4_lut_adj_1125 (.I0(n46150), .I1(n28022), .I2(\data_out_frame[17] [2]), 
            .I3(n46190), .O(n58));   // verilog/coms.v(85[17:28])
    defparam i20_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut_adj_1126 (.I0(n45990), .I1(n60), .I2(n42_adj_4413), 
            .I3(\data_out_frame[17] [4]), .O(n68_adj_4414));   // verilog/coms.v(85[17:28])
    defparam i30_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut_adj_1127 (.I0(n45704), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[8] [1]), .I3(n28418), .O(n66_adj_4415));   // verilog/coms.v(85[17:28])
    defparam i28_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i29_3_lut (.I0(\data_out_frame[16] [3]), .I1(n58), .I2(\data_out_frame[8] [2]), 
            .I3(GND_net), .O(n67_adj_4416));   // verilog/coms.v(85[17:28])
    defparam i29_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i27_4_lut_adj_1128 (.I0(n45972), .I1(n45764), .I2(n45939), 
            .I3(n45710), .O(n65));   // verilog/coms.v(85[17:28])
    defparam i27_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1129 (.I0(n45990), .I1(n42923), .I2(n43876), 
            .I3(\data_out_frame[18] [1]), .O(n24_adj_4417));
    defparam i10_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1130 (.I0(\data_out_frame[11] [2]), .I1(n46307), 
            .I2(\data_out_frame[14] [7]), .I3(n46003), .O(n62));   // verilog/coms.v(85[17:28])
    defparam i24_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1131 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [15]), .O(n44979));
    defparam i1_2_lut_4_lut_adj_1131.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1132 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [23]), .O(n44973));
    defparam i1_2_lut_4_lut_adj_1132.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1133 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [25]), .O(n44925));
    defparam i1_2_lut_4_lut_adj_1133.LUT_INIT = 16'hba00;
    SB_LUT4 i26_4_lut_adj_1134 (.I0(\data_out_frame[13] [4]), .I1(n46159), 
            .I2(n46350), .I3(n46006), .O(n64));   // verilog/coms.v(85[17:28])
    defparam i26_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1135 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [26]), .O(n44947));
    defparam i1_2_lut_4_lut_adj_1135.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1136 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [27]), .O(n45015));
    defparam i1_2_lut_4_lut_adj_1136.LUT_INIT = 16'hba00;
    SB_LUT4 i25_4_lut_adj_1137 (.I0(n45788), .I1(\data_out_frame[10] [7]), 
            .I2(n45707), .I3(n28486), .O(n63_adj_4418));   // verilog/coms.v(85[17:28])
    defparam i25_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_19_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n40474), .O(n2_adj_4304)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i36_4_lut (.I0(n65), .I1(n67_adj_4416), .I2(n66_adj_4415), 
            .I3(n68_adj_4414), .O(n74_adj_4419));   // verilog/coms.v(85[17:28])
    defparam i36_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1817_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[17] [1]), .O(n6577));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7_4_lut_adj_1138 (.I0(\data_in_frame[2] [1]), .I1(n14_adj_4412), 
            .I2(n10_adj_4408), .I3(\data_in_frame[0] [2]), .O(Kp_23__N_1195));   // verilog/coms.v(78[16:27])
    defparam i7_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n45773));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_LUT4 i31_4_lut_adj_1140 (.I0(n45_adj_4420), .I1(n62), .I2(n46371), 
            .I3(n45942), .O(n69_adj_4421));   // verilog/coms.v(85[17:28])
    defparam i31_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1141 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [28]), .O(n45013));
    defparam i1_2_lut_4_lut_adj_1141.LUT_INIT = 16'hba00;
    SB_LUT4 i8_4_lut_adj_1142 (.I0(n46133), .I1(n45916), .I2(\data_out_frame[18] [0]), 
            .I3(n43235), .O(n22_adj_4422));
    defparam i8_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n46092));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1144 (.I0(\data_in_frame[0] [4]), .I1(n46092), 
            .I2(n45773), .I3(\data_in_frame[0] [3]), .O(n28992));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1145 (.I0(n45979), .I1(n24_adj_4417), .I2(n18_adj_4423), 
            .I3(n45697), .O(n26_adj_4424));
    defparam i12_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1146 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [1]), .O(n28771));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1147 (.I0(\data_in_frame[5] [4]), .I1(n28771), 
            .I2(GND_net), .I3(GND_net), .O(n45648));
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_LUT4 i37_4_lut (.I0(n69_adj_4421), .I1(n74_adj_4419), .I2(n63_adj_4418), 
            .I3(n64), .O(n48223));   // verilog/coms.v(85[17:28])
    defparam i37_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1148 (.I0(n48223), .I1(n26_adj_4424), .I2(n22_adj_4422), 
            .I3(\data_out_frame[18] [5]), .O(n42875));
    defparam i13_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1149 (.I0(\data_in_frame[5] [2]), .I1(n46291), 
            .I2(GND_net), .I3(GND_net), .O(n45791));
    defparam i1_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1150 (.I0(Kp_23__N_1020), .I1(n46119), .I2(n45791), 
            .I3(n28857), .O(n28_adj_4425));   // verilog/coms.v(70[16:69])
    defparam i10_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1151 (.I0(n7_adj_4409), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n9_adj_4410), .I3(\FRAME_MATCHER.state [31]), .O(n45011));
    defparam i1_2_lut_4_lut_adj_1151.LUT_INIT = 16'hba00;
    SB_LUT4 i14_3_lut_adj_1152 (.I0(\data_in_frame[5] [3]), .I1(n28_adj_4425), 
            .I2(\data_in_frame[4] [7]), .I3(GND_net), .O(n32_adj_4426));   // verilog/coms.v(70[16:69])
    defparam i14_3_lut_adj_1152.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1153 (.I0(n28120), .I1(n46067), .I2(n46297), 
            .I3(n45794), .O(n30_adj_4427));   // verilog/coms.v(70[16:69])
    defparam i12_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_CARRY add_43_19 (.CI(n40474), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n40475));
    SB_LUT4 i11_4_lut_adj_1154 (.I0(n29005), .I1(n45679), .I2(n46027), 
            .I3(\data_in_frame[3] [5]), .O(n29_adj_4428));   // verilog/coms.v(70[16:69])
    defparam i11_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1817_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[17] [2]), .O(n6578));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17_4_lut_adj_1155 (.I0(n29_adj_4428), .I1(n31_adj_4429), .I2(n30_adj_4427), 
            .I3(n32_adj_4426), .O(n43663));   // verilog/coms.v(70[16:69])
    defparam i17_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_18_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n40473), .O(n2_adj_4306)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1156 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n45936));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1156.LUT_INIT = 16'h6666;
    SB_CARRY add_43_18 (.CI(n40473), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n40474));
    SB_LUT4 i1_2_lut_adj_1157 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28213));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1158 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28645));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1159 (.I0(n28645), .I1(n28213), .I2(\data_in_frame[6] [6]), 
            .I3(GND_net), .O(n45726));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1159.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37658 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n53137));
    defparam byte_transmit_counter_0__bdd_4_lut_37658.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1160 (.I0(\data_in_frame[6] [0]), .I1(n43663), 
            .I2(n6_adj_4430), .I3(\data_in_frame[6] [2]), .O(n11_adj_4364));   // verilog/coms.v(85[17:63])
    defparam i1_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_17_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n40472), .O(n2_adj_4308)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_17 (.CI(n40472), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n40473));
    SB_LUT4 i1_2_lut_3_lut_adj_1161 (.I0(n63_c), .I1(n63_adj_4213), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n123));   // verilog/coms.v(139[7:80])
    defparam i1_2_lut_3_lut_adj_1161.LUT_INIT = 16'h8080;
    SB_LUT4 mux_1817_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[17] [3]), .O(n6579));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i21806_2_lut_3_lut (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n35309));
    defparam i21806_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1162 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28035));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1162.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_16_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n40471), .O(n2_adj_4310)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_16 (.CI(n40471), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n40472));
    SB_LUT4 i1_2_lut_3_lut_adj_1163 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n45061));
    defparam i1_2_lut_3_lut_adj_1163.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1164 (.I0(n28035), .I1(n46285), .I2(n45782), 
            .I3(\data_out_frame[7] [7]), .O(n1516));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1165 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n45065));
    defparam i1_2_lut_3_lut_adj_1165.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_15_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n40470), .O(n2_adj_4312)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1166 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n45926));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1166.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1167 (.I0(n45926), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[10] [2]), .I3(n46059), .O(n10_adj_4433));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1168 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n45069));
    defparam i1_2_lut_3_lut_adj_1168.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_3_lut_adj_1169 (.I0(\data_out_frame[10] [1]), .I1(n10_adj_4433), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n1513));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1170 (.I0(n28299), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4434));   // verilog/coms.v(75[16:27])
    defparam i2_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1171 (.I0(n4_adj_4435), .I1(\data_in_frame[5] [6]), 
            .I2(n8_adj_4434), .I3(n46014), .O(n45969));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n45758));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1173 (.I0(n28219), .I1(n45969), .I2(GND_net), 
            .I3(GND_net), .O(n45971));
    defparam i1_2_lut_adj_1173.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n45797));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1175 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n46342));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1175.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1176 (.I0(Kp_23__N_1183), .I1(\data_in_frame[7] [0]), 
            .I2(Kp_23__N_1195), .I3(n29001), .O(n10_adj_4436));
    defparam i4_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_CARRY add_43_15 (.CI(n40470), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n40471));
    SB_LUT4 n53137_bdd_4_lut (.I0(n53137), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n53140));
    defparam n53137_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_43_14_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n40469), .O(n2_adj_4314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1177 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n7_adj_4264));
    defparam i1_2_lut_3_lut_adj_1177.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_1178 (.I0(\data_out_frame[14] [2]), .I1(n46056), 
            .I2(\data_out_frame[12] [1]), .I3(n46342), .O(n16_adj_4437));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_adj_1179 (.I0(n28226), .I1(Kp_23__N_1214), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4438));
    defparam i3_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1180 (.I0(n46049), .I1(Kp_23__N_1237), .I2(n9_adj_4438), 
            .I3(n10_adj_4436), .O(n45993));
    defparam i2_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1181 (.I0(\data_in_frame[7] [6]), .I1(n28299), 
            .I2(n28120), .I3(GND_net), .O(n28264));
    defparam i2_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1182 (.I0(n28264), .I1(n45993), .I2(n45971), 
            .I3(n28657), .O(n46234));
    defparam i3_4_lut_adj_1182.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1183 (.I0(\data_out_frame[9] [5]), .I1(n46266), 
            .I2(\data_out_frame[9] [6]), .I3(n45797), .O(n17_adj_4439));   // verilog/coms.v(85[17:28])
    defparam i7_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1184 (.I0(n17_adj_4439), .I1(\data_out_frame[10] [0]), 
            .I2(n16_adj_4437), .I3(\data_out_frame[12] [0]), .O(n42805));   // verilog/coms.v(85[17:28])
    defparam i9_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1185 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n45073));
    defparam i1_2_lut_3_lut_adj_1185.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(\data_out_frame[16] [4]), .I1(n42805), 
            .I2(GND_net), .I3(GND_net), .O(n46003));
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_out_frame[16] [6]), .I1(n45807), 
            .I2(GND_net), .I3(GND_net), .O(n28176));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1817_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[17] [4]), .O(n6580));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n45801));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4440));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1190 (.I0(n45719), .I1(n45644), .I2(n46234), 
            .I3(n6_adj_4440), .O(n46331));
    defparam i4_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1191 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46095));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1191.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1192 (.I0(n45923), .I1(\data_in_frame[8] [0]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n46116));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1192.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1193 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n45939));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1194 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46288));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1194.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1195 (.I0(\data_in_frame[3] [6]), .I1(n46116), 
            .I2(n45811), .I3(\data_in_frame[6] [0]), .O(n28219));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1196 (.I0(n45939), .I1(n46095), .I2(\data_out_frame[7] [4]), 
            .I3(\data_out_frame[10] [0]), .O(n12_adj_4441));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1197 (.I0(\data_in_frame[5] [5]), .I1(n46237), 
            .I2(GND_net), .I3(GND_net), .O(n45713));
    defparam i1_2_lut_adj_1197.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1198 (.I0(\data_out_frame[10] [1]), .I1(n12_adj_4441), 
            .I2(n46288), .I3(\data_out_frame[5] [2]), .O(n1510));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i21807_2_lut_3_lut (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n35311));
    defparam i21807_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1199 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n45077));
    defparam i1_2_lut_3_lut_adj_1199.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1200 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n46269));
    defparam i1_2_lut_adj_1200.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1201 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n45661));
    defparam i2_3_lut_adj_1201.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1202 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[3] [6]), .I3(GND_net), .O(n45679));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_adj_1202.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n46266));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1204 (.I0(n45652), .I1(\data_in_frame[10] [1]), 
            .I2(n45679), .I3(n6_adj_4442), .O(n46359));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_in_frame[9] [7]), .I1(n46359), 
            .I2(GND_net), .I3(GND_net), .O(n46310));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i21808_2_lut_3_lut (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n35313));
    defparam i21808_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_4_lut_adj_1206 (.I0(n45661), .I1(n45713), .I2(\data_in_frame[10] [3]), 
            .I3(\data_in_frame[8] [2]), .O(n12_adj_4443));
    defparam i5_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1207 (.I0(\data_in_frame[7] [7]), .I1(n12_adj_4443), 
            .I2(n45845), .I3(\data_in_frame[5] [7]), .O(n28287));
    defparam i6_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1208 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n7_adj_4262));
    defparam i1_2_lut_3_lut_adj_1208.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28414));
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1210 (.I0(\data_in_frame[5] [4]), .I1(n28414), 
            .I2(n26983), .I3(\data_in_frame[7] [5]), .O(n45815));
    defparam i3_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(n29005), .I1(n45815), .I2(GND_net), 
            .I3(GND_net), .O(n28368));
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1212 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n7_adj_4260));
    defparam i1_2_lut_3_lut_adj_1212.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1213 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[12] [4]), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n45905));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_CARRY add_43_14 (.CI(n40469), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n40470));
    SB_LUT4 i4_4_lut_adj_1214 (.I0(n46331), .I1(n45801), .I2(\data_in_frame[14] [3]), 
            .I3(n46359), .O(n10_adj_4444));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1215 (.I0(n46257), .I1(n10_adj_4444), .I2(\data_in_frame[12] [2]), 
            .I3(GND_net), .O(n28275));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_adj_1215.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1216 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n45081));
    defparam i1_2_lut_3_lut_adj_1216.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4445));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n45710));
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(CLK_c), 
           .D(n29679));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1219 (.I0(n45710), .I1(n46059), .I2(\data_out_frame[11] [7]), 
            .I3(\data_out_frame[5] [1]), .O(n12_adj_4446));
    defparam i5_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1220 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n7_adj_4258));
    defparam i1_2_lut_3_lut_adj_1220.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_13_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n40468), .O(n2_adj_4316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i21809_2_lut_3_lut (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n35315));
    defparam i21809_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_1221 (.I0(\data_out_frame[10] [0]), .I1(n12_adj_4446), 
            .I2(n46269), .I3(\data_out_frame[7] [3]), .O(n27502));
    defparam i6_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\data_out_frame[12] [1]), .I1(n27502), 
            .I2(GND_net), .I3(GND_net), .O(n46086));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1817_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[17] [5]), .O(n6581));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1223 (.I0(n28146), .I1(n28275), .I2(n45905), 
            .I3(n6_adj_4445), .O(n45933));   // verilog/coms.v(76[16:43])
    defparam i4_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1224 (.I0(\data_in_frame[16] [7]), .I1(n46310), 
            .I2(n46175), .I3(n45905), .O(n14_adj_4447));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1225 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n35317));
    defparam i1_2_lut_3_lut_adj_1225.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1226 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n7_adj_4256));
    defparam i1_2_lut_3_lut_adj_1226.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1227 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n7_adj_4254));
    defparam i1_2_lut_3_lut_adj_1227.LUT_INIT = 16'he0e0;
    SB_LUT4 i7_4_lut_adj_1228 (.I0(\data_in_frame[14] [7]), .I1(n14_adj_4447), 
            .I2(n10_adj_4448), .I3(n45722), .O(n28540));   // verilog/coms.v(76[16:43])
    defparam i7_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1817_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[17] [6]), .O(n6582));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1229 (.I0(n45807), .I1(\data_out_frame[16] [5]), 
            .I2(n42799), .I3(GND_net), .O(n46136));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1229.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1230 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n7_adj_4252));
    defparam i1_2_lut_3_lut_adj_1230.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1231 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[14] [5]), 
            .I2(n28176), .I3(n28584), .O(n10_adj_4449));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_CARRY add_43_13 (.CI(n40468), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n40469));
    SB_LUT4 i4_4_lut_adj_1232 (.I0(n45833), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[18] [5]), .I3(n46136), .O(n10_adj_4450));
    defparam i4_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1233 (.I0(n42795), .I1(n10_adj_4450), .I2(n42875), 
            .I3(GND_net), .O(n27578));
    defparam i5_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1234 (.I0(n42875), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42909));
    defparam i1_2_lut_adj_1234.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1235 (.I0(n42923), .I1(\data_out_frame[23] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n45848));
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_0__3__I_0_2_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_979));   // verilog/coms.v(74[16:27])
    defparam data_in_frame_0__3__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1236 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [7]), .I3(GND_net), .O(n46356));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1236.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1237 (.I0(\data_out_frame[23] [5]), .I1(\data_out_frame[23] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28149));
    defparam i1_2_lut_adj_1237.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1238 (.I0(n42913), .I1(n45859), .I2(GND_net), 
            .I3(GND_net), .O(n45860));
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1239 (.I0(\data_out_frame[25] [5]), .I1(n45860), 
            .I2(n28149), .I3(n43943), .O(n45956));
    defparam i3_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1240 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n7_adj_4250));
    defparam i1_2_lut_3_lut_adj_1240.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1241 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n45085));
    defparam i1_2_lut_3_lut_adj_1241.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1242 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n45652));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1243 (.I0(\data_out_frame[25] [6]), .I1(n45956), 
            .I2(GND_net), .I3(GND_net), .O(n45957));
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_988), 
            .I2(GND_net), .I3(GND_net), .O(n45694));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_in_frame[7] [3]), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4451));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1246 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n7_adj_4248));
    defparam i1_2_lut_3_lut_adj_1246.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1247 (.I0(Kp_23__N_988), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[0] [7]), .I3(n6_adj_4451), .O(n45818));
    defparam i4_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\data_in_frame[5] [2]), .I1(n28937), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4452));
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1249 (.I0(n45818), .I1(n26983), .I2(n28673), 
            .I3(n6_adj_4452), .O(n42840));
    defparam i4_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(\data_in_frame[7] [1]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4453));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h6666;
    SB_LUT4 i21811_2_lut_3_lut (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n35319));
    defparam i21811_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1251 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[4] [5]), .I3(n6_adj_4453), .O(n45836));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_in_frame[0] [1]), .I1(n45656), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1020));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i21812_2_lut_3_lut (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n35321));
    defparam i21812_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1253 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n45089));
    defparam i1_2_lut_3_lut_adj_1253.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1254 (.I0(Kp_23__N_1020), .I1(n45836), .I2(\data_in_frame[6] [7]), 
            .I3(n28673), .O(n28544));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1255 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n45093));
    defparam i1_2_lut_3_lut_adj_1255.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37649 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n53131));
    defparam byte_transmit_counter_0__bdd_4_lut_37649.LUT_INIT = 16'he4aa;
    SB_LUT4 i21814_2_lut_3_lut (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n35325));
    defparam i21814_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1817_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[17] [7]), .O(n6583));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1256 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n7_adj_4246));
    defparam i1_2_lut_3_lut_adj_1256.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1257 (.I0(n49), .I1(n2_adj_4432), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n45097));
    defparam i1_2_lut_3_lut_adj_1257.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1817_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35344), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[19] [0]), .O(n6560));   // verilog/coms.v(127[12] 300[6])
    defparam mux_1817_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1258 (.I0(n46067), .I1(\data_in_frame[4] [6]), 
            .I2(Kp_23__N_977), .I3(\data_in_frame[6] [7]), .O(n14_adj_4454));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1259 (.I0(\data_in_frame[0] [4]), .I1(n14_adj_4454), 
            .I2(n10_adj_4455), .I3(\data_in_frame[0] [2]), .O(Kp_23__N_1217));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1260 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n4_adj_4357));   // verilog/coms.v(70[16:27])
    defparam i1_3_lut_adj_1260.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_0__5__I_0_2_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_981));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_0__5__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1261 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n28937));
    defparam i1_3_lut_adj_1261.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n45794));
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(\data_in_frame[11] [4]), .I1(Kp_23__N_1217), 
            .I2(GND_net), .I3(GND_net), .O(n46368));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1264 (.I0(Kp_23__N_979), .I1(n12_adj_4456), .I2(n46291), 
            .I3(\data_in_frame[2] [4]), .O(Kp_23__N_1237));
    defparam i6_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(\data_in_frame[9] [4]), .I1(n28544), 
            .I2(GND_net), .I3(GND_net), .O(n46036));
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 select_622_Select_1_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4327));
    defparam select_622_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_2_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4326));
    defparam select_622_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n45729));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n29014));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1268 (.I0(\data_in_frame[6] [4]), .I1(n46297), 
            .I2(\data_in_frame[4] [1]), .I3(GND_net), .O(n46024));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_adj_1268.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_0__1__I_0_2_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_977));   // verilog/coms.v(72[16:27])
    defparam data_in_frame_0__1__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n46386));
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1270 (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n45671), .I3(n6_adj_4457), .O(n28232));   // verilog/coms.v(70[16:69])
    defparam i4_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 select_622_Select_3_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4325));
    defparam select_622_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_4_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4324));
    defparam select_622_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i5_4_lut_adj_1271 (.I0(\data_in_frame[1] [7]), .I1(n45656), 
            .I2(\data_in_frame[4] [3]), .I3(\data_in_frame[4] [5]), .O(n12_adj_4458));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 select_622_Select_5_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4323));
    defparam select_622_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 n53131_bdd_4_lut (.I0(n53131), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n53134));
    defparam n53131_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1272 (.I0(\data_in_frame[2] [1]), .I1(n12_adj_4458), 
            .I2(n45729), .I3(\data_in_frame[6] [5]), .O(Kp_23__N_1214));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 select_622_Select_6_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4322));
    defparam select_622_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1273 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_1214), 
            .I2(GND_net), .I3(GND_net), .O(n28537));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1273.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1274 (.I0(\data_in_frame[9] [0]), .I1(n45716), 
            .I2(n28537), .I3(GND_net), .O(n28581));
    defparam i2_3_lut_adj_1274.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1275 (.I0(\data_in_frame[15] [5]), .I1(n28581), 
            .I2(\data_in_frame[13] [3]), .I3(GND_net), .O(n45975));
    defparam i2_3_lut_adj_1275.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1276 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46365));
    defparam i1_2_lut_adj_1276.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1277 (.I0(n43591), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46322));
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'h6666;
    SB_LUT4 select_622_Select_7_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4321));
    defparam select_622_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_4_lut_adj_1278 (.I0(n27974), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state_31__N_2724 [3]), .I3(n47441), .O(n44983));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_1278.LUT_INIT = 16'hdc50;
    SB_LUT4 i3_4_lut_adj_1279 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[5] [6]), .O(n45845));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1280 (.I0(\FRAME_MATCHER.state [4]), .I1(n34776), 
            .I2(GND_net), .I3(GND_net), .O(n44963));
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1281 (.I0(n4_adj_4435), .I1(n45845), .I2(n8_adj_4459), 
            .I3(\data_in_frame[6] [1]), .O(Kp_23__N_1183));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 equal_2054_i3_2_lut (.I0(Kp_23__N_1183), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4267));   // verilog/coms.v(236[9:81])
    defparam equal_2054_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1282 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4435));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1282.LUT_INIT = 16'h6666;
    SB_LUT4 select_622_Select_8_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4320));
    defparam select_622_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1283 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28857));
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n45667));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1285 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n46119));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h6666;
    SB_LUT4 select_622_Select_9_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4319));
    defparam select_622_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1286 (.I0(n34776), .I1(\FRAME_MATCHER.state [8]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4265));
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n46027));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46128));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1289 (.I0(n46119), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[6] [1]), .I3(n46247), .O(n10_adj_4460));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1289.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1290 (.I0(n45811), .I1(n10_adj_4460), .I2(\data_in_frame[8] [3]), 
            .I3(GND_net), .O(n28226));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1291 (.I0(n45671), .I1(n46247), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4461));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h6666;
    SB_LUT4 select_622_Select_10_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4318));
    defparam select_622_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i4_4_lut_adj_1292 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n46027), .I3(n6_adj_4461), .O(n28657));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(n28226), .I1(n45825), .I2(GND_net), 
            .I3(GND_net), .O(n28676));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1294 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n46181));
    defparam i1_2_lut_adj_1294.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1295 (.I0(n46075), .I1(n28902), .I2(\data_in_frame[17] [4]), 
            .I3(GND_net), .O(n42817));
    defparam i2_3_lut_adj_1295.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1296 (.I0(n42817), .I1(n46181), .I2(\data_in_frame[19] [5]), 
            .I3(n28881), .O(n16_adj_4462));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1297 (.I0(n46219), .I1(n46322), .I2(n46365), 
            .I3(GND_net), .O(n8_adj_4463));
    defparam i3_3_lut_adj_1297.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1298 (.I0(\data_in_frame[21] [3]), .I1(n28540), 
            .I2(n45933), .I3(GND_net), .O(n8_adj_4464));   // verilog/coms.v(72[16:41])
    defparam i3_3_lut_adj_1298.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1299 (.I0(\data_in_frame[16] [6]), .I1(n46197), 
            .I2(n45933), .I3(\data_in_frame[21] [1]), .O(n47492));
    defparam i3_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1300 (.I0(n34776), .I1(\FRAME_MATCHER.state [13]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4263));
    defparam i1_2_lut_adj_1300.LUT_INIT = 16'h8888;
    SB_LUT4 select_622_Select_11_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4317));
    defparam select_622_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i6_4_lut_adj_1301 (.I0(n46319), .I1(n28129), .I2(\data_in_frame[19] [7]), 
            .I3(n42817), .O(n14_adj_4465));
    defparam i6_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1302 (.I0(n46254), .I1(\data_in_frame[20] [1]), 
            .I2(\data_in_frame[13] [3]), .I3(n28129), .O(n14_adj_4466));
    defparam i6_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1303 (.I0(\data_in_frame[20] [0]), .I1(n46219), 
            .I2(\data_in_frame[13] [4]), .I3(n45738), .O(n13_adj_4467));
    defparam i5_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1304 (.I0(n34776), .I1(\FRAME_MATCHER.state [14]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4261));
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1305 (.I0(n46338), .I1(n46039), .I2(n28581), 
            .I3(\data_in_frame[19] [7]), .O(n13_adj_4468));
    defparam i5_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1306 (.I0(\data_in_frame[21] [2]), .I1(\data_in_frame[14] [6]), 
            .I2(n45950), .I3(GND_net), .O(n14_adj_4469));
    defparam i5_3_lut_adj_1306.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1307 (.I0(n46277), .I1(\data_in_frame[18] [6]), 
            .I2(n42881), .I3(n46077), .O(n15_adj_4470));
    defparam i6_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1308 (.I0(n46260), .I1(n45975), .I2(\data_in_frame[20] [3]), 
            .I3(n46338), .O(n10_adj_4471));
    defparam i4_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1309 (.I0(n15_adj_4470), .I1(n45896), .I2(n14_adj_4469), 
            .I3(\data_in_frame[19] [0]), .O(n48007));
    defparam i8_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1310 (.I0(n28140), .I1(\data_in_frame[18] [2]), 
            .I2(n8_adj_4472), .I3(n45982), .O(n6_adj_4473));
    defparam i2_4_lut_adj_1310.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_adj_1311 (.I0(\data_in_frame[21] [7]), .I1(\data_in_frame[19] [5]), 
            .I2(n28084), .I3(n46319), .O(n47431));
    defparam i2_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut (.I0(\data_in_frame[19] [4]), .I1(n16_adj_4462), .I2(\data_in_frame[14] [6]), 
            .I3(GND_net), .O(n18_adj_4474));   // verilog/coms.v(78[16:27])
    defparam i8_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1312 (.I0(n46272), .I1(n28881), .I2(\data_in_frame[19] [3]), 
            .I3(\data_in_frame[19] [2]), .O(n14_adj_4475));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1313 (.I0(\data_in_frame[21] [6]), .I1(\data_in_frame[14] [7]), 
            .I2(n45910), .I3(n42881), .O(n17_adj_4476));   // verilog/coms.v(78[16:27])
    defparam i7_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1314 (.I0(\data_in_frame[21] [4]), .I1(n46072), 
            .I2(\data_in_frame[15] [1]), .I3(n28279), .O(n13_adj_4477));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1315 (.I0(n46046), .I1(n46225), .I2(\data_in_frame[18] [4]), 
            .I3(\data_in_frame[13] [5]), .O(n12_adj_4478));
    defparam i5_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1316 (.I0(\data_in_frame[20] [5]), .I1(n43819), 
            .I2(\data_in_frame[16] [3]), .I3(\data_in_frame[18] [3]), .O(n11_adj_4479));
    defparam i4_4_lut_adj_1316.LUT_INIT = 16'h9669;
    SB_LUT4 i79_2_lut (.I0(n34776), .I1(\FRAME_MATCHER.state [16]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4259));
    defparam i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_622_Select_12_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4315));
    defparam select_622_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i8_4_lut_adj_1317 (.I0(n13_adj_4477), .I1(n17_adj_4476), .I2(n14_adj_4475), 
            .I3(n18_adj_4474), .O(n24_adj_4480));
    defparam i8_4_lut_adj_1317.LUT_INIT = 16'h7bde;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37644 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n53125));
    defparam byte_transmit_counter_0__bdd_4_lut_37644.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1318 (.I0(\data_in_frame[21] [5]), .I1(n46009), 
            .I2(n28540), .I3(n28084), .O(n48304));
    defparam i3_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1319 (.I0(n34776), .I1(\FRAME_MATCHER.state [19]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4257));
    defparam i1_2_lut_adj_1319.LUT_INIT = 16'h8888;
    SB_LUT4 i3_3_lut_adj_1320 (.I0(\data_in_frame[18] [5]), .I1(n28275), 
            .I2(n46153), .I3(GND_net), .O(n8_adj_4481));
    defparam i3_3_lut_adj_1320.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1321 (.I0(n34776), .I1(\FRAME_MATCHER.state [20]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4255));
    defparam i1_2_lut_adj_1321.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1322 (.I0(n46263), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[16] [3]), .I3(n43819), .O(n14_adj_4482));
    defparam i6_4_lut_adj_1322.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1323 (.I0(\data_in_frame[20] [7]), .I1(\data_in_frame[19] [0]), 
            .I2(n46197), .I3(GND_net), .O(n7_adj_4483));
    defparam i2_3_lut_adj_1323.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1324 (.I0(n34776), .I1(\FRAME_MATCHER.state [21]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4253));
    defparam i1_2_lut_adj_1324.LUT_INIT = 16'h8888;
    SB_LUT4 select_622_Select_13_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4313));
    defparam select_622_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i5_4_lut_adj_1325 (.I0(\data_in_frame[20] [6]), .I1(n46153), 
            .I2(n45953), .I3(\data_in_frame[16] [2]), .O(n13_adj_4484));
    defparam i5_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1326 (.I0(n28651), .I1(\data_in_frame[18] [0]), 
            .I2(n8_adj_4463), .I3(n46338), .O(n6_adj_4485));
    defparam i2_4_lut_adj_1326.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_adj_1327 (.I0(\data_in_frame[19] [0]), .I1(n46156), 
            .I2(n46197), .I3(\data_in_frame[21] [0]), .O(n47374));
    defparam i2_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1328 (.I0(\data_in_frame[19] [2]), .I1(n47492), 
            .I2(n8_adj_4464), .I3(n45896), .O(n20_adj_4486));
    defparam i4_4_lut_adj_1328.LUT_INIT = 16'hdeed;
    SB_LUT4 i2_4_lut_adj_1329 (.I0(n13_adj_4468), .I1(n13_adj_4467), .I2(n14_adj_4466), 
            .I3(n14_adj_4465), .O(n18_adj_4487));
    defparam i2_4_lut_adj_1329.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1330 (.I0(n46046), .I1(n48007), .I2(n10_adj_4471), 
            .I3(\data_in_frame[17] [7]), .O(n19_adj_4488));
    defparam i3_4_lut_adj_1330.LUT_INIT = 16'hedde;
    SB_LUT4 i1_4_lut_adj_1331 (.I0(n47374), .I1(\data_in_frame[18] [1]), 
            .I2(n6_adj_4485), .I3(\data_in_frame[20] [2]), .O(n17_adj_4489));
    defparam i1_4_lut_adj_1331.LUT_INIT = 16'hd77d;
    SB_LUT4 i34659_4_lut (.I0(n47431), .I1(\data_in_frame[18] [3]), .I2(n6_adj_4473), 
            .I3(\data_in_frame[20] [4]), .O(n50031));
    defparam i34659_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12_4_lut_adj_1332 (.I0(n48304), .I1(n24_adj_4480), .I2(n11_adj_4479), 
            .I3(n12_adj_4478), .O(n28_adj_4490));
    defparam i12_4_lut_adj_1332.LUT_INIT = 16'hfeef;
    SB_LUT4 i1_2_lut_adj_1333 (.I0(n34776), .I1(\FRAME_MATCHER.state [22]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4251));
    defparam i1_2_lut_adj_1333.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1334 (.I0(n13_adj_4484), .I1(n7_adj_4483), .I2(n14_adj_4482), 
            .I3(n8_adj_4481), .O(n21_adj_4491));
    defparam i5_4_lut_adj_1334.LUT_INIT = 16'h7bde;
    SB_LUT4 i13_4_lut_adj_1335 (.I0(n17_adj_4489), .I1(n19_adj_4488), .I2(n18_adj_4487), 
            .I3(n20_adj_4486), .O(n29_adj_4492));
    defparam i13_4_lut_adj_1335.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1336 (.I0(n29_adj_4492), .I1(n21_adj_4491), .I2(n28_adj_4490), 
            .I3(n50031), .O(n31_adj_4272));
    defparam i15_4_lut_adj_1336.LUT_INIT = 16'hfeff;
    SB_LUT4 select_622_Select_14_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4311));
    defparam select_622_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_15_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4309));
    defparam select_622_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1337 (.I0(n34776), .I1(\FRAME_MATCHER.state [24]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4249));
    defparam i1_2_lut_adj_1337.LUT_INIT = 16'h8888;
    SB_LUT4 select_622_Select_16_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4307));
    defparam select_622_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_17_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4305));
    defparam select_622_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i4_4_lut_adj_1338 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4493));   // verilog/coms.v(238[12:32])
    defparam i4_4_lut_adj_1338.LUT_INIT = 16'h7bde;
    SB_LUT4 i21813_2_lut (.I0(\FRAME_MATCHER.state [29]), .I1(n34776), .I2(GND_net), 
            .I3(GND_net), .O(n35323));
    defparam i21813_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1339 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4494));   // verilog/coms.v(238[12:32])
    defparam i2_4_lut_adj_1339.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1340 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_4495));   // verilog/coms.v(238[12:32])
    defparam i3_4_lut_adj_1340.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1341 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_4496));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut_adj_1341.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1342 (.I0(n9_adj_4496), .I1(n11_adj_4495), .I2(n10_adj_4494), 
            .I3(n12_adj_4493), .O(n25302));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut_adj_1342.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1343 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n126), .I3(\FRAME_MATCHER.state [2]), .O(n5_adj_4219));
    defparam i1_4_lut_adj_1343.LUT_INIT = 16'hfeff;
    SB_LUT4 select_622_Select_18_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4303));
    defparam select_622_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_19_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4301));
    defparam select_622_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1344 (.I0(n34776), .I1(\FRAME_MATCHER.state [30]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4247));
    defparam i1_2_lut_adj_1344.LUT_INIT = 16'h8888;
    SB_LUT4 i3_3_lut_adj_1345 (.I0(n5_adj_4219), .I1(n25302), .I2(n31_adj_4272), 
            .I3(GND_net), .O(n48426));
    defparam i3_3_lut_adj_1345.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1346 (.I0(\FRAME_MATCHER.state [12]), .I1(\FRAME_MATCHER.state [9]), 
            .I2(\FRAME_MATCHER.state [15]), .I3(\FRAME_MATCHER.state [10]), 
            .O(n10_adj_4497));
    defparam i4_4_lut_adj_1346.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1347 (.I0(\FRAME_MATCHER.state [8]), .I1(n10_adj_4497), 
            .I2(\FRAME_MATCHER.state [11]), .I3(GND_net), .O(n45517));
    defparam i5_3_lut_adj_1347.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1348 (.I0(\FRAME_MATCHER.state [5]), .I1(\FRAME_MATCHER.state [6]), 
            .I2(\FRAME_MATCHER.state [7]), .I3(\FRAME_MATCHER.state [4]), 
            .O(n36131));
    defparam i3_4_lut_adj_1348.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1349 (.I0(\FRAME_MATCHER.state [26]), .I1(\FRAME_MATCHER.state [25]), 
            .I2(\FRAME_MATCHER.state [20]), .I3(\FRAME_MATCHER.state [18]), 
            .O(n45610));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1349.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1350 (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [30]), 
            .I2(\FRAME_MATCHER.state [23]), .I3(\FRAME_MATCHER.state [29]), 
            .O(n20_adj_4498));
    defparam i8_4_lut_adj_1350.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1351 (.I0(\FRAME_MATCHER.state [24]), .I1(\FRAME_MATCHER.state [28]), 
            .I2(\FRAME_MATCHER.state [19]), .I3(\FRAME_MATCHER.state [21]), 
            .O(n19_adj_4499));
    defparam i7_4_lut_adj_1351.LUT_INIT = 16'hfffe;
    SB_LUT4 select_622_Select_20_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4299));
    defparam select_622_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i9_4_lut_adj_1352 (.I0(\FRAME_MATCHER.state [16]), .I1(\FRAME_MATCHER.state [17]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [27]), 
            .O(n21_adj_4500));
    defparam i9_4_lut_adj_1352.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut_adj_1353 (.I0(n21_adj_4500), .I1(n19_adj_4499), .I2(n20_adj_4498), 
            .I3(GND_net), .O(n45638));
    defparam i11_3_lut_adj_1353.LUT_INIT = 16'hfefe;
    SB_LUT4 select_622_Select_21_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4297));
    defparam select_622_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1354 (.I0(n25059), .I1(n3684), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4409));
    defparam i1_2_lut_adj_1354.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_1355 (.I0(\FRAME_MATCHER.i_31__N_2626 ), .I1(n25059), 
            .I2(n4452), .I3(GND_net), .O(n2_adj_4432));
    defparam i1_3_lut_adj_1355.LUT_INIT = 16'h0808;
    SB_LUT4 i4_4_lut_adj_1356 (.I0(n45610), .I1(n36131), .I2(n45517), 
            .I3(n6_adj_4501), .O(n39679));
    defparam i4_4_lut_adj_1356.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1357 (.I0(\FRAME_MATCHER.state[0] ), .I1(n39679), 
            .I2(GND_net), .I3(GND_net), .O(n126));
    defparam i1_2_lut_adj_1357.LUT_INIT = 16'heeee;
    SB_LUT4 select_622_Select_22_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4295));
    defparam select_622_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1358 (.I0(n25059), .I1(n3303), .I2(GND_net), 
            .I3(GND_net), .O(n25249));
    defparam i1_2_lut_adj_1358.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1359 (.I0(n771), .I1(n25059), .I2(GND_net), .I3(GND_net), 
            .O(n25262));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_adj_1359.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1360 (.I0(n39685), .I1(n25262), .I2(n25249), 
            .I3(n33), .O(n9_adj_4410));
    defparam i1_4_lut_adj_1360.LUT_INIT = 16'h50dc;
    SB_LUT4 select_622_Select_23_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4293));
    defparam select_622_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_24_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4291));
    defparam select_622_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_25_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4289));
    defparam select_622_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_26_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4287));
    defparam select_622_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 n53125_bdd_4_lut (.I0(n53125), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n53128));
    defparam n53125_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_622_Select_27_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4285));
    defparam select_622_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_28_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4283));
    defparam select_622_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_29_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4281));
    defparam select_622_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_30_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4279));
    defparam select_622_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_31_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4276));
    defparam select_622_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_622_Select_0_i3_2_lut_4_lut (.I0(n36137), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27968), .I3(\FRAME_MATCHER.i [0]), .O(n3));
    defparam select_622_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_4_lut_adj_1361 (.I0(\FRAME_MATCHER.state [2]), .I1(n126), 
            .I2(\FRAME_MATCHER.state [3]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n27974));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_4_lut_adj_1361.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(n45638), .I3(GND_net), .O(n6_adj_4501));
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(n45517), .I3(GND_net), .O(n36340));
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut_3_lut_adj_1364 (.I0(n34_adj_4502), .I1(n45_adj_4503), 
            .I2(n49), .I3(GND_net), .O(n47441));   // verilog/coms.v(115[11:12])
    defparam i2_2_lut_3_lut_adj_1364.LUT_INIT = 16'hfefe;
    SB_LUT4 i16214_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45612), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n29736));
    defparam i16214_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16215_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45612), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n29737));
    defparam i16215_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16216_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45612), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n29738));
    defparam i16216_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16217_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45612), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n29739));
    defparam i16217_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16218_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45612), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n29740));
    defparam i16218_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2660_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_4218));
    defparam i2660_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i16219_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45612), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n29741));
    defparam i16219_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16220_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45612), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n29742));
    defparam i16220_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16221_3_lut_4_lut (.I0(n8_adj_4328), .I1(n45612), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n29743));
    defparam i16221_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1365 (.I0(\FRAME_MATCHER.state [3]), .I1(n39679), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n39684));
    defparam i2_3_lut_adj_1365.LUT_INIT = 16'hefef;
    SB_LUT4 i36890_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n27916), .I3(n36614), .O(n27917));
    defparam i36890_3_lut_4_lut.LUT_INIT = 16'h010f;
    SB_LUT4 i22622_2_lut_4_lut (.I0(n45_adj_4503), .I1(n34_adj_4502), .I2(n7_adj_4409), 
            .I3(\FRAME_MATCHER.state [10]), .O(n36142));
    defparam i22622_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(n5389), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n36614), .I3(GND_net), .O(n27916));
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'haeae;
    SB_LUT4 i37607_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n29367));
    defparam i37607_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n1), .O(n5_adj_4504));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h1d11;
    SB_LUT4 i22594_2_lut_4_lut (.I0(n25302), .I1(n31_adj_4272), .I2(n31), 
            .I3(\FRAME_MATCHER.state [1]), .O(n1));
    defparam i22594_2_lut_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i22623_2_lut_4_lut (.I0(n45_adj_4503), .I1(n34_adj_4502), .I2(n7_adj_4409), 
            .I3(\FRAME_MATCHER.state [12]), .O(n36144));
    defparam i22623_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i36903_3_lut_4_lut (.I0(n46585), .I1(n5389), .I2(n39678), 
            .I3(n39690), .O(n48025));
    defparam i36903_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i22624_2_lut_4_lut (.I0(n45_adj_4503), .I1(n34_adj_4502), .I2(n7_adj_4409), 
            .I3(\FRAME_MATCHER.state [17]), .O(n36146));
    defparam i22624_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1367 (.I0(n45_adj_4503), .I1(n34_adj_4502), 
            .I2(n7_adj_4409), .I3(\FRAME_MATCHER.state [18]), .O(n36148));
    defparam i1_2_lut_4_lut_adj_1367.LUT_INIT = 16'hfe00;
    SB_LUT4 i16206_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45612), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n29728));
    defparam i16206_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34677_3_lut_4_lut (.I0(n4_adj_4357), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(\data_in_frame[2] [2]), .O(n50049));
    defparam i34677_3_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i16207_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45612), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n29729));
    defparam i16207_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16208_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45612), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n29730));
    defparam i16208_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16209_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45612), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n29731));
    defparam i16209_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [5]), 
            .I2(n28992), .I3(GND_net), .O(n45770));   // verilog/coms.v(70[16:62])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1369 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(n45833), .I3(n46178), .O(n42897));
    defparam i1_2_lut_3_lut_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1370 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[5] [7]), .I3(\data_out_frame[6] [1]), .O(n1241));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1371 (.I0(n28219), .I1(n45969), .I2(n46328), 
            .I3(n46374), .O(n45893));
    defparam i1_2_lut_3_lut_4_lut_adj_1371.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1372 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[6] [2]), .I3(n45926), .O(n46187));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut_4_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[6] [2]), .I3(\data_out_frame[15] [0]), .O(n16_adj_4386));   // verilog/coms.v(73[16:42])
    defparam i5_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16210_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45612), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n29732));
    defparam i16210_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16211_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45612), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n29733));
    defparam i16211_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_2_lut_3_lut_4_lut (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[17] [1]), .I3(\data_out_frame[17] [0]), 
            .O(n42_adj_4413));   // verilog/coms.v(74[16:43])
    defparam i4_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i44_1_lut_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n39684), .I3(GND_net), .O(n2987));
    defparam i44_1_lut_2_lut_3_lut.LUT_INIT = 16'h0707;
    SB_LUT4 i16212_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45612), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n29734));
    defparam i16212_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16213_3_lut_4_lut (.I0(n8_adj_4336), .I1(n45612), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n29735));
    defparam i16213_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1373 (.I0(\data_in_frame[19] [5]), .I1(n28651), 
            .I2(n45738), .I3(\data_in_frame[19] [6]), .O(n45913));
    defparam i1_2_lut_3_lut_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(n28299), .I1(\data_in_frame[6] [0]), 
            .I2(n28219), .I3(GND_net), .O(n6_adj_4442));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1375 (.I0(tx_active), .I1(r_SM_Main_2__N_3616[0]), 
            .I2(tx_transmit_N_3513), .I3(n39686), .O(n45588));
    defparam i1_2_lut_3_lut_4_lut_adj_1375.LUT_INIT = 16'h00fe;
    SB_LUT4 i2_2_lut_3_lut_adj_1376 (.I0(n28299), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[3] [6]), .I3(GND_net), .O(n8_adj_4459));   // verilog/coms.v(76[16:43])
    defparam i2_2_lut_3_lut_adj_1376.LUT_INIT = 16'h9696;
    SB_LUT4 i13_3_lut_4_lut (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(n28992), .I3(n28937), .O(n31_adj_4429));
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1377 (.I0(n28651), .I1(\data_in_frame[17] [5]), 
            .I2(n46075), .I3(\data_in_frame[19] [6]), .O(n46319));
    defparam i1_2_lut_3_lut_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i22341_2_lut_3_lut (.I0(n36137), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n35859));
    defparam i22341_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[6] [6]), .I3(\data_in_frame[2] [2]), .O(n10_adj_4455));   // verilog/coms.v(73[16:27])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n28299));
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n39684), .I3(GND_net), .O(n36137));
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'hf8f8;
    SB_LUT4 i16198_3_lut_4_lut (.I0(n36193), .I1(n45612), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n29720));
    defparam i16198_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16199_3_lut_4_lut (.I0(n36193), .I1(n45612), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n29721));
    defparam i16199_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1380 (.I0(n34_adj_4502), .I1(n45_adj_4503), 
            .I2(n25059), .I3(n3684), .O(n34776));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_3_lut_4_lut_adj_1380.LUT_INIT = 16'hfeee;
    SB_LUT4 i16200_3_lut_4_lut (.I0(n36193), .I1(n45612), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n29722));
    defparam i16200_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1381 (.I0(\FRAME_MATCHER.state [2]), 
            .I1(\FRAME_MATCHER.state[0] ), .I2(n39679), .I3(\FRAME_MATCHER.state [1]), 
            .O(n27968));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1381.LUT_INIT = 16'hfffe;
    SB_LUT4 i16201_3_lut_4_lut (.I0(n36193), .I1(n45612), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n29723));
    defparam i16201_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16202_3_lut_4_lut (.I0(n36193), .I1(n45612), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n29724));
    defparam i16202_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16203_3_lut_4_lut (.I0(n36193), .I1(n45612), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n29725));
    defparam i16203_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16204_3_lut_4_lut (.I0(n36193), .I1(n45612), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n29726));
    defparam i16204_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16205_3_lut_4_lut (.I0(n36193), .I1(n45612), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n29727));
    defparam i16205_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_4_lut_adj_1382 (.I0(n35330), .I1(tx_transmit_N_3513), 
            .I2(n25059), .I3(n39686), .O(n49));
    defparam i1_3_lut_4_lut_adj_1382.LUT_INIT = 16'h00e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1383 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[4] [4]), .O(n46067));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n45656));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i71_2_lut_3_lut (.I0(n113), .I1(n25059), .I2(n3303), .I3(GND_net), 
            .O(n34_adj_4502));   // verilog/coms.v(115[11:12])
    defparam i71_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_adj_1385 (.I0(\data_in_frame[11] [5]), .I1(n42840), 
            .I2(n45719), .I3(GND_net), .O(n42915));
    defparam i1_2_lut_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1386 (.I0(\data_in_frame[11] [5]), .I1(n42840), 
            .I2(n45684), .I3(n46036), .O(n43591));
    defparam i2_3_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i74_2_lut_3_lut (.I0(n114), .I1(n771), .I2(n25059), .I3(GND_net), 
            .O(n45_adj_4503));   // verilog/coms.v(115[11:12])
    defparam i74_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[14] [1]), .I3(GND_net), .O(n46345));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1388 (.I0(n28226), .I1(n45825), .I2(n45722), 
            .I3(GND_net), .O(n28881));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1388.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1389 (.I0(n28657), .I1(n28226), .I2(\data_in_frame[10] [5]), 
            .I3(\data_in_frame[12] [6]), .O(n45722));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1390 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[9] [2]), .I3(GND_net), .O(n28074));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1391 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [5]), .I3(GND_net), .O(n45811));   // verilog/coms.v(75[16:27])
    defparam i2_2_lut_3_lut_adj_1391.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1392 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[6] [2]), .I3(GND_net), .O(n46247));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1392.LUT_INIT = 16'h9696;
    SB_LUT4 i16190_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45628), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n29712));
    defparam i16190_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1393 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(\data_in_frame[3] [7]), .O(n45671));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1394 (.I0(\data_in_frame[10] [4]), .I1(Kp_23__N_1183), 
            .I2(\data_in_frame[8] [2]), .I3(GND_net), .O(n45825));   // verilog/coms.v(74[16:43])
    defparam i2_2_lut_3_lut_adj_1394.LUT_INIT = 16'h9696;
    SB_LUT4 i16191_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45628), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n29713));
    defparam i16191_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1395 (.I0(\FRAME_MATCHER.state [3]), .I1(n25059), 
            .I2(n3684), .I3(n2_adj_4432), .O(n44957));
    defparam i1_3_lut_4_lut_adj_1395.LUT_INIT = 16'haa80;
    SB_LUT4 i16192_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45628), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n29714));
    defparam i16192_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16193_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45628), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n29715));
    defparam i16193_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1396 (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[15] [5]), 
            .I2(n28581), .I3(\data_in_frame[13] [3]), .O(n46219));
    defparam i1_2_lut_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1397 (.I0(n28232), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[11] [1]), .I3(GND_net), .O(n45716));
    defparam i1_2_lut_3_lut_adj_1397.LUT_INIT = 16'h9696;
    SB_LUT4 i16194_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45628), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n29716));
    defparam i16194_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1398 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n123_c));   // verilog/coms.v(102[12:33])
    defparam i1_2_lut_adj_1398.LUT_INIT = 16'h8888;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1399 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(n46024), .I3(GND_net), .O(n6_adj_4457));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_3_lut_adj_1399.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1400 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[2] [0]), .I3(GND_net), .O(n46297));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_3_lut_adj_1400.LUT_INIT = 16'h9696;
    SB_LUT4 i16195_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45628), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n29717));
    defparam i16195_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16196_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45628), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n29718));
    defparam i16196_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1401 (.I0(Kp_23__N_1237), .I1(\data_in_frame[11] [4]), 
            .I2(Kp_23__N_1217), .I3(n28074), .O(n45684));
    defparam i2_3_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[5] [0]), 
            .I2(n28673), .I3(n28937), .O(n12_adj_4456));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1402 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(n4_adj_4357), .I3(GND_net), .O(n28673));   // verilog/coms.v(70[16:27])
    defparam i2_2_lut_3_lut_adj_1402.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1403 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[1] [0]), 
            .I2(Kp_23__N_988), .I3(GND_net), .O(n26983));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 i16197_3_lut_4_lut (.I0(n8_adj_4217), .I1(n45628), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n29719));
    defparam i16197_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n46585), .O(n29243));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_3_lut_4_lut_adj_1404 (.I0(\data_out_frame[23] [3]), .I1(n42923), 
            .I2(\data_out_frame[23] [4]), .I3(n42958), .O(n43943));
    defparam i2_3_lut_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(n42875), .I1(\data_out_frame[20] [7]), 
            .I2(n27578), .I3(GND_net), .O(n42958));
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1406 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[1] [6]), .O(n19_adj_4505));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1406.LUT_INIT = 16'h6900;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1407 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [2]), 
            .I2(n46356), .I3(n45652), .O(Kp_23__N_988));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1408 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[0] [7]), .O(n46237));   // verilog/coms.v(73[16:34])
    defparam i2_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1409 (.I0(\data_in_frame[15] [0]), .I1(n29005), 
            .I2(n45815), .I3(GND_net), .O(n10_adj_4448));   // verilog/coms.v(76[16:43])
    defparam i2_2_lut_3_lut_adj_1409.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1410 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n46059));
    defparam i1_2_lut_3_lut_adj_1410.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1411 (.I0(n45652), .I1(n46356), .I2(\data_in_frame[3] [1]), 
            .I3(\data_in_frame[3] [3]), .O(n29005));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_3_lut_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1412 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n10_adj_4506));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_adj_1412.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(n29005), .I1(n45815), .I2(n45851), 
            .I3(GND_net), .O(n28146));
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1414 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(n45997), .I3(n45694), .O(n8_adj_4355));   // verilog/coms.v(70[16:27])
    defparam i3_3_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1415 (.I0(n28287), .I1(\data_in_frame[9] [7]), 
            .I2(n46359), .I3(GND_net), .O(n45851));
    defparam i1_2_lut_3_lut_adj_1415.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1416 (.I0(\data_in_frame[5] [5]), .I1(n46237), 
            .I2(\data_in_frame[7] [7]), .I3(n28299), .O(n45923));
    defparam i2_3_lut_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1417 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [4]), 
            .I2(n28544), .I3(GND_net), .O(n45719));
    defparam i1_2_lut_3_lut_adj_1417.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1418 (.I0(n42799), .I1(\data_out_frame[16] [4]), 
            .I2(n42805), .I3(GND_net), .O(n28584));
    defparam i1_2_lut_3_lut_adj_1418.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[4] [6]), .O(n46056));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1420 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[10] [1]), 
            .I2(n10_adj_4433), .I3(\data_out_frame[5] [7]), .O(n28014));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[0] [1]), 
            .I2(n45656), .I3(n11_adj_4364), .O(n46014));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[0] [1]), 
            .I2(n45656), .I3(GND_net), .O(n46244));
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1422 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n46285));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1422.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1423 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[4] [0]), .I3(\data_out_frame[6] [1]), .O(n45782));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1424 (.I0(n28645), .I1(n28213), .I2(\data_in_frame[6] [6]), 
            .I3(\data_in_frame[6] [1]), .O(n6_adj_4430));   // verilog/coms.v(85[17:28])
    defparam i2_2_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1425 (.I0(\data_out_frame[13] [7]), .I1(n46203), 
            .I2(n42805), .I3(\data_out_frame[16] [3]), .O(n42795));
    defparam i2_3_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1426 (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[5] [4]), 
            .I2(n28771), .I3(GND_net), .O(n28120));
    defparam i1_2_lut_3_lut_adj_1426.LUT_INIT = 16'h9696;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[12] [6]), .I3(\data_out_frame[12] [5]), 
            .O(n45_adj_4420));   // verilog/coms.v(85[17:28])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(n42822), .I3(\data_out_frame[13] [5]), .O(n18_adj_4423));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1427 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n46291));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1427.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1428 (.I0(\data_out_frame[13] [4]), .I1(n28800), 
            .I2(n42820), .I3(\data_out_frame[15] [5]), .O(n43923));
    defparam i2_3_lut_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1429 (.I0(n1510), .I1(\data_out_frame[12] [2]), 
            .I2(\data_out_frame[14] [3]), .I3(n46086), .O(n42799));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1430 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[5] [2]), .I3(n46291), .O(n8_adj_4407));
    defparam i2_2_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1431 (.I0(n1510), .I1(\data_out_frame[12] [2]), 
            .I2(n28014), .I3(\data_out_frame[14] [4]), .O(n45807));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i16182_3_lut_4_lut (.I0(n10_adj_4506), .I1(n45606), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n29704));
    defparam i16182_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_2053_i7_2_lut_3_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n7_adj_4406));   // verilog/coms.v(166[9:87])
    defparam equal_2053_i7_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1432 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[9] [5]), .I3(GND_net), .O(n45688));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_adj_1432.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1433 (.I0(n35859), .I1(n10_adj_4506), .I2(GND_net), 
            .I3(GND_net), .O(n45628));
    defparam i1_2_lut_adj_1433.LUT_INIT = 16'hdddd;
    SB_LUT4 i16183_3_lut_4_lut (.I0(n10_adj_4506), .I1(n45606), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n29705));
    defparam i16183_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1434 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(n46122), .I3(\data_out_frame[6] [5]), .O(n45788));
    defparam i2_3_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1435 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[11] [2]), .I3(n45785), .O(n46163));   // verilog/coms.v(71[16:62])
    defparam i2_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i16184_3_lut_4_lut (.I0(n10_adj_4506), .I1(n45606), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n29706));
    defparam i16184_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16185_3_lut_4_lut (.I0(n10_adj_4506), .I1(n45606), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n29707));
    defparam i16185_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut_adj_1436 (.I0(n28533), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[13] [4]), .I3(n46133), .O(n8_adj_4401));
    defparam i3_3_lut_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1437 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[11] [0]), .I3(n46111), .O(n6_adj_4402));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i16186_3_lut_4_lut (.I0(n10_adj_4506), .I1(n45606), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n29708));
    defparam i16186_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16187_3_lut_4_lut (.I0(n10_adj_4506), .I1(n45606), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n29709));
    defparam i16187_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1438 (.I0(\data_out_frame[15] [7]), .I1(n45807), 
            .I2(\data_out_frame[16] [5]), .I3(n42799), .O(n45990));
    defparam i1_2_lut_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i16188_3_lut_4_lut (.I0(n10_adj_4506), .I1(n45606), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n29710));
    defparam i16188_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16189_3_lut_4_lut (.I0(n10_adj_4506), .I1(n45606), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n29711));
    defparam i16189_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1439 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[11] [0]), .I3(GND_net), .O(n45741));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1439.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1440 (.I0(\data_out_frame[12] [6]), .I1(n27527), 
            .I2(\data_out_frame[14] [6]), .I3(\data_out_frame[14] [7]), 
            .O(n6_adj_4388));
    defparam i1_2_lut_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1441 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n28456));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1442 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[6] [1]), 
            .I2(n45704), .I3(n45926), .O(n6_adj_4381));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1443 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n22_adj_4373));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_3_lut_adj_1443.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1444 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[16] [6]), 
            .I2(n45807), .I3(GND_net), .O(n46350));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1444.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1445 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n6_adj_4376));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1445.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1446 (.I0(n28287), .I1(n28226), .I2(n45825), 
            .I3(\data_in_frame[12] [5]), .O(n46077));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1447 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[9] [0]), .I3(GND_net), .O(n46304));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1447.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1448 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[13] [6]), .I3(\data_out_frame[16] [2]), 
            .O(n46371));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i16174_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45628), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n29696));
    defparam i16174_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16175_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45628), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n29697));
    defparam i16175_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16176_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45628), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n29698));
    defparam i16176_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16177_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45628), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n29699));
    defparam i16177_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1449 (.I0(n28259), .I1(\data_in_frame[9] [6]), 
            .I2(n28264), .I3(\data_in_frame[9] [7]), .O(n42581));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1450 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[8] [6]), 
            .I2(Kp_23__N_1195), .I3(n45804), .O(n46338));
    defparam i1_2_lut_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(\data_in_frame[8] [6]), .I1(Kp_23__N_1195), 
            .I2(n45804), .I3(GND_net), .O(n28140));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1452 (.I0(\data_in_frame[7] [2]), .I1(n28259), 
            .I2(Kp_23__N_1217), .I3(n46377), .O(n6_adj_4354));
    defparam i1_2_lut_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1453 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [3]), 
            .I2(n28912), .I3(GND_net), .O(n46153));
    defparam i1_2_lut_3_lut_adj_1453.LUT_INIT = 16'h9696;
    SB_LUT4 i16178_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45628), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n29700));
    defparam i16178_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1454 (.I0(\data_out_frame[17] [4]), .I1(n27527), 
            .I2(\data_out_frame[13] [0]), .I3(n28526), .O(n45872));
    defparam i2_3_lut_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1455 (.I0(\data_out_frame[15] [3]), .I1(n45878), 
            .I2(n10_adj_4393), .I3(\data_out_frame[12] [7]), .O(n45674));
    defparam i1_2_lut_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1456 (.I0(n45707), .I1(n46056), .I2(n10_adj_4348), 
            .I3(\data_out_frame[16] [2]), .O(n45749));
    defparam i5_3_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(n42875), .I1(\data_out_frame[20] [7]), 
            .I2(n45744), .I3(GND_net), .O(n46178));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'h9696;
    SB_LUT4 i16179_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45628), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n29701));
    defparam i16179_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1458 (.I0(n28342), .I1(n46348), .I2(\data_out_frame[20] [4]), 
            .I3(n46082), .O(n6_adj_4347));
    defparam i1_2_lut_4_lut_adj_1458.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1459 (.I0(n45959), .I1(n43593), .I2(n46362), 
            .I3(n45840), .O(n47585));
    defparam i2_3_lut_4_lut_adj_1459.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1460 (.I0(\data_out_frame[20] [1]), .I1(n43883), 
            .I2(\data_out_frame[20] [2]), .I3(n43850), .O(n45959));
    defparam i1_2_lut_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1461 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[25] [6]), .I3(n45956), .O(n6_adj_4344));
    defparam i2_2_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1462 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[25] [6]), .I3(GND_net), .O(n46316));
    defparam i1_2_lut_3_lut_adj_1462.LUT_INIT = 16'h9696;
    SB_LUT4 i9_3_lut_4_lut (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(\data_out_frame[23] [2]), .I3(\data_out_frame[23] [1]), 
            .O(n26));
    defparam i9_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1463 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[17] [6]), 
            .I2(n28526), .I3(GND_net), .O(n46335));
    defparam i1_2_lut_3_lut_adj_1463.LUT_INIT = 16'h9696;
    SB_LUT4 i16180_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45628), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n29702));
    defparam i16180_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16181_3_lut_4_lut (.I0(n8_adj_4274), .I1(n45628), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n29703));
    defparam i16181_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1464 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[17] [6]), 
            .I2(n43923), .I3(GND_net), .O(n6_adj_4339));
    defparam i1_2_lut_3_lut_adj_1464.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1465 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n35859), .O(n45606));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1465.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_1466 (.I0(\data_out_frame[20] [1]), .I1(n43883), 
            .I2(\data_out_frame[24] [3]), .I3(GND_net), .O(n45862));
    defparam i1_2_lut_3_lut_adj_1466.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1467 (.I0(n1516), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n45972));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1467.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1468 (.I0(n43866), .I1(n42781), .I2(n43437), 
            .I3(\data_out_frame[19] [5]), .O(n45884));
    defparam i2_3_lut_4_lut_adj_1468.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1469 (.I0(n1516), .I1(\data_out_frame[12] [4]), 
            .I2(n10_adj_4449), .I3(n28014), .O(n45833));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1470 (.I0(n43876), .I1(\data_out_frame[19] [3]), 
            .I2(n45867), .I3(\data_out_frame[23] [6]), .O(n6_adj_4334));
    defparam i1_2_lut_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i16166_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45628), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29688));
    defparam i16166_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16167_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45628), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29689));
    defparam i16167_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16168_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45628), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n29690));
    defparam i16168_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16169_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45628), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29691));
    defparam i16169_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16170_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45628), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29692));
    defparam i16170_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16171_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45628), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29693));
    defparam i16171_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16172_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45628), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29694));
    defparam i16172_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16173_3_lut_4_lut (.I0(n8_adj_4277), .I1(n45628), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29695));
    defparam i16173_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1471 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[16] [0]), 
            .I2(n28800), .I3(GND_net), .O(n6_adj_4346));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 i16158_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45628), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n29680));
    defparam i16158_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16159_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45628), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n29681));
    defparam i16159_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16160_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45628), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n29682));
    defparam i16160_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16161_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45628), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n29683));
    defparam i16161_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16162_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45628), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n29684));
    defparam i16162_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16163_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45628), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n29685));
    defparam i16163_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4395));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16164_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45628), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n29686));
    defparam i16164_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16165_3_lut_4_lut (.I0(n8_adj_4332), .I1(n45628), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n29687));
    defparam i16165_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4394));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36039_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n51338));
    defparam i36039_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36036_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n51337));
    defparam i36036_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1472 (.I0(\data_in_frame[7] [2]), .I1(n28259), 
            .I2(Kp_23__N_1217), .I3(GND_net), .O(n46049));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1472.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1473 (.I0(\data_in_frame[7] [2]), .I1(n28259), 
            .I2(n46225), .I3(\data_in_frame[11] [6]), .O(n8_adj_4472));   // verilog/coms.v(74[16:43])
    defparam i3_3_lut_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i34882_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50364));
    defparam i34882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34883_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50365));
    defparam i34883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1474 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[11] [2]), .I3(n4_adj_4271), .O(n45804));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1475 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[9] [2]), .I3(\data_in_frame[11] [7]), .O(n45644));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1476 (.I0(\data_out_frame[4] [5]), .I1(n45785), 
            .I2(\data_out_frame[6] [4]), .I3(n45821), .O(n28447));   // verilog/coms.v(71[16:62])
    defparam i2_3_lut_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1477 (.I0(\data_out_frame[4] [5]), .I1(n45785), 
            .I2(\data_out_frame[6] [7]), .I3(GND_net), .O(n45887));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_3_lut_adj_1477.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1478 (.I0(tx_active), .I1(r_SM_Main_2__N_3616[0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n6_adj_4333));
    defparam i2_2_lut_3_lut_adj_1478.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1479 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n39684), .I3(GND_net), .O(n39686));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1479.LUT_INIT = 16'hf7f7;
    SB_LUT4 i4_3_lut_4_lut (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[9] [2]), .O(n11_adj_4370));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1480 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[7] [3]), .I3(n45887), .O(n8_adj_4398));
    defparam i3_3_lut_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1481 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n6935));
    defparam i1_2_lut_3_lut_adj_1481.LUT_INIT = 16'h0202;
    SB_LUT4 i4_2_lut_4_lut_adj_1482 (.I0(\data_out_frame[4] [0]), .I1(n45902), 
            .I2(\data_out_frame[6] [2]), .I3(n28466), .O(n18_adj_4350));   // verilog/coms.v(75[16:43])
    defparam i4_2_lut_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1483 (.I0(\data_out_frame[4] [0]), .I1(n45902), 
            .I2(\data_out_frame[6] [2]), .I3(n45640), .O(n28068));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1484 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n36614), .I3(n35330), .O(n8_adj_4331));
    defparam i3_3_lut_4_lut_adj_1484.LUT_INIT = 16'h0080;
    SB_LUT4 i2_3_lut_4_lut_adj_1485 (.I0(n45971), .I1(n46328), .I2(\data_in_frame[12] [4]), 
            .I3(n28287), .O(n42881));
    defparam i2_3_lut_4_lut_adj_1485.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_adj_1486 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[13] [2]), .I3(GND_net), .O(n10_adj_4375));   // verilog/coms.v(73[16:42])
    defparam i2_2_lut_3_lut_adj_1486.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1487 (.I0(n2076), .I1(n45833), .I2(\data_out_frame[19] [1]), 
            .I3(n26083), .O(n45859));
    defparam i2_3_lut_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1488 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(Kp_23__N_1195), .I3(n45969), .O(n11));
    defparam i1_3_lut_4_lut_adj_1488.LUT_INIT = 16'h7dbe;
    SB_LUT4 i1_2_lut_adj_1489 (.I0(\data_in_frame[0] [5]), .I1(n28992), 
            .I2(GND_net), .I3(GND_net), .O(n28108));   // verilog/coms.v(70[16:62])
    defparam i1_2_lut_adj_1489.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1490 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[1] [7]), 
            .I2(n45773), .I3(n45770), .O(n22_adj_4507));
    defparam i5_4_lut_adj_1490.LUT_INIT = 16'h1248;
    SB_LUT4 i1_2_lut_adj_1491 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4508));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1491.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1492 (.I0(n25302), .I1(n22_adj_4507), .I2(\data_in_frame[2] [0]), 
            .I3(n45770), .O(n28_adj_4509));
    defparam i11_4_lut_adj_1492.LUT_INIT = 16'h4004;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37639 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n53119));
    defparam byte_transmit_counter_0__bdd_4_lut_37639.LUT_INIT = 16'he4aa;
    SB_LUT4 n53119_bdd_4_lut (.I0(n53119), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n53122));
    defparam n53119_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i23081_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n36612), .O(n36614));   // verilog/coms.v(127[12] 300[6])
    defparam i23081_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37634 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n53113));
    defparam byte_transmit_counter_0__bdd_4_lut_37634.LUT_INIT = 16'he4aa;
    SB_LUT4 i34679_4_lut (.I0(Kp_23__N_979), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[2] [4]), .I3(n4_adj_4508), .O(n50051));
    defparam i34679_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i13_4_lut_adj_1493 (.I0(n50049), .I1(n7_adj_4406), .I2(\data_in_frame[1] [4]), 
            .I3(\data_in_frame[1] [5]), .O(n30_adj_4510));
    defparam i13_4_lut_adj_1493.LUT_INIT = 16'h1000;
    SB_LUT4 i6_4_lut_adj_1494 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[1] [1]), .I3(n28108), .O(n23));
    defparam i6_4_lut_adj_1494.LUT_INIT = 16'h2184;
    SB_LUT4 i14_4_lut_adj_1495 (.I0(n19_adj_4505), .I1(n28_adj_4509), .I2(\data_in_frame[1] [2]), 
            .I3(\data_in_frame[1] [3]), .O(n31_adj_4511));
    defparam i14_4_lut_adj_1495.LUT_INIT = 16'h8000;
    SB_LUT4 i16_4_lut_adj_1496 (.I0(n31_adj_4511), .I1(n23), .I2(n30_adj_4510), 
            .I3(n50051), .O(\FRAME_MATCHER.state_31__N_2724 [3]));
    defparam i16_4_lut_adj_1496.LUT_INIT = 16'h0080;
    SB_LUT4 i3_3_lut_adj_1497 (.I0(n5_adj_4269), .I1(n36131), .I2(n36340), 
            .I3(GND_net), .O(n46585));
    defparam i3_3_lut_adj_1497.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1498 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state_31__N_2724 [3]), 
            .O(n6_adj_4512));
    defparam i2_4_lut_adj_1498.LUT_INIT = 16'hccdc;
    SB_LUT4 i36925_4_lut (.I0(n27916), .I1(n36614), .I2(n5_adj_4504), 
            .I3(n6_adj_4512), .O(n45554));
    defparam i36925_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i2_2_lut_3_lut_adj_1499 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4217));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_adj_1499.LUT_INIT = 16'hfefe;
    SB_LUT4 n53113_bdd_4_lut (.I0(n53113), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n53116));
    defparam n53113_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1500 (.I0(\FRAME_MATCHER.state [3]), .I1(n5389), 
            .I2(n36614), .I3(GND_net), .O(n48518));
    defparam i2_3_lut_adj_1500.LUT_INIT = 16'h0101;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37629 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n53101));
    defparam byte_transmit_counter_0__bdd_4_lut_37629.LUT_INIT = 16'he4aa;
    SB_LUT4 n53101_bdd_4_lut (.I0(n53101), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n53104));
    defparam n53101_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_4_lut (.I0(\data_out_frame[5] [6]), .I1(n28068), .I2(\data_out_frame[10] [5]), 
            .I3(n45782), .O(n45664));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1501 (.I0(\data_out_frame[19] [3]), .I1(n45867), 
            .I2(\data_out_frame[19] [2]), .I3(n43916), .O(n42913));
    defparam i2_3_lut_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1502 (.I0(\data_out_frame[19] [3]), .I1(n45867), 
            .I2(\data_out_frame[23] [6]), .I3(GND_net), .O(n46141));
    defparam i1_2_lut_3_lut_adj_1502.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1503 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n39684), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2626 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1503.LUT_INIT = 16'h0202;
    SB_LUT4 i1_3_lut_4_lut_adj_1504 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n27908), .I3(\FRAME_MATCHER.i [1]), .O(n5));
    defparam i1_3_lut_4_lut_adj_1504.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_2_lut_adj_1505 (.I0(n35859), .I1(n10_adj_4245), .I2(GND_net), 
            .I3(GND_net), .O(n45620));
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_3_lut_4_lut_adj_1506 (.I0(\data_out_frame[19] [3]), .I1(n45867), 
            .I2(n46210), .I3(\data_out_frame[25] [7]), .O(n14_adj_4337));
    defparam i5_3_lut_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1507 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n39684), .I3(GND_net), .O(n113));
    defparam i1_2_lut_3_lut_adj_1507.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_4_lut_adj_1508 (.I0(n43235), .I1(n42795), .I2(\data_out_frame[20] [5]), 
            .I3(\data_out_frame[23] [1]), .O(n46082));
    defparam i1_2_lut_4_lut_adj_1508.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1509 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n39684), .I3(GND_net), .O(n114));
    defparam i1_2_lut_3_lut_adj_1509.LUT_INIT = 16'hfefe;
    uart_tx tx (.CLK_c(CLK_c), .n29165(n29165), .tx_o(tx_o), .tx_data({tx_data}), 
            .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3616[0] (r_SM_Main_2__N_3616[0]), 
            .\r_SM_Main_2__N_3613[1] (\r_SM_Main_2__N_3613[1] ), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .GND_net(GND_net), .n45528(n45528), .n29578(n29578), .n29579(n29579), 
            .tx_active(tx_active), .n53403(n53403), .VCC_net(VCC_net), 
            .n20247(n20247), .n4(n4), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.CLK_c(CLK_c), .n29175(n29175), .r_SM_Main({r_SM_Main_adj_18}), 
            .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), .\r_SM_Main_2__N_3542[2] (\r_SM_Main_2__N_3542[2] ), 
            .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_14 ), .n27903(n27903), 
            .GND_net(GND_net), .n4(n4_adj_15), .n45526(n45526), .n29587(n29587), 
            .rx_data({rx_data}), .n29582(n29582), .n45179(n45179), .rx_data_ready(rx_data_ready), 
            .n29561(n29561), .n29560(n29560), .n29559(n29559), .n29558(n29558), 
            .n29557(n29557), .n29556(n29556), .n29555(n29555), .n45591(n45591), 
            .VCC_net(VCC_net), .n4_adj_8(n4_adj_16), .n4_adj_9(n4_adj_17), 
            .n27898(n27898), .n35507(n35507)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (CLK_c, n29165, tx_o, tx_data, r_SM_Main, \r_SM_Main_2__N_3616[0] , 
            \r_SM_Main_2__N_3613[1] , \r_Bit_Index[0] , GND_net, n45528, 
            n29578, n29579, tx_active, n53403, VCC_net, n20247, 
            n4, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    output n29165;
    output tx_o;
    input [7:0]tx_data;
    output [2:0]r_SM_Main;
    input \r_SM_Main_2__N_3616[0] ;
    output \r_SM_Main_2__N_3613[1] ;
    output \r_Bit_Index[0] ;
    input GND_net;
    output n45528;
    input n29578;
    input n29579;
    output tx_active;
    input n53403;
    input VCC_net;
    output n20247;
    output n4;
    output tx_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [8:0]n41;
    
    wire n6852;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n29450;
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n29414, n3, n25082;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n21442;
    wire [2:0]r_SM_Main_2__N_3610;
    
    wire n50388, n50389, n50299, n50298, n3_adj_4212, n21441, o_Tx_Serial_N_3644, 
        n53203, n48013, n10, n41864, n41863, n41862, n41861, n41860, 
        n41859, n41858, n41857;
    
    SB_DFFESR r_Clock_Count_2065__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n6852), 
            .D(n41[3]), .R(n29450));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n6852), 
            .D(n41[2]), .R(n29450));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n6852), 
            .D(n41[1]), .R(n29450));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n6852), 
            .D(n41[0]), .R(n29450));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n29165), 
            .D(n307[1]), .R(n29414));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n29165), 
            .D(n307[2]), .R(n29414));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .E(n6852), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n25082), .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n21442), .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_2065__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n6852), 
            .D(n41[4]), .R(n29450));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3616[0] ), 
            .I3(r_SM_Main[1]), .O(n25082));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3610[0]), .O(n29414));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_870 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_3613[1] ), .O(n29165));
    defparam i1_3_lut_4_lut_adj_870.LUT_INIT = 16'h1101;
    SB_LUT4 i34906_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n50388));
    defparam i34906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34907_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n50389));
    defparam i34907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34817_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n50299));
    defparam i34817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34816_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n50298));
    defparam i34816_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n3_adj_4212), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n25082), .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n25082), .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n25082), .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n25082), .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n25082), .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n25082), .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n25082), .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_2065__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .E(n6852), 
            .D(n41[8]), .R(n29450));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i8054_3_lut (.I0(n21441), .I1(\r_SM_Main_2__N_3613[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n21442));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i8054_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3644), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFESR r_Clock_Count_2065__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n6852), 
            .D(n41[7]), .R(n29450));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n6852), 
            .D(n41[6]), .R(n29450));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n6852), 
            .D(n41[5]), .R(n29450));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i11338_2_lut_3_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4212));
    defparam i11338_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2200_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i2200_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n45528));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(n45528), .I1(\r_SM_Main_2__N_3613[1] ), .I2(GND_net), 
            .I3(GND_net), .O(r_SM_Main_2__N_3610[0]));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2193_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i2193_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n50298), 
            .I2(n50299), .I3(r_Bit_Index[2]), .O(n53203));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n53203_bdd_4_lut (.I0(n53203), .I1(n50389), .I2(n50388), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3644));
    defparam n53203_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n29578));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[2]), .O(n48013));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), .I2(n48013), 
            .I3(r_Clock_Count[8]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3613[1] ));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i36860_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3613[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n29450));
    defparam i36860_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1985_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n6852));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1985_1_lut.LUT_INIT = 16'h5555;
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n29579));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n53403));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_2065_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n41864), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2065_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n41863), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_9 (.CI(n41863), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n41864));
    SB_LUT4 r_Clock_Count_2065_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n41862), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_8 (.CI(n41862), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n41863));
    SB_LUT4 r_Clock_Count_2065_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n41861), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_7 (.CI(n41861), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n41862));
    SB_LUT4 r_Clock_Count_2065_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n41860), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_6 (.CI(n41860), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n41861));
    SB_LUT4 r_Clock_Count_2065_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n41859), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_5 (.CI(n41859), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n41860));
    SB_LUT4 r_Clock_Count_2065_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n41858), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_4 (.CI(n41858), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n41859));
    SB_LUT4 r_Clock_Count_2065_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n41857), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_3 (.CI(n41857), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n41858));
    SB_LUT4 r_Clock_Count_2065_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n41857));
    SB_LUT4 i6864_2_lut (.I0(\r_SM_Main_2__N_3616[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n20247));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i6864_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i8053_3_lut_4_lut (.I0(\r_SM_Main_2__N_3616[0] ), .I1(n45528), 
            .I2(\r_SM_Main_2__N_3613[1] ), .I3(r_SM_Main[1]), .O(n21441));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i8053_3_lut_4_lut.LUT_INIT = 16'hc0aa;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (CLK_c, n29175, r_SM_Main, r_Rx_Data, RX_N_10, \r_SM_Main_2__N_3542[2] , 
            \r_Bit_Index[0] , n27903, GND_net, n4, n45526, n29587, 
            rx_data, n29582, n45179, rx_data_ready, n29561, n29560, 
            n29559, n29558, n29557, n29556, n29555, n45591, VCC_net, 
            n4_adj_8, n4_adj_9, n27898, n35507) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    output n29175;
    output [2:0]r_SM_Main;
    output r_Rx_Data;
    input RX_N_10;
    output \r_SM_Main_2__N_3542[2] ;
    output \r_Bit_Index[0] ;
    output n27903;
    input GND_net;
    output n4;
    output n45526;
    input n29587;
    output [7:0]rx_data;
    input n29582;
    input n45179;
    output rx_data_ready;
    input n29561;
    input n29560;
    input n29559;
    input n29558;
    input n29557;
    input n29556;
    input n29555;
    input n45591;
    input VCC_net;
    output n4_adj_8;
    output n4_adj_9;
    output n27898;
    output n35507;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]n37;
    
    wire n29244;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n29448;
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n29416, n3, r_Rx_Data_R;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n27775, n36314;
    wire [2:0]r_SM_Main_2__N_3548;
    
    wire n1, n36198, n9, n27763, n6, n41856, n41855, n41854, 
        n41853, n41852, n41851, n41850, n51349, n51347, n6_adj_4209, 
        n51315;
    
    SB_DFFESR r_Clock_Count_2063__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n29244), 
            .D(n37[7]), .R(n29448));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n29244), 
            .D(n37[6]), .R(n29448));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n29244), 
            .D(n37[5]), .R(n29448));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n29244), 
            .D(n37[4]), .R(n29448));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n29244), 
            .D(n37[3]), .R(n29448));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n29244), 
            .D(n37[2]), .R(n29448));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n29244), 
            .D(n37[1]), .R(n29448));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n29244), 
            .D(n37[0]), .R(n29448));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n29175), 
            .D(n326[1]), .R(n29416));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n29175), 
            .D(n326[2]), .R(n29416));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3545[0]), .O(n29416));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_866 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_3542[2] ), .O(n29175));
    defparam i1_3_lut_4_lut_adj_866.LUT_INIT = 16'h1101;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3542[2] ), .O(n27775));
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut (.I0(n27775), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n27903));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_312_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_312_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n36314), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3548[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n36198), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2178_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i2178_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n45526));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i22735_2_lut (.I0(n45526), .I1(\r_SM_Main_2__N_3542[2] ), .I2(GND_net), 
            .I3(GND_net), .O(r_SM_Main_2__N_3545[0]));
    defparam i22735_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2171_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i2171_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n29587));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n29582));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n45179));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i4_4_lut (.I0(n9), .I1(n27763), .I2(r_Clock_Count[3]), .I3(r_Clock_Count[1]), 
            .O(r_SM_Main_2__N_3548[0]));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i3_4_lut_adj_867 (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(r_Clock_Count[5]), .O(n27763));   // verilog/uart_rx.v(118[17:47])
    defparam i3_4_lut_adj_867.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n29561));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n29560));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n29559));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n29558));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n29557));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n29556));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n29555));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n45591));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i22511_4_lut (.I0(r_Clock_Count[0]), .I1(n27763), .I2(n6), 
            .I3(r_Clock_Count[1]), .O(\r_SM_Main_2__N_3542[2] ));
    defparam i22511_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i3_2_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(GND_net), .O(n9));
    defparam i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 r_Clock_Count_2063_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n41856), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2063_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n41855), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_8 (.CI(n41855), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n41856));
    SB_LUT4 r_Clock_Count_2063_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n41854), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_7 (.CI(n41854), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n41855));
    SB_LUT4 r_Clock_Count_2063_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n41853), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_6 (.CI(n41853), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n41854));
    SB_LUT4 r_Clock_Count_2063_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n41852), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_5 (.CI(n41852), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n41853));
    SB_LUT4 r_Clock_Count_2063_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n41851), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_4 (.CI(n41851), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n41852));
    SB_LUT4 r_Clock_Count_2063_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n41850), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_3 (.CI(n41850), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n41851));
    SB_LUT4 r_Clock_Count_2063_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n41850));
    SB_LUT4 i36077_4_lut (.I0(r_Rx_Data), .I1(r_Clock_Count[1]), .I2(n27763), 
            .I3(r_Clock_Count[3]), .O(n51349));
    defparam i36077_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i36096_3_lut (.I0(n51349), .I1(r_SM_Main[0]), .I2(n9), .I3(GND_net), 
            .O(n51347));
    defparam i36096_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n51347), .I2(\r_SM_Main_2__N_3542[2] ), 
            .I3(r_SM_Main[1]), .O(n29448));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2_2_lut_adj_868 (.I0(r_SM_Main_2__N_3548[0]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4209));
    defparam i2_2_lut_adj_868.LUT_INIT = 16'h4444;
    SB_LUT4 i36857_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6_adj_4209), 
            .I3(r_Rx_Data), .O(n29244));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i36857_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 equal_310_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_8));   // verilog/uart_rx.v(97[17:39])
    defparam equal_310_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_308_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_9));   // verilog/uart_rx.v(97[17:39])
    defparam equal_308_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_869 (.I0(n27775), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n27898));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_869.LUT_INIT = 16'hbbbb;
    SB_LUT4 i21994_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35507));
    defparam i21994_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35923_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3548[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n51315));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i35923_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n51315), .I1(\r_SM_Main_2__N_3542[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n36314));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_3_lut (.I0(n45526), .I1(\r_SM_Main_2__N_3542[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n36198));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_3_lut.LUT_INIT = 16'hc7c7;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (CLK_c, enable_slow_N_4190, \state[1] , n5740, \state[0] , 
            GND_net, \state[3] , \state[0]_adj_4 , read, \state[2] , 
            n29575, rw, n45289, data_ready, n6387, sda_enable, \state_7__N_4087[0] , 
            n51345, n10, n27911, n27954, scl_enable, n29607, data, 
            n35513, n4, n29598, n29597, n29596, n29595, VCC_net, 
            \state_7__N_4103[3] , n6935, \saved_addr[0] , n10_adj_5, 
            n10_adj_6, n8, scl, n30125, sda_out, n29583, n29563, 
            n29538, n4_adj_7) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input CLK_c;
    output enable_slow_N_4190;
    output \state[1] ;
    output [0:0]n5740;
    output \state[0] ;
    input GND_net;
    output \state[3] ;
    output \state[0]_adj_4 ;
    input read;
    output \state[2] ;
    input n29575;
    output rw;
    input n45289;
    output data_ready;
    output n6387;
    output sda_enable;
    output \state_7__N_4087[0] ;
    output n51345;
    output n10;
    output n27911;
    output n27954;
    output scl_enable;
    input n29607;
    output [7:0]data;
    output n35513;
    output n4;
    input n29598;
    input n29597;
    input n29596;
    input n29595;
    input VCC_net;
    input \state_7__N_4103[3] ;
    input n6935;
    output \saved_addr[0] ;
    input n10_adj_5;
    output n10_adj_6;
    input n8;
    output scl;
    input n30125;
    output sda_out;
    input n29583;
    input n29563;
    input n29538;
    output n4_adj_7;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [15:0]delay_counter_15__N_3989;
    
    wire n29213;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    
    wire n29431, n42412, n15, n51340, enable, n7, n27773, n47167, 
        n13, n45151;
    wire [15:0]n4132;
    
    wire n28, n26, n27, n25, n40572, n40571, n40570, n40569, 
        n40568, n40567, n40566, n40565, n40564, n40563;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n40562, n40561, n40560, n40559, n40558, n45153;
    
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[1]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[2]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[3]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[4]), .S(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[5]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[6]), .S(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[7]), .S(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[8]), .S(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[9]), .S(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[10]), .S(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[11]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[12]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[13]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[14]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[15]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i35976_4_lut (.I0(n42412), .I1(enable_slow_N_4190), .I2(\state[1] ), 
            .I3(n15), .O(n51340));   // verilog/eeprom.v(23[11:16])
    defparam i35976_4_lut.LUT_INIT = 16'hfaee;
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n5740[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 state_7__I_0_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/eeprom.v(51[5:9])
    defparam state_7__I_0_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut (.I0(n7), .I1(\state[3] ), .I2(\state[0]_adj_4 ), 
            .I3(n27773), .O(n42412));   // verilog/eeprom.v(42[12:28])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(n15), .I1(n47167), .I2(enable_slow_N_4190), 
            .I3(n13), .O(n45151));   // verilog/coms.v(145[4] 299[11])
    defparam i1_4_lut.LUT_INIT = 16'hfac8;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n29213), 
            .D(delay_counter_15__N_3989[0]), .R(n29431));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i36898_2_lut (.I0(n27773), .I1(enable_slow_N_4190), .I2(GND_net), 
            .I3(GND_net), .O(n4132[14]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i36898_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n27773));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1366_Mux_0_i1_4_lut (.I0(read), .I1(n27773), .I2(\state[0] ), 
            .I3(enable_slow_N_4190), .O(n5740[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_1366_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 add_908_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n4132[14]), 
            .I3(n40572), .O(delay_counter_15__N_3989[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_908_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n4132[14]), 
            .I3(n40571), .O(delay_counter_15__N_3989[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_16 (.CI(n40571), .I0(delay_counter[14]), .I1(n4132[14]), 
            .CO(n40572));
    SB_LUT4 add_908_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n4132[14]), 
            .I3(n40570), .O(delay_counter_15__N_3989[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_15 (.CI(n40570), .I0(delay_counter[13]), .I1(n4132[14]), 
            .CO(n40571));
    SB_LUT4 add_908_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n4132[14]), 
            .I3(n40569), .O(delay_counter_15__N_3989[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_14 (.CI(n40569), .I0(delay_counter[12]), .I1(n4132[14]), 
            .CO(n40570));
    SB_LUT4 add_908_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n4132[14]), 
            .I3(n40568), .O(delay_counter_15__N_3989[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_13 (.CI(n40568), .I0(delay_counter[11]), .I1(n4132[14]), 
            .CO(n40569));
    SB_LUT4 add_908_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n4132[14]), 
            .I3(n40567), .O(delay_counter_15__N_3989[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_12 (.CI(n40567), .I0(delay_counter[10]), .I1(n4132[14]), 
            .CO(n40568));
    SB_LUT4 add_908_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n4132[14]), 
            .I3(n40566), .O(delay_counter_15__N_3989[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_11 (.CI(n40566), .I0(delay_counter[9]), .I1(n4132[14]), 
            .CO(n40567));
    SB_LUT4 add_908_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n4132[14]), 
            .I3(n40565), .O(delay_counter_15__N_3989[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_10 (.CI(n40565), .I0(delay_counter[8]), .I1(n4132[14]), 
            .CO(n40566));
    SB_LUT4 add_908_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n4132[14]), 
            .I3(n40564), .O(delay_counter_15__N_3989[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_9 (.CI(n40564), .I0(delay_counter[7]), .I1(n4132[14]), 
            .CO(n40565));
    SB_LUT4 add_908_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n4132[14]), 
            .I3(n40563), .O(delay_counter_15__N_3989[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(\state[2] ), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_908_8 (.CI(n40563), .I0(delay_counter[6]), .I1(n4132[14]), 
            .CO(n40564));
    SB_LUT4 add_908_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n4132[14]), 
            .I3(n40562), .O(delay_counter_15__N_3989[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_7 (.CI(n40562), .I0(delay_counter[5]), .I1(n4132[14]), 
            .CO(n40563));
    SB_LUT4 add_908_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n4132[14]), 
            .I3(n40561), .O(delay_counter_15__N_3989[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_6 (.CI(n40561), .I0(delay_counter[4]), .I1(n4132[14]), 
            .CO(n40562));
    SB_LUT4 add_908_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n4132[14]), 
            .I3(n40560), .O(delay_counter_15__N_3989[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_5 (.CI(n40560), .I0(delay_counter[3]), .I1(n4132[14]), 
            .CO(n40561));
    SB_LUT4 add_908_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n4132[14]), 
            .I3(n40559), .O(delay_counter_15__N_3989[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_4 (.CI(n40559), .I0(delay_counter[2]), .I1(n4132[14]), 
            .CO(n40560));
    SB_LUT4 add_908_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n4132[14]), 
            .I3(n40558), .O(delay_counter_15__N_3989[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_3 (.CI(n40558), .I0(delay_counter[1]), .I1(n4132[14]), 
            .CO(n40559));
    SB_LUT4 add_908_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n4132[14]), 
            .I3(GND_net), .O(delay_counter_15__N_3989[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n4132[14]), 
            .CO(n40558));
    SB_LUT4 i15922_2_lut (.I0(n29213), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29431));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15922_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n29213));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n45151));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n45153));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n29575));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n45289));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i24_4_lut_4_lut (.I0(\state[1] ), .I1(read), .I2(\state[0] ), 
            .I3(n51340), .O(n45153));   // verilog/eeprom.v(23[11:16])
    defparam i24_4_lut_4_lut.LUT_INIT = 16'hf404;
    SB_LUT4 i2_4_lut_4_lut (.I0(n42412), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(GND_net), .O(n47167));   // verilog/coms.v(145[4] 299[11])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[1] ), .I1(enable_slow_N_4190), .I2(read), 
            .I3(\state[0] ), .O(n13));   // verilog/coms.v(145[4] 299[11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'haa8a;
    i2c_controller i2c (.CLK_c(CLK_c), .n6387(n6387), .\state[1] (state[1]), 
            .\state[2] (\state[2] ), .\state[3] (\state[3] ), .sda_enable(sda_enable), 
            .enable_slow_N_4190(enable_slow_N_4190), .\state_7__N_4087[0] (\state_7__N_4087[0] ), 
            .n51345(n51345), .\state[0] (\state[0]_adj_4 ), .GND_net(GND_net), 
            .n10(n10), .n27911(n27911), .n27954(n27954), .scl_enable(scl_enable), 
            .n29607(n29607), .data({data}), .n35513(n35513), .n4(n4), 
            .n29598(n29598), .n29597(n29597), .n29596(n29596), .n29595(n29595), 
            .VCC_net(VCC_net), .\state_7__N_4103[3] (\state_7__N_4103[3] ), 
            .n6935(n6935), .\saved_addr[0] (\saved_addr[0] ), .n10_adj_1(n10_adj_5), 
            .enable(enable), .n10_adj_2(n10_adj_6), .n8(n8), .scl(scl), 
            .n30125(n30125), .sda_out(sda_out), .n29583(n29583), .n29563(n29563), 
            .n29538(n29538), .n4_adj_3(n4_adj_7)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (CLK_c, n6387, \state[1] , \state[2] , \state[3] , 
            sda_enable, enable_slow_N_4190, \state_7__N_4087[0] , n51345, 
            \state[0] , GND_net, n10, n27911, n27954, scl_enable, 
            n29607, data, n35513, n4, n29598, n29597, n29596, 
            n29595, VCC_net, \state_7__N_4103[3] , n6935, \saved_addr[0] , 
            n10_adj_1, enable, n10_adj_2, n8, scl, n30125, sda_out, 
            n29583, n29563, n29538, n4_adj_3) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input CLK_c;
    output n6387;
    output \state[1] ;
    output \state[2] ;
    output \state[3] ;
    output sda_enable;
    output enable_slow_N_4190;
    output \state_7__N_4087[0] ;
    output n51345;
    output \state[0] ;
    input GND_net;
    output n10;
    output n27911;
    output n27954;
    output scl_enable;
    input n29607;
    output [7:0]data;
    output n35513;
    output n4;
    input n29598;
    input n29597;
    input n29596;
    input n29595;
    input VCC_net;
    input \state_7__N_4103[3] ;
    input n6935;
    output \saved_addr[0] ;
    input n10_adj_1;
    input enable;
    output n10_adj_2;
    input n8;
    output scl;
    input n30125;
    output sda_out;
    input n29583;
    input n29563;
    input n29538;
    output n4_adj_3;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n29451, n5, n35595, n35650, n36202, n45353, n47752, n20040, 
        n6809, n29404;
    wire [0:0]n6094;
    
    wire n45223, sda_out_adj_4194;
    wire [7:0]n119;
    
    wire n29287;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n29486, n11, n11_adj_4195, n17, enable_slow_N_4189, i2c_clk_N_4176, 
        n29041, n9, scl_enable_N_4177, n29160, n6058, n40748, n40747, 
        n40746, n40745, n40744, n40743, n40742, n46494, n6380, 
        n37, n51319, n51272, n33, n34, n39, n7, n51375, n11_adj_4197, 
        n12, n35305, n11_adj_4199, n10_adj_4200, n41900, n41899, 
        n41898, n41897, n41896;
    
    SB_DFFSR counter2_2067_2068__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n29451));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6387), .D(n5), 
            .S(n35595));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6387), .D(n35650), 
            .S(n36202));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6387), .D(n45353), 
            .S(n47752));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n6809), 
            .D(n20040), .S(n29404));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4194), .C(i2c_clk), .E(n45223), 
            .D(n6094[0]));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n29287), .D(n119[0]), 
            .S(n29486));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i35958_3_lut_4_lut (.I0(n11), .I1(n11_adj_4195), .I2(enable_slow_N_4190), 
            .I3(\state_7__N_4087[0] ), .O(n51345));
    defparam i35958_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 i36984_3_lut_4_lut (.I0(n11), .I1(n11_adj_4195), .I2(n17), 
            .I3(n6387), .O(n35595));
    defparam i36984_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11_adj_4195));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i36880_2_lut (.I0(\state_7__N_4087[0] ), .I1(enable_slow_N_4190), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4189));   // verilog/i2c_controller.v(62[6:32])
    defparam i36880_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n29451), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4176));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n29041));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i36936_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11_adj_4195), 
            .I3(n6387), .O(n36202));   // verilog/i2c_controller.v(151[5:14])
    defparam i36936_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n29287), .D(n119[3]), 
            .R(n29486));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10), .I2(counter[0]), .I3(GND_net), 
            .O(n27911));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n29287), .D(n119[2]), 
            .S(n29486));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_3_lut_adj_860 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n27954));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_860.LUT_INIT = 16'hefef;
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_4176));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4177));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_120 (.Q(\state_7__N_4087[0] ), .C(CLK_c), .E(n29160), 
            .D(enable_slow_N_4189));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n29287), .D(n119[1]), 
            .S(n29486));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_3_lut_4_lut_adj_861 (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(n17), .O(scl_enable_N_4177));
    defparam i1_3_lut_4_lut_adj_861.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_4_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[3] ), 
            .I3(\state[2] ), .O(n6058));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h001c;
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29607));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i22000_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35513));
    defparam i22000_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_316_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_316_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29598));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29597));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29596));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29595));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n40748), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n40747), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n40747), .I0(counter[6]), .I1(VCC_net), 
            .CO(n40748));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n40746), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n40746), .I0(counter[5]), .I1(VCC_net), 
            .CO(n40747));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n40745), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n40745), .I0(counter[4]), .I1(VCC_net), 
            .CO(n40746));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n40744), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n40744), .I0(counter[3]), .I1(VCC_net), 
            .CO(n40745));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n40743), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n40743), .I0(counter[2]), .I1(VCC_net), 
            .CO(n40744));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n40742), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31130_2_lut (.I0(\state_7__N_4103[3] ), .I1(n17), .I2(GND_net), 
            .I3(GND_net), .O(n46494));
    defparam i31130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(n6380), .I1(n46494), .I2(n6935), .I3(n37), 
            .O(n29287));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i35904_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n51319));   // verilog/i2c_controller.v(198[28:35])
    defparam i35904_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i35916_4_lut (.I0(n51319), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n51272));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i35916_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 mux_1503_i1_4_lut (.I0(n51272), .I1(\state[0] ), .I2(n6058), 
            .I3(\state[2] ), .O(n6094[0]));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam mux_1503_i1_4_lut.LUT_INIT = 16'h303a;
    SB_CARRY sub_39_add_2_3 (.CI(n40742), .I0(counter[1]), .I1(VCC_net), 
            .CO(n40743));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n40742));
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33), .I2(n37), .I3(GND_net), 
            .O(n29404));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_862 (.I0(n34), .I1(n37), .I2(GND_net), .I3(GND_net), 
            .O(n39));
    defparam i1_2_lut_adj_862.LUT_INIT = 16'heeee;
    SB_LUT4 i36910_4_lut (.I0(n6058), .I1(n39), .I2(\state[2] ), .I3(\state[1] ), 
            .O(n6809));
    defparam i36910_4_lut.LUT_INIT = 16'hc8cc;
    SB_LUT4 i36874_2_lut (.I0(\state[0] ), .I1(n6058), .I2(GND_net), .I3(GND_net), 
            .O(n20040));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i36874_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_863 (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_863.LUT_INIT = 16'h4444;
    SB_LUT4 i36051_4_lut (.I0(n10_adj_1), .I1(n10), .I2(\state_7__N_4103[3] ), 
            .I3(enable), .O(n51375));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i36051_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(n7), .I2(n51375), .I3(\state[0] ), 
            .O(n45353));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i36992_2_lut (.I0(\state_7__N_4103[3] ), .I1(n11_adj_4197), 
            .I2(GND_net), .I3(GND_net), .O(n35650));
    defparam i36992_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_2));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10_adj_2), 
            .O(n6380));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i36872_4_lut (.I0(n29041), .I1(n6380), .I2(n11), .I3(n35305), 
            .O(n6387));
    defparam i36872_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_864 (.I0(n11_adj_4199), .I1(n11_adj_4197), .I2(\state_7__N_4103[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_864.LUT_INIT = 16'h5755;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i21907_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i21907_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4200));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4200), .I2(counter2[0]), 
            .I3(GND_net), .O(n29451));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n30125));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i2367_2_lut (.I0(sda_out_adj_4194), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2367_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n29287), .D(n119[7]), 
            .R(n29486));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n29287), .D(n119[6]), 
            .R(n29486));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n29287), .D(n119[5]), 
            .R(n29486));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n29287), .D(n119[4]), 
            .R(n29486));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29583));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n29563));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2067_2068__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n29451));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2067_2068__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n29451));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2067_2068__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n29451));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2067_2068__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n29451));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2067_2068__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n29451));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29538));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 counter2_2067_2068_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n41900), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2067_2068_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n41899), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_6 (.CI(n41899), .I0(GND_net), .I1(counter2[4]), 
            .CO(n41900));
    SB_LUT4 counter2_2067_2068_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n41898), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_5 (.CI(n41898), .I0(GND_net), .I1(counter2[3]), 
            .CO(n41899));
    SB_LUT4 counter2_2067_2068_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n41897), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_4 (.CI(n41897), .I0(GND_net), .I1(counter2[2]), 
            .CO(n41898));
    SB_LUT4 counter2_2067_2068_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n41896), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_3 (.CI(n41896), .I0(GND_net), .I1(counter2[1]), 
            .CO(n41897));
    SB_LUT4 counter2_2067_2068_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n41896));
    SB_LUT4 equal_318_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_318_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i21803_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n35305));
    defparam i21803_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i36934_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n6387), .O(n47752));
    defparam i36934_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0554;
    SB_LUT4 i31098_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n46494), .O(n29486));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i31098_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 equal_2051_i19_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4190));
    defparam equal_2051_i19_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4197));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n17));   // verilog/i2c_controller.v(77[27:43])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4199));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i36908_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n45223));
    defparam i36908_4_lut_4_lut.LUT_INIT = 16'h0156;
    SB_LUT4 i1_2_lut_3_lut_adj_865 (.I0(enable), .I1(\state_7__N_4087[0] ), 
            .I2(enable_slow_N_4190), .I3(GND_net), .O(n29160));
    defparam i1_2_lut_3_lut_adj_865.LUT_INIT = 16'heaea;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000) 
//

module \quadrature_decoder(1,500000)  (encoder1_position, GND_net, \a_new[1] , 
            ENCODER1_B_N_keep, n1653, ENCODER1_A_N_keep, VCC_net, b_prev, 
            direction_N_3907, n29591, n1658) /* synthesis lattice_noprune=1 */ ;
    output [31:0]encoder1_position;
    input GND_net;
    output \a_new[1] ;
    input ENCODER1_B_N_keep;
    input n1653;
    input ENCODER1_A_N_keep;
    input VCC_net;
    output b_prev;
    output direction_N_3907;
    input n29591;
    output n1658;
    
    wire [31:0]n133;
    
    wire direction_N_3906, n41844, n41845, n41843, n41842, n41841, 
        n41840, n41839, n41838, n41837, n41836, n41835, n41834;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire a_prev_N_3913, n41833, n41832, n41831, n41830, n41829, 
        n41828, n41827, n41826, n41825, n41824, n41823, n41822, 
        n41821, n41820, n41819, debounce_cnt, n29599, a_prev, n29588, 
        direction_N_3910, n41849, n41848, n41847, n41846;
    
    SB_LUT4 position_2061_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[26]), .I3(n41844), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_28 (.CI(n41844), .I0(direction_N_3906), 
            .I1(encoder1_position[26]), .CO(n41845));
    SB_LUT4 position_2061_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[25]), .I3(n41843), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_27 (.CI(n41843), .I0(direction_N_3906), 
            .I1(encoder1_position[25]), .CO(n41844));
    SB_LUT4 position_2061_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[24]), .I3(n41842), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_26 (.CI(n41842), .I0(direction_N_3906), 
            .I1(encoder1_position[24]), .CO(n41843));
    SB_LUT4 position_2061_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[23]), .I3(n41841), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_25 (.CI(n41841), .I0(direction_N_3906), 
            .I1(encoder1_position[23]), .CO(n41842));
    SB_LUT4 position_2061_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[22]), .I3(n41840), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_24 (.CI(n41840), .I0(direction_N_3906), 
            .I1(encoder1_position[22]), .CO(n41841));
    SB_LUT4 position_2061_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[21]), .I3(n41839), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_23 (.CI(n41839), .I0(direction_N_3906), 
            .I1(encoder1_position[21]), .CO(n41840));
    SB_LUT4 position_2061_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[20]), .I3(n41838), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_22 (.CI(n41838), .I0(direction_N_3906), 
            .I1(encoder1_position[20]), .CO(n41839));
    SB_LUT4 position_2061_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[19]), .I3(n41837), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_21 (.CI(n41837), .I0(direction_N_3906), 
            .I1(encoder1_position[19]), .CO(n41838));
    SB_LUT4 position_2061_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[18]), .I3(n41836), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_20 (.CI(n41836), .I0(direction_N_3906), 
            .I1(encoder1_position[18]), .CO(n41837));
    SB_LUT4 position_2061_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[17]), .I3(n41835), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_19 (.CI(n41835), .I0(direction_N_3906), 
            .I1(encoder1_position[17]), .CO(n41836));
    SB_LUT4 position_2061_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[16]), .I3(n41834), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_18 (.CI(n41834), .I0(direction_N_3906), 
            .I1(encoder1_position[16]), .CO(n41835));
    SB_LUT4 i36896_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i36896_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 position_2061_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[15]), .I3(n41833), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_17 (.CI(n41833), .I0(direction_N_3906), 
            .I1(encoder1_position[15]), .CO(n41834));
    SB_LUT4 position_2061_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[14]), .I3(n41832), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_16 (.CI(n41832), .I0(direction_N_3906), 
            .I1(encoder1_position[14]), .CO(n41833));
    SB_LUT4 position_2061_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[13]), .I3(n41831), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_15 (.CI(n41831), .I0(direction_N_3906), 
            .I1(encoder1_position[13]), .CO(n41832));
    SB_LUT4 position_2061_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[12]), .I3(n41830), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_14 (.CI(n41830), .I0(direction_N_3906), 
            .I1(encoder1_position[12]), .CO(n41831));
    SB_LUT4 position_2061_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[11]), .I3(n41829), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1653), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1653), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_CARRY position_2061_add_4_13 (.CI(n41829), .I0(direction_N_3906), 
            .I1(encoder1_position[11]), .CO(n41830));
    SB_LUT4 position_2061_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[10]), .I3(n41828), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_12 (.CI(n41828), .I0(direction_N_3906), 
            .I1(encoder1_position[10]), .CO(n41829));
    SB_LUT4 position_2061_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[9]), .I3(n41827), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_11 (.CI(n41827), .I0(direction_N_3906), 
            .I1(encoder1_position[9]), .CO(n41828));
    SB_LUT4 position_2061_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[8]), .I3(n41826), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_10 (.CI(n41826), .I0(direction_N_3906), 
            .I1(encoder1_position[8]), .CO(n41827));
    SB_LUT4 position_2061_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[7]), .I3(n41825), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_9 (.CI(n41825), .I0(direction_N_3906), 
            .I1(encoder1_position[7]), .CO(n41826));
    SB_LUT4 position_2061_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[6]), .I3(n41824), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_8 (.CI(n41824), .I0(direction_N_3906), 
            .I1(encoder1_position[6]), .CO(n41825));
    SB_LUT4 position_2061_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[5]), .I3(n41823), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_7 (.CI(n41823), .I0(direction_N_3906), 
            .I1(encoder1_position[5]), .CO(n41824));
    SB_LUT4 position_2061_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[4]), .I3(n41822), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_6 (.CI(n41822), .I0(direction_N_3906), 
            .I1(encoder1_position[4]), .CO(n41823));
    SB_LUT4 position_2061_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[3]), .I3(n41821), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_5 (.CI(n41821), .I0(direction_N_3906), 
            .I1(encoder1_position[3]), .CO(n41822));
    SB_LUT4 position_2061_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[2]), .I3(n41820), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_4 (.CI(n41820), .I0(direction_N_3906), 
            .I1(encoder1_position[2]), .CO(n41821));
    SB_LUT4 position_2061_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[1]), .I3(n41819), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_3 (.CI(n41819), .I0(direction_N_3906), 
            .I1(encoder1_position[1]), .CO(n41820));
    SB_LUT4 position_2061_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n41819));
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1653), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1653), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1653), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 i16077_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n29599));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16077_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16066_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n29588));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE position_2061__i0 (.Q(encoder1_position[0]), .C(n1653), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1653), .D(n29599));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1658), .C(n1653), .D(n29591));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(\a_new[1] ), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1653), .D(n29588));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2061__i1 (.Q(encoder1_position[1]), .C(n1653), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i2 (.Q(encoder1_position[2]), .C(n1653), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i3 (.Q(encoder1_position[3]), .C(n1653), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i4 (.Q(encoder1_position[4]), .C(n1653), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i5 (.Q(encoder1_position[5]), .C(n1653), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i6 (.Q(encoder1_position[6]), .C(n1653), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i7 (.Q(encoder1_position[7]), .C(n1653), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i8 (.Q(encoder1_position[8]), .C(n1653), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i9 (.Q(encoder1_position[9]), .C(n1653), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i10 (.Q(encoder1_position[10]), .C(n1653), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i11 (.Q(encoder1_position[11]), .C(n1653), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i12 (.Q(encoder1_position[12]), .C(n1653), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i13 (.Q(encoder1_position[13]), .C(n1653), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i14 (.Q(encoder1_position[14]), .C(n1653), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i15 (.Q(encoder1_position[15]), .C(n1653), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i16 (.Q(encoder1_position[16]), .C(n1653), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i17 (.Q(encoder1_position[17]), .C(n1653), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i18 (.Q(encoder1_position[18]), .C(n1653), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i19 (.Q(encoder1_position[19]), .C(n1653), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i20 (.Q(encoder1_position[20]), .C(n1653), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i21 (.Q(encoder1_position[21]), .C(n1653), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i22 (.Q(encoder1_position[22]), .C(n1653), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i23 (.Q(encoder1_position[23]), .C(n1653), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i24 (.Q(encoder1_position[24]), .C(n1653), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i25 (.Q(encoder1_position[25]), .C(n1653), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i26 (.Q(encoder1_position[26]), .C(n1653), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i27 (.Q(encoder1_position[27]), .C(n1653), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i28 (.Q(encoder1_position[28]), .C(n1653), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i29 (.Q(encoder1_position[29]), .C(n1653), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i30 (.Q(encoder1_position[30]), .C(n1653), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i31 (.Q(encoder1_position[31]), .C(n1653), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 position_2061_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[31]), .I3(n41849), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2061_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[30]), .I3(n41848), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_32 (.CI(n41848), .I0(direction_N_3906), 
            .I1(encoder1_position[30]), .CO(n41849));
    SB_LUT4 position_2061_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[29]), .I3(n41847), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_31 (.CI(n41847), .I0(direction_N_3906), 
            .I1(encoder1_position[29]), .CO(n41848));
    SB_LUT4 position_2061_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[28]), .I3(n41846), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_30 (.CI(n41846), .I0(direction_N_3906), 
            .I1(encoder1_position[28]), .CO(n41847));
    SB_LUT4 position_2061_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[27]), .I3(n41845), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_29 (.CI(n41845), .I0(direction_N_3906), 
            .I1(encoder1_position[27]), .CO(n41846));
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (pwm_setpoint, GND_net, pwm_out, clk32MHz, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input [23:0]pwm_setpoint;
    input GND_net;
    output pwm_out;
    input clk32MHz;
    input VCC_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n24, n8, n45, n51435, n52105, n52034, n25, n51762;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n4, pwm_out_N_797, n27, n52031, n29, n52032, n33, n31, 
        n51459, n51454, n30, n10, n35, n51450, n52284, n51764, 
        n52312, n37, n52313, n39, n52307, n43, n41, n52255, 
        n51443, n51438, n52199, n40, n52201;
    wire [23:0]n101;
    
    wire n41809, n41808, n41807, n41806, n41805, n41804, n41803, 
        n41802, n41801, n41800, n41799, n41798, n41797, n41796, 
        n41795, n41794, n41793, n41792, n41791, n41790, n41789, 
        n41788, n41787, pwm_counter_23__N_795, n48043, n6, n48066, 
        n14, n13, n15, n51514, n6_adj_4191, n23, n11, n13_adj_4192, 
        n15_adj_4193, n9, n17, n19, n21, n51480, n12, n51814, 
        n51810, n52211, n51989, n52033, n16;
    
    SB_LUT4 i36622_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n51435), 
            .O(n52105));   // verilog/pwm.v(21[8:24])
    defparam i36622_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36280_3_lut (.I0(n52034), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n51762));   // verilog/pwm.v(21[8:24])
    defparam i36280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_DFF pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .D(pwm_out_N_797));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i36548_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n52031));   // verilog/pwm.v(21[8:24])
    defparam i36548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36549_3_lut (.I0(n52031), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n52032));   // verilog/pwm.v(21[8:24])
    defparam i36549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35972_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n51459), 
            .O(n51454));
    defparam i35972_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36801_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n51450), 
            .O(n52284));   // verilog/pwm.v(21[8:24])
    defparam i36801_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36282_3_lut (.I0(n52032), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n51764));   // verilog/pwm.v(21[8:24])
    defparam i36282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36829_4_lut (.I0(n51764), .I1(n52284), .I2(n35), .I3(n51454), 
            .O(n52312));   // verilog/pwm.v(21[8:24])
    defparam i36829_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36830_3_lut (.I0(n52312), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n52313));   // verilog/pwm.v(21[8:24])
    defparam i36830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36824_3_lut (.I0(n52313), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n52307));   // verilog/pwm.v(21[8:24])
    defparam i36824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35961_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n52255), 
            .O(n51443));
    defparam i35961_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36716_4_lut (.I0(n51762), .I1(n52105), .I2(n45), .I3(n51438), 
            .O(n52199));   // verilog/pwm.v(21[8:24])
    defparam i36716_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36806_3_lut (.I0(n52307), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n40));   // verilog/pwm.v(21[8:24])
    defparam i36806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36718_4_lut (.I0(n40), .I1(n52199), .I2(n45), .I3(n51443), 
            .O(n52201));   // verilog/pwm.v(21[8:24])
    defparam i36718_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36719_3_lut (.I0(n52201), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_797));   // verilog/pwm.v(21[8:24])
    defparam i36719_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 pwm_counter_2059_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n41809), .O(n101[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_2059_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n41808), .O(n101[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_24 (.CI(n41808), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n41809));
    SB_LUT4 pwm_counter_2059_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n41807), .O(n101[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_23 (.CI(n41807), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n41808));
    SB_LUT4 pwm_counter_2059_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n41806), .O(n101[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_22 (.CI(n41806), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n41807));
    SB_LUT4 pwm_counter_2059_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n41805), .O(n101[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_21 (.CI(n41805), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n41806));
    SB_LUT4 pwm_counter_2059_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n41804), .O(n101[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_20 (.CI(n41804), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n41805));
    SB_LUT4 pwm_counter_2059_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n41803), .O(n101[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_19 (.CI(n41803), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n41804));
    SB_LUT4 pwm_counter_2059_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n41802), .O(n101[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_18 (.CI(n41802), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n41803));
    SB_LUT4 pwm_counter_2059_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n41801), .O(n101[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_17 (.CI(n41801), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n41802));
    SB_LUT4 pwm_counter_2059_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n41800), .O(n101[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_16 (.CI(n41800), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n41801));
    SB_LUT4 pwm_counter_2059_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n41799), .O(n101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_15 (.CI(n41799), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n41800));
    SB_LUT4 pwm_counter_2059_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n41798), .O(n101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_14 (.CI(n41798), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n41799));
    SB_LUT4 pwm_counter_2059_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n41797), .O(n101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_13 (.CI(n41797), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n41798));
    SB_LUT4 pwm_counter_2059_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n41796), .O(n101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_12 (.CI(n41796), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n41797));
    SB_LUT4 pwm_counter_2059_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n41795), .O(n101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_11 (.CI(n41795), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n41796));
    SB_LUT4 pwm_counter_2059_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n41794), .O(n101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_10 (.CI(n41794), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n41795));
    SB_LUT4 pwm_counter_2059_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n41793), .O(n101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_9 (.CI(n41793), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n41794));
    SB_LUT4 pwm_counter_2059_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n41792), .O(n101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_8 (.CI(n41792), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n41793));
    SB_LUT4 pwm_counter_2059_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n41791), .O(n101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_7 (.CI(n41791), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n41792));
    SB_LUT4 pwm_counter_2059_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n41790), .O(n101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_6 (.CI(n41790), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n41791));
    SB_LUT4 pwm_counter_2059_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n41789), .O(n101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_5 (.CI(n41789), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n41790));
    SB_LUT4 pwm_counter_2059_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n41788), .O(n101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_4 (.CI(n41788), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n41789));
    SB_LUT4 pwm_counter_2059_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n41787), .O(n101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_3 (.CI(n41787), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n41788));
    SB_LUT4 pwm_counter_2059_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n41787));
    SB_DFFSR pwm_counter_2059__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n101[0]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n48043));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[21]), .I1(n48043), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n6));
    defparam i1_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut (.I0(pwm_counter[12]), .I1(pwm_counter[13]), .I2(pwm_counter[20]), 
            .I3(n6), .O(n48066));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(pwm_counter[17]), .I1(n48066), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_2_lut (.I0(pwm_counter[19]), .I1(pwm_counter[14]), .I2(GND_net), 
            .I3(GND_net), .O(n13));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[22]), .I1(pwm_counter[16]), .I2(pwm_counter[18]), 
            .I3(pwm_counter[15]), .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37610_4_lut (.I0(pwm_counter[23]), .I1(n15), .I2(n13), .I3(n14), 
            .O(pwm_counter_23__N_795));   // verilog/pwm.v(18[8:40])
    defparam i37610_4_lut.LUT_INIT = 16'h5554;
    SB_DFFSR pwm_counter_2059__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n101[1]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n101[2]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n101[3]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n101[4]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n101[5]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n101[6]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n101[7]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n101[8]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n101[9]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n101[10]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n101[11]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n101[12]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n101[13]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n101[14]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n101[15]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n101[16]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n101[17]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n101[18]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n101[19]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n101[20]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n101[21]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n101[22]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n101[23]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i36032_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n51514));   // verilog/pwm.v(21[8:24])
    defparam i36032_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6_adj_4191));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4192));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4193));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35998_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n51480));
    defparam i35998_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35977_4_lut (.I0(n27), .I1(n15_adj_4193), .I2(n13_adj_4192), 
            .I3(n11), .O(n51459));
    defparam i35977_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36332_4_lut (.I0(n13_adj_4192), .I1(n11), .I2(n9), .I3(n51514), 
            .O(n51814));
    defparam i36332_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36328_4_lut (.I0(n19), .I1(n17), .I2(n15_adj_4193), .I3(n51814), 
            .O(n51810));
    defparam i36328_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36728_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n51810), 
            .O(n52211));
    defparam i36728_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36506_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n52211), 
            .O(n51989));
    defparam i36506_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36772_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n51989), 
            .O(n52255));
    defparam i36772_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36550_3_lut (.I0(n6_adj_4191), .I1(pwm_setpoint[10]), .I2(n21), 
            .I3(GND_net), .O(n52033));   // verilog/pwm.v(21[8:24])
    defparam i36550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36551_3_lut (.I0(n52033), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n52034));   // verilog/pwm.v(21[8:24])
    defparam i36551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35956_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n51480), 
            .O(n51438));
    defparam i35956_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35953_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n51435));
    defparam i35953_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35968_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n51450));
    defparam i35968_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
