// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Feb 26 21:17:16 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(48[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(94[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(95[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    
    wire n43615, n43614;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    
    wire n15;
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(280[22:33])
    
    wire n48672, n29428, n27281, n43613;
    wire [7:0]data;   // verilog/TinyFPGA_B.v(337[14:18])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(361[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(369[15:20])
    
    wire pwm_setpoint_23__N_263, n209, n211, n249, n250, n251, n252, 
        n253, n254, n255, n256, n257, n258, n259, n260, n261, 
        n262, n263, n264, n265, n266, n267, n268, n269, n270, 
        n296, n43612, n330, n334, n335, n336, n337, n338, n339, 
        n340, n341, n342, n343, n344, n345;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire n356, n56518, n56506, n56500, n379, n43611, n43610, n43160, 
        n418, n419, n420, n421, n422, n423, n424, n425, n426, 
        n427, n428, n429, n430, n431, n432, n433, n434, n435, 
        n436, n437, n438, n439, n440, n441;
    wire [23:0]pwm_setpoint_23__N_11;
    wire [7:0]commutation_state_7__N_264;
    
    wire commutation_state_7__N_272, n29426, n29425;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n29424, GHA_N_478, GLA_N_495, GHB_N_500, GLB_N_509, GHC_N_514, 
        GLC_N_523, dti_N_527, n43609, n29423, n29422, n29421, n29420, 
        n29419, n29418, RX_N_10;
    wire [31:0]motor_state_23__N_123;
    wire [31:0]encoder0_position_scaled_23__N_327;
    wire [32:0]encoder0_position_scaled_23__N_51;
    
    wire encoder1_position_scaled_23__N_359;
    wire [31:0]encoder1_position_scaled_23__N_75;
    wire [23:0]displacement_23__N_99;
    
    wire n2274, n8584, n8585, n8586, n8587, n1532, n1533, n1534, 
        n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
        n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, 
        n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
        n1559, n1560, n1561, n1562, n1563, n43608, n43607, n43606, 
        n43605, n8588, n8589, n1650, n43604, n43603, n43602, n43601, 
        n43600, n56362, n56356, n56350, n56344, n56338, n2091, 
        n2233;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n43599, n5, n36748, n43598, n43597, n43596;
    wire [3:0]state_3__N_639;
    
    wire n24, n20, n56458, n4, n8, n29417, n15_adj_5457, n7936, 
        n43595, n43594, n43593, n43592, n43591, n4929, n43590, 
        n5_adj_5458, n52732, n29416, n29415, n43589, n29411, n4928, 
        n4927, n43159, n20976, n43588, n43587, n43586, n43158, 
        n43585, n4926, n4925, n4924, n4923, n43584, n4922, n43583, 
        n4921, n4920, n4919, n4918, n4917, n4599, n4916, n4915, 
        n4914, n29410, n29409, n43156, n4_adj_5459, n55474, n625, 
        n623, n622, n621, n55375, n55333, n4913, n43582, n29408, 
        n29407, n29406, n29405, n29404, n29403, n55935, n43157, 
        n43581, n54784, n29402, n4748, n43580, n43104, n43579, 
        n43578, n43577, n3, n4_adj_5460, n5_adj_5461, n6, n7, 
        n8_adj_5462, n9, n10, n11, n12, n13, n14, n15_adj_5463, 
        n16, n17, n18, n19, n20_adj_5464, n21, n22, n23, n24_adj_5465, 
        n25, n2, n29401, n14_adj_5466, n15_adj_5467, n16_adj_5468, 
        n17_adj_5469, n18_adj_5470, n19_adj_5471, n20_adj_5472, n21_adj_5473, 
        n22_adj_5474, n23_adj_5475, n24_adj_5476, n25_adj_5477, n4_adj_5478, 
        n29400, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(92[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(96[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(96[12:19])
    
    wire n49469;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(97[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(98[12:26])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(113[11:16])
    
    wire n43576, n49781, n43088, n43575, n43574, n43573, n43572, 
        n43571, n4_adj_5479, n43570, n122, n43569, n43568, n43567, 
        n43566, n43565, n43564, n43563, n43562, n43561, n43560, 
        n43559, n43558, n43557, n43556, n43555, n43103, n43554, 
        n36740, n43553, n43087, n36736, n43552, n43102, n43551, 
        n4912, n4911, n43550, n43549, n43548, n43101, n43547, 
        n43546, n56702, n56452, n56700, n56446, n56440, n56410, 
        n43545, n43544, n43100, n43543, n43099, n43542, n43541, 
        n43540, n43539, n43538, n43537, n43536, n43993, n43535, 
        n43992, n43534, n4_adj_5480, n43991, n43533, n43990, n43532, 
        n43989, n43988, n43531, n43530, n43987, n43529, n43528, 
        n43986, n43985, n49436, n544, n543, n542, n541, n540, 
        n539, n538, n537, n536, n535, n534, n533, n532, n531, 
        n530, n529, n528, n527, n526, n525, n43527, n43526, 
        n43984, n43983, n43525, n43086, n43524, n43982, n43085, 
        n43098, n43981, n43523, n43084, n43522, n43521, n43980, 
        n43520, n43519, n43979, n43978, n43518, n43977, n43517, 
        n43516, n43976, n55263, n43975, n43515, n43514, n43974, 
        n43513, n43512, n43973, n43511, n43972, n43510, n55332, 
        n43509, n54780, n43971, n43970, n43508, n27117, n43969, 
        n43097, n43968, n43967, n43966, n43965, n43964, n43963, 
        n43962, n43961, n36728, n43960, n43959, n43500, n43958, 
        n43957, n43956, n43955, n43954, n43953, n43952, n36718, 
        n43951, n43499, n43950, n43498, n43949, n43948, n43947, 
        n49707, n43497, n43496, n43946, n43945, n43944, n43943, 
        n43942, n43495, n43941, n43940, n43939, n43938, n51094, 
        n36712, n36710, n43937, n43936, n43494, n43493, n43935, 
        n43934, n43933, n43932, n43083, n43492, n43931, n43930, 
        n43929, n36704, n43491, n54721, n43928, n43927, n43490, 
        n43926, n43925, n43924, n57092, n43923, n524, n29396, 
        n29395, n54718, n523, n522, n521, n43922, n29394, n520, 
        n519, n27222, n29393, n518, n516, n43489, n3303, n43488, 
        n43487, n43921, n50654, n43486, n36694, n43920, n43919, 
        n43918, n43917, n43485, n43916, n43484, n43483, n43915, 
        n43482, n43481, n49611, n43914, n43480, n43913, n43479, 
        n43912, n43911, n43478, n36672, n43910, n43909, n43908, 
        n43907, n43906, n43905, n54709, n36668, n36666, n36664, 
        n43124, n43904, n43903, n43902, n43123, n43901, n43468, 
        n43900, n43899, n43096, n43467, n43466, n43465, n43095, 
        n43898, n43897, n43464, n36660, n43463, n36658, n36510, 
        n36656, n43896, n43895, n43462, n43122, n43461, n43894, 
        n43460, n43893, n43892, n43891, n43459, n43458, n43890, 
        n43457, n43121, n36654, n43456, n49594, n36650, n36648, 
        n43889, n43455, n43094, n43888, n43887, n43454, n43453, 
        n43452, n43886, n43885, n43884, n43451, n43883, n43450, 
        n43449, n43882, n15_adj_5481, n54704, n29392, n29391, n51177, 
        n43881, n43448, n54702, n29390, n29389, n4452, n36642, 
        n36640, n49681, n43880, n43120, n43879, n43447, n43878, 
        n43446, n43877, n43445, n43876, n43119, n43082, n43875, 
        n43118, n43444, n36636, n43874, n36634, n36632, n43443, 
        n43873, n43872, n43871, n43870, n43869, n43868, n49501, 
        n43117, n5_adj_5482, n43442, n43867, n43866, n43865, n43864, 
        n36630, n43441, n43863, n43440, n43862, n43861, n43860, 
        n43859, n43858, n43857, n43856, n54692, n49689, n43855, 
        n43854, n43116, n43853, n43852, n43115, n43851, n43850, 
        n43849, n43848, n43114, n43847, n43846, n43845, n43844, 
        n43843, n49477, n43842, n43841, n49475, n49473, n35841, 
        n49471, n49468, n36626, n35837, n43840, n54688, n54686, 
        n43839, n43838, n43837, n43836, n43835, n43834, n43833, 
        n43832, n43831, n43830, n43829, n43828, n43827, n43439, 
        n43826, n43825, n43824, n43438, n43823, n43822, n43437, 
        n35823, n43821, n43820, n43819, n35819, n35803, n35728, 
        n43436, n29388, n29387, n43435, n43818, n43817, n43434, 
        n43816, n43815, n43814, n43813, n43433, n43812, n43811, 
        n15_adj_5483, n29386, n29385, n29384, n14_adj_5484, n15_adj_5485, 
        \FRAME_MATCHER.i_31__N_2843 , \FRAME_MATCHER.i_31__N_2845 , n43432, 
        n43810, n48264, n43809, n33, n32, n31, n30, n29, n28, 
        n27, n26, n25_adj_5486, n24_adj_5487, n23_adj_5488, n22_adj_5489, 
        n21_adj_5490, n20_adj_5491, n19_adj_5492, n18_adj_5493, n17_adj_5494, 
        n16_adj_5495, n15_adj_5496, n14_adj_5497, n13_adj_5498, n12_adj_5499, 
        n11_adj_5500, n10_adj_5501, n9_adj_5502, n8_adj_5503, n7_adj_5504, 
        n6_adj_5505, n5_adj_5506, n4_adj_5507, n3_adj_5508, n2_adj_5509, 
        n12_adj_5510, n49533, n9_adj_5511, n25_adj_5512, n24_adj_5513, 
        n23_adj_5514, n22_adj_5515, n21_adj_5516, n20_adj_5517, n19_adj_5518, 
        n18_adj_5519, n17_adj_5520, n16_adj_5521, n15_adj_5522, n14_adj_5523, 
        n13_adj_5524, n12_adj_5525, n11_adj_5526, n10_adj_5527, n9_adj_5528, 
        n8_adj_5529, n7_adj_5530, n6_adj_5531, n5_adj_5532, n4_adj_5533, 
        n3_adj_5534, n2_adj_5535, n36101, n10_adj_5536, n43808, n43431, 
        n43430, n43807, n2573, n49790, n43429, n29966, n29965, 
        n6272, n29959, n29958, n29957, n29956, n29955, n6_adj_5537, 
        n29954, n29953, n29952, n29378, n43806, n43805, n29951, 
        n29950, n29949, n29948, n29377, n29947, n29946, n5_adj_5538, 
        n43804, n29945, n29944, n29943, n29942, n29941, n29940, 
        n43803, n43802, n43428, n43801, n43800, n43427, n43426, 
        n43799, n43798, n43425, n43797, n43796, n43795, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(37[23:31])
    
    wire n4_adj_5539, n43794, n43793, n29939, n29938, n29376, n29937, 
        n29375, n29374, n29936, n29373, n43792, n29372, n43791, 
        n29371, n29370, n29369, n43790, n29935, n43789, n43788, 
        n29934;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3996 ;
    
    wire n55554, n29933, n40, n32_adj_5540, n24_adj_5541, n55879, 
        n43787, n43786, n26_adj_5542, n19_adj_5543, n29932;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev, n29931, n29930, n29929, n29928, n29927, position_31__N_4108, 
        n29926, n29925, n29924, n29923, n29922, n29921, n29920, 
        n29919, n29918, n29917, n29916, n29915, n24565, n29914, 
        n29913, n29912, n29911, n29910, n29909, n29908, n29907, 
        n29906, n29905, n29904, n29903, n29902, n29901, n29900, 
        n29899, n4910, n4909, n4908, n4907, n4906, n4904, n4903, 
        n4902, n4901, n4900, n4899, n4898, n4897, n4896, n4895, 
        n4894, n4893, n4892, n4891, n4890, n4889, n4888, n4887, 
        n4886, n4885, n4884, n4883, n29898, n29897, n43785, n29368, 
        n29896, n29895, n29366, n29894, n29893, n29892, n29891, 
        n29890, n29889;
    wire [1:0]a_new_adj_5703;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev_adj_5545, n29888, n29887, n29886, n29885, n29884, 
        position_31__N_4108_adj_5546, n29883, n29882, n29881, n29880, 
        n29879, n29878, n29877, n29876, n29875, n29874, n29186, 
        n29873, n29872, n29184, n29871, n29870, n29869, n51089, 
        n29868, n29867, n43784, n29859, n29365, n29364, n29858, 
        n29857, n29856, n29855, n29854, n29853, n29363, n43783, 
        rw;
    wire [7:0]state_adj_5716;   // verilog/eeprom.v(23[11:16])
    
    wire n43782, n43781, n55556, n43780, n29852, n29851, n28795, 
        n29850, n29849, n29848, n29847, n29846, n17_adj_5549, n16_adj_5550, 
        n15_adj_5551, n13_adj_5552, n11_adj_5553, n55756, n9_adj_5554, 
        n8_adj_5555, n7_adj_5556, n6_adj_5557, n5_adj_5558, n4_adj_5559, 
        n29845, clk_out;
    wire [15:0]data_adj_5722;   // verilog/tli4970.v(27[14:18])
    wire [7:0]state_adj_5724;   // verilog/tli4970.v(29[13:18])
    
    wire n43779, n29844, n29843, n29362, n29361, n29360, n29358, 
        n29357, n29842, n29841, n29840, n29839, n29838, n5_adj_5570, 
        n43778, n63, n43777, n6_adj_5571, n29837, n29836, n29835, 
        n43776, n29834, n29833, n29832, n29831, n29830, n29829, 
        n29828, n29827, n29826, n29825, n29824, n29823, n29822, 
        n29821, n29820, n29819, n43775, n43774, n29818, n29817, 
        n29816, n29815, n28762, n43773, n29814, n29813, n29812, 
        n28758, n29811, n29810, n29809, n29808, n29807, n29805, 
        n29804, state_7__N_4499, n29803, n29355, n29354, n29353, 
        n29802, n29801, n29800, n29799, n29798, n29797, n29796, 
        n29795, n29794, n29793, n29792, n29791, n29790, n29789, 
        n29788, n24_adj_5572, n55472, n19_adj_5573, n17_adj_5574, 
        n16_adj_5575, n15_adj_5576, n13_adj_5577, n11_adj_5578, n29787, 
        n19_adj_5579, n17_adj_5580, n16_adj_5581, n15_adj_5582, n13_adj_5583, 
        n11_adj_5584, n9_adj_5585, n29786, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n29785, n29784, n29783, n29782, n29781, n29780, n8_adj_5586, 
        n43210, n29779, n29778, n29777, n29776, n29775, n29774, 
        n29773, n29772, n43772, n43209, n43771, n43770, n43769, 
        n29771, n36808, n29770, n29769, n7_adj_5587, n6_adj_5588, 
        n29768, n5_adj_5589, n29767;
    wire [2:0]r_SM_Main_2__N_3777;
    
    wire n52856, n29766, n29352, n29763, n29762, n29761, n29760, 
        n29759, n29758, n29757, n29756, n29755, n29754, n29753, 
        n29752, n29751;
    wire [2:0]r_SM_Main_adj_5734;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5736;   // verilog/uart_tx.v(33[16:27])
    
    wire n43768, n43767, n43766;
    wire [2:0]r_SM_Main_2__N_3848;
    
    wire n29750, n26_adj_5594, n29749, n29748, n29351, n29747, n43765, 
        n29741, n4_adj_5595, n29740, n29736, n29735, n29732, n29727;
    wire [7:0]state_adj_5747;   // verilog/i2c_controller.v(33[12:17])
    
    wire n29726, n29725;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n29349, n29724, n29723, enable_slow_N_4393, n29722, n7_adj_5597, 
        n43764, n43763, n43762, n29721, n43208, n29720, n29719;
    wire [7:0]state_7__N_4290;
    
    wire n4_adj_5598, n29718, n29717, n29716, n7354, n29714, n29713, 
        n29347, n43761, n43760, n29712, n29711, n29710, n29346, 
        n29709;
    wire [7:0]state_7__N_4306;
    
    wire n29345, n29708, n43759, n55330, n29707, n29706, n29705, 
        n29704, n29703, n29702, n29701, n43758, n43757, n43207, 
        n29700, n29049, n9_adj_5599, n8_adj_5600, n7_adj_5601, n6_adj_5602, 
        n5_adj_5603, n4_adj_5604, n29699, n50454, n29698, n29697, 
        n29696, n29343, n29341, n29340, n29339, n29338, n29337, 
        n7974, n29695, n29694, n29693, n29692, n50462, n43756, 
        n29691, n29690, n29689, n29336, n29335, n29334, n29333, 
        n29332, n29331, n29330, n29329, n29328, n29327, n29326, 
        n29688, n29687, n29325, n29324, n50464, n29686, n29685, 
        n43755, n29684, n29683, n29682, n29323, n29681, n29680, 
        n29679, n29678, n29677, n29676, n29256, n29675, n29674, 
        n29673, n29672, n29671, n29670, n29669, n29668, n29667, 
        n29666, n29665, n29664, n28689, n29663, n29662, n29661, 
        n29660, n29659, n50497, n29658, n29657, n29656, n7593, 
        n29655, n29654, n29653, n29652, n29651, n29322, n29650, 
        n833, n832, n831, n830, n829, n828, n861, n50867, n896, 
        n897, n898, n899, n900, n901, n50765, n927, n928, n929, 
        n930, n931, n932, n933, n960, n29649, n50786, n56404, 
        n995, n996, n997, n998, n999, n1000, n1001, n51036, 
        n50620, n50602, n1026, n1027, n1028, n1029, n1030, n1031, 
        n1032, n1033, n1059, n28664, n1093, n1094, n1095, n1096, 
        n1097, n1098, n1099, n1100, n1101, n1125, n1126, n1127, 
        n1128, n1129, n1130, n1131, n1132, n1133, n1158, n43206, 
        n4_adj_5605, n43754, n1193, n1194, n1195, n1196, n1197, 
        n1198, n1199, n1200, n1201, n4_adj_5606, n1224, n1225, 
        n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, 
        n1257, n9_adj_5607, n1292, n1293, n1294, n1295, n1296, 
        n1297, n1298, n1299, n1300, n1301, n1323, n1324, n1325, 
        n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, 
        n1356, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
        n1397, n1398, n1399, n1400, n1401, n1422, n1423, n1424, 
        n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
        n1433, n1455, n1490, n1491, n1492, n1493, n1494, n1495, 
        n1496, n1497, n1498, n1499, n1500, n1501, n1521, n1522, 
        n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, 
        n1531, n1532_adj_5608, n1533_adj_5609, n1554_adj_5610, n43205, 
        n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
        n1597, n1598, n1599, n1600, n1601, n1620, n1621, n1622, 
        n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
        n1631, n1632, n1633, n56120, n1653, n43204, n43203, n43753, 
        n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
        n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1719, 
        n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, 
        n1728, n1729, n1730, n1731, n1732, n1733, n1752, n43113, 
        n29648, n1787, n1788, n1789, n1790, n1791, n1792, n1793, 
        n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
        n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
        n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
        n1851, n43752, n1886, n1887, n1888, n1889, n1890, n1891, 
        n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
        n1900, n1901, n1917, n1918, n1919, n1920, n1921, n1922, 
        n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, 
        n1931, n1932, n1933, n1950, n1985, n1986, n1987, n1988, 
        n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
        n1997, n1998, n1999, n2000, n2001, n2016, n2017, n2018, 
        n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
        n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2049, 
        n56392, n2084, n2085, n2086, n2087, n2088, n2089, n2090, 
        n2091_adj_5611, n2092, n2093, n2094, n2095, n2096, n2097, 
        n2098, n2099, n2100, n2101, n43751, n2115, n2116, n2117, 
        n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2126, 
        n2127, n2128, n2129, n2130, n2131, n2132, n2133, n43750, 
        n43749, n43748, n2148, n29647, n43202, n43747, n2183, 
        n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, 
        n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, 
        n2200, n2201, n2214, n2215, n2216, n2217, n2218, n2219, 
        n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, 
        n2228, n2229, n2230, n2231, n2232, n2233_adj_5612, n2247, 
        n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, 
        n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
        n2298, n2299, n2300, n2301, n2313, n2314, n2315, n2316, 
        n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, 
        n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
        n2333, n2346, n2381, n2382, n2383, n2384, n2385, n2386, 
        n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, 
        n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2412, 
        n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, 
        n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, 
        n2429, n2430, n2431, n2432, n2433, n2445, n48368, n2479, 
        n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, 
        n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, 
        n2496, n2497, n2498, n2499, n2500, n2501, n2511, n2512, 
        n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
        n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, 
        n2529, n2530, n2531, n2532, n2533, n2544, n29646, n2579, 
        n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, 
        n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, 
        n2596, n2597, n2598, n2599, n2600, n2601, n2610, n2611, 
        n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
        n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, 
        n2628, n2629, n2630, n2631, n2632, n2633, n24373, n55883, 
        n2643, n43746, n2678, n2679, n2680, n2681, n2682, n2683, 
        n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, 
        n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
        n2700, n2701, n2709, n2710, n2711, n2712, n2713, n2714, 
        n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
        n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, 
        n2731, n2732, n2733, n2742, n43201, n28640, n2777, n2778, 
        n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
        n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, 
        n2795, n2796, n2797, n2798, n2799, n2800, n2801, n29645, 
        n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
        n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
        n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, 
        n2832, n2833, n2841, n27227, n55374, n56270, n2876, n2877, 
        n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
        n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
        n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
        n27284, n47754, n2907, n2908, n2909, n2910, n2911, n2912, 
        n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
        n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
        n2929, n2930, n2931, n2932, n2933, n2940, n2975, n2976, 
        n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, 
        n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
        n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
        n3001, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
        n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, 
        n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
        n3029, n3030, n3031, n3032, n3033, n3039, n49729, n3073, 
        n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
        n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
        n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, 
        n3098, n3099, n3100, n3101, n3105, n3106, n3107, n3108, 
        n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
        n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, 
        n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
        n3133, n48646, n3138, n3173, n3174, n3175, n3176, n3177, 
        n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, 
        n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
        n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
        n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
        n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
        n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, 
        n3228, n3229, n3230, n3231, n3232, n3233, n3237, n3271, 
        n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
        n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, 
        n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, 
        n3296, n3298, n3299, n3300, n3301, n29644, n52032, n48638, 
        n56332, n56314, n56308, n56302, n29643, n24_adj_5613, n48616, 
        n62, n52004, n27140, n27143, n29146, n28583, n50546, n50549, 
        n51996, n27267, n29321, n44246, n44245, n51988, n28559, 
        n51982, n5_adj_5614, n51976, n51970, n56209, n55850, n55505, 
        n51964, n51962, n63_adj_5615, n51954, n51950, n51948, n29320, 
        n50597, n27294, n27287, n56195, n51940, n51938, n22902, 
        n54328, n51932, n51924, n48016, n27137, n55724, n56181, 
        n55470, n55819, n51918, n51912, n51908, n51906, n43200, 
        n51892, n56167, n51886, n43199, n44244, n43745, n43744, 
        n51880, n43198, n51874, n51872, n29319, n51864, n54311, 
        n56150, n51856, n50599, n51850, n51844, n5_adj_5616, n51838, 
        n29318, n29317, n29316, n29315, n29314, n29313, n29312, 
        n54298, n10_adj_5617, n51834, n44243, n44242, n44241, n44240, 
        n44239, n51832, n29311, n48, n49, n50, n51, n52, n53, 
        n54, n55, n29310, n44238, n44237, n44236, n56237, n44235, 
        n10832, n51818, n51812, n54294, n43197, n43743, n44234, 
        n44233, n43742, n49684, n51806, n43741, n44232, n43196, 
        n51802, n44231, n44230, n44229, n44228, n44227, n54290, 
        n43740, n43739, n43738, n43195, n44226, n48226, n36692, 
        n51794, n56116, n51780, n51774, n29308, n29307, n29306, 
        n29305, n29304, n29303, n29301, n29300, n29299, n29298, 
        n29297, n29296, n29295, n29294, n29293, n29292, n29291, 
        n29290, n29289, n29288, n29287, n29286, n29284, n29283, 
        n29282, n29280, n29279, n29278, n29277, n51768, n51766, 
        n43737, n43736, n43194, n44225, n43735, n43112, n51752, 
        n44224, n44223, n43734, n43193, n43733, n51748, n43732, 
        n43731, n43730, n43729, n51746, n50777, n44222, n43192, 
        n43191, n43190, n43728, n44221, n44220, n44219, n44218, 
        n44217, n43727, n43726, n43111, n51740, n56554, n49830, 
        n55331, n51730, n29276, n29275, n29274, n29273, n29269, 
        n56096, n51724, n29268, n29267, n29266, n29265, n29264, 
        n29263, n29261, n29260, n29483, n29482, n29481, n29480, 
        n29479, n29478, n29477, n29476, n51720, n43725, n43189, 
        n44216, n49802, n29468, n29467, n29466, n29465, n29464, 
        n29463, n29462, n29461, n29460, n29459, n29458, n29457, 
        n29456, n29455, n29454, n29453, n29452, n29451, n29450, 
        n29449, n29448, n29447, n29446, n29445, n29442, n29441, 
        n29440, n29439, n29438, n29437, n43188, n51708, n29259, 
        n29258, n29257, n29436, n29434, n29433, n29432, n29431, 
        n29430, n29429, n51706, n56075, n51696, n43187, n51684, 
        n2_adj_5618, n3_adj_5619, n4_adj_5620, n5_adj_5621, n6_adj_5622, 
        n7_adj_5623, n8_adj_5624, n9_adj_5625, n10_adj_5626, n11_adj_5627, 
        n12_adj_5628, n13_adj_5629, n14_adj_5630, n15_adj_5631, n16_adj_5632, 
        n17_adj_5633, n18_adj_5634, n19_adj_5635, n20_adj_5636, n21_adj_5637, 
        n22_adj_5638, n23_adj_5639, n24_adj_5640, n25_adj_5641, n26_adj_5642, 
        n27_adj_5643, n28_adj_5644, n29_adj_5645, n30_adj_5646, n31_adj_5647, 
        n32_adj_5648, n33_adj_5649, n51678, n51672, n43186, n43185, 
        n43724, n43723, n56524, n43722, n43721, n51662, n52838, 
        n51654, n56548, n51652, n56055, n51646, n51644, n43720, 
        n48565, n52805, n43184, n43719, n43718, n51630, n43183, 
        n43182, n43717, n43181, n43180, n6_adj_5650, n43716, n43093, 
        n51618, n43715, n43110, n43714, n43713, n51612, n43179, 
        n43109, n43108, n51606, n43712, n43092, n27232, n54253, 
        n43178, n51600, n43177, n43711, n54252, n51594, n43710, 
        n43107, n43709, n51592, n54251, n43708, n43707, n43706, 
        n43176, n43705, n51590, n43175, n56033, n43340, n43704, 
        n43174, n43173, n43703, n43091, n43090, n43702, n43339, 
        n51576, n43701, n51570, n43338, n43172, n43700, n43089, 
        n49816, n43699, n51564, n43171, n43106, n43105, n43698, 
        n43697, n43696, n43695, n43694, n43337, n51560, n43336, 
        n43693, n43692, n43691, n43690, n43335, n43689, n54250, 
        n43688, n43687, n43334, n43686, n43685, n50459, n43684, 
        n54249, n43683, n43682, n49761, n43681, n43680, n43679, 
        n43678, n43333, n43677, n27256, n43332, n43676, n43170, 
        n43675, n43674, n43673, n43672, n27262, n43671, n43169, 
        n54248, n43670, n43081, n43669, n43668, n43667, n51550, 
        n43666, n43665, n43331, n54247, n43330, n43664, n43663, 
        n43329, n43662, n43661, n43660, n43168, n43328, n43659, 
        n43658, n43167, n43657, n49772, n43656, n43655, n43654, 
        n43327, n43166, n51544, n43653, n19731, n43652, n43651, 
        n43650, n43649, n43648, n43326, n43647, n43646, n43325, 
        n51538, n43645, n43324, n43644, n43643, n43642, n43641, 
        n43640, n51532, n43323, n43322, n43639, n43638, n43637, 
        n51530, n43165, n43321, n43636, n43635, n43634, n43164, 
        n43320, n43319, n43633, n43632, n43318, n43163, n43631, 
        n43630, n43162, n43629, n43628, n43627, n43626, n43625, 
        n43624, n43623, n43622, n43621, n43620, n27118, n13_adj_5651, 
        n15_adj_5652, n21_adj_5653, n27_adj_5654, n43161, n29_adj_5655, 
        n43619, n33_adj_5656, n43618, n35, n43617, n43, n43616, 
        n48270, n51520, n52823, n56010, n51518, n51516, n49746, 
        n8_adj_5657, n51514, n51512, n51510, n51508, n51506, n51504, 
        n51502, n54237, n51498, n51496, n51494, n51490, n56542, 
        n51484, n51482, n14_adj_5658, n51478, n51476, n51474, n51472, 
        n55986, n10_adj_5659, n14_adj_5660, n10_adj_5661, n51466, 
        n51460, n51454, n51444, n51438, n51432, n49744, n51428, 
        n51422, n51420, n49704, n49699, n51406, n55788, n6_adj_5662, 
        n51402, n51394, n54231, n51220, n51386, n51380, n7_adj_5663, 
        n4_adj_5664, n8_adj_5665, n7_adj_5666, n51372, n51366, n51360, 
        n51354, n51348, n51212, n51342, n12_adj_5667, n56288, n48472, 
        n52728, n51338, n55557, n55555, n55960, n51334, n55533, 
        n55532, n56536, n6_adj_5668;
    
    VCC i2 (.Y(VCC_net));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_22 (.CI(n43817), 
            .I0(n2714), .I1(VCC_net), .CO(n43818));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_21_lut (.I0(GND_net), 
            .I1(n2715), .I2(VCC_net), .I3(n43816), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40167_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55960));
    defparam i40167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_1039_17_lut (.I0(GND_net), .I1(n4889), .I2(n4914), .I3(n43332), 
            .O(n426)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF dir_205 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_263));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_4_lut (.I0(GND_net), 
            .I1(n1432), .I2(GND_net), .I3(n43565), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1377_3_lut (.I0(n2022), 
            .I1(n2089), .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_281_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[22]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i23_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_123[22]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_18_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_5465));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40357_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56150));
    defparam i40357_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE dti_207 (.Q(dti), .C(clk16MHz), .E(n28559), .D(dti_N_527));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i902_3_lut (.I0(n1323), .I1(n1390), 
            .I2(n1356), .I3(GND_net), .O(n1422));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i902_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(control_mode[3]), .I1(control_mode[4]), .I2(control_mode[2]), 
            .I3(control_mode[6]), .O(n52032));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[0]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 i1_3_lut (.I0(n52032), .I1(control_mode[7]), .I2(control_mode[5]), 
            .I3(GND_net), .O(n27284));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_21 (.CI(n43816), 
            .I0(n2715), .I1(VCC_net), .CO(n43817));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_20_lut (.I0(GND_net), 
            .I1(n2716), .I2(VCC_net), .I3(n43815), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_4 (.CI(n43565), 
            .I0(n1432), .I1(GND_net), .CO(n43566));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_20 (.CI(n43815), 
            .I0(n2716), .I1(VCC_net), .CO(n43816));
    SB_CARRY add_1039_17 (.CI(n43332), .I0(n4889), .I1(n4914), .CO(n43333));
    SB_CARRY add_175_31 (.CI(n43184), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n43185));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_3_lut (.I0(GND_net), 
            .I1(n1433), .I2(VCC_net), .I3(n43564), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_19_lut (.I0(GND_net), 
            .I1(n2717), .I2(VCC_net), .I3(n43814), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_3 (.CI(n43564), 
            .I0(n1433), .I1(VCC_net), .CO(n43565));
    SB_LUT4 add_1039_16_lut (.I0(GND_net), .I1(n4890), .I2(n4915), .I3(n43331), 
            .O(n427)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_1039_16 (.CI(n43331), .I0(n4890), .I1(n4915), .CO(n43332));
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[0]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4306[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_99[0]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_2_lut (.I0(GND_net), 
            .I1(n525), .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_2 (.CI(VCC_net), 
            .I0(n525), .I1(GND_net), .CO(n43564));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_13_lut (.I0(GND_net), 
            .I1(n1323), .I2(VCC_net), .I3(n43563), .O(n1390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_15_lut (.I0(GND_net), .I1(n4891), .I2(n4916), .I3(n43330), 
            .O(n428)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_15_lut.LUT_INIT = 16'hC33C;
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_1039_15 (.CI(n43330), .I0(n4891), .I1(n4916), .CO(n43331));
    SB_LUT4 add_175_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n43183), .O(n1535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_30_lut.LUT_INIT = 16'hC33C;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .GND_net(GND_net), .neopxl_color({neopxl_color}), .\state[1] (state[1]), 
            .\state[0] (state[0]), .n28689(n28689), .\state_3__N_639[1] (state_3__N_639[1]), 
            .timer({timer}), .n49594(n49594), .VCC_net(VCC_net), .LED_c(LED_c), 
            .n29258(n29258), .n29700(n29700), .n29699(n29699), .n29698(n29698), 
            .n29697(n29697), .n29696(n29696), .n29695(n29695), .n29694(n29694), 
            .n29693(n29693), .n29692(n29692), .n29691(n29691), .n29690(n29690), 
            .n29689(n29689), .n29688(n29688), .n29684(n29684), .n29683(n29683), 
            .n29682(n29682), .n29681(n29681), .n29680(n29680), .n29679(n29679), 
            .n29678(n29678), .n29677(n29677), .n29676(n29676), .n29675(n29675), 
            .n29674(n29674), .n29673(n29673), .n29672(n29672), .n29671(n29671), 
            .n29670(n29670), .n29669(n29669), .n29668(n29668), .n29667(n29667), 
            .NEOPXL_c(NEOPXL_c), .n29436(n29436)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(50[24] 56[2])
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_19 (.CI(n43814), 
            .I0(n2717), .I1(VCC_net), .CO(n43815));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_18_lut (.I0(GND_net), 
            .I1(n2718), .I2(VCC_net), .I3(n43813), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_30 (.CI(n43183), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n43184));
    SB_LUT4 add_175_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n43182), .O(n1536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_12_lut (.I0(GND_net), 
            .I1(n1324), .I2(VCC_net), .I3(n43562), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1730 (.I0(control_mode[0]), .I1(n27284), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(284[5:22])
    defparam i1_3_lut_adj_1730.LUT_INIT = 16'hfdfd;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_12 (.CI(n43562), 
            .I0(n1324), .I1(VCC_net), .CO(n43563));
    SB_LUT4 mux_281_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[23]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_18 (.CI(n43813), 
            .I0(n2718), .I1(VCC_net), .CO(n43814));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_11_lut (.I0(GND_net), 
            .I1(n1325), .I2(VCC_net), .I3(n43561), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_17_lut (.I0(GND_net), 
            .I1(n2719), .I2(VCC_net), .I3(n43812), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_17 (.CI(n43812), 
            .I0(n2719), .I1(VCC_net), .CO(n43813));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_16_lut (.I0(GND_net), 
            .I1(n2720), .I2(VCC_net), .I3(n43811), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_16 (.CI(n43811), 
            .I0(n2720), .I1(VCC_net), .CO(n43812));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_15_lut (.I0(GND_net), 
            .I1(n2721), .I2(VCC_net), .I3(n43810), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_15 (.CI(n43810), 
            .I0(n2721), .I1(VCC_net), .CO(n43811));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_11 (.CI(n43561), 
            .I0(n1325), .I1(VCC_net), .CO(n43562));
    SB_LUT4 mux_276_i24_3_lut (.I0(encoder0_position_scaled[23]), .I1(motor_state_23__N_123[23]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i24_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_14_lut (.I0(GND_net), 
            .I1(n2722), .I2(VCC_net), .I3(n43809), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_14 (.CI(n43809), 
            .I0(n2722), .I1(VCC_net), .CO(n43810));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_13_lut (.I0(GND_net), 
            .I1(n2723), .I2(VCC_net), .I3(n43808), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_13 (.CI(n43808), 
            .I0(n2723), .I1(VCC_net), .CO(n43809));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_12_lut (.I0(GND_net), 
            .I1(n2724), .I2(VCC_net), .I3(n43807), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_14_lut (.I0(GND_net), .I1(n4892), .I2(n4917), .I3(n43329), 
            .O(n429)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_12 (.CI(n43807), 
            .I0(n2724), .I1(VCC_net), .CO(n43808));
    SB_CARRY add_1039_14 (.CI(n43329), .I0(n4892), .I1(n4917), .CO(n43330));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_11_lut (.I0(GND_net), 
            .I1(n2725), .I2(VCC_net), .I3(n43806), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_29 (.CI(n43182), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n43183));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_11 (.CI(n43806), 
            .I0(n2725), .I1(VCC_net), .CO(n43807));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_10_lut (.I0(GND_net), 
            .I1(n2726), .I2(VCC_net), .I3(n43805), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_10 (.CI(n43805), 
            .I0(n2726), .I1(VCC_net), .CO(n43806));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_9_lut (.I0(GND_net), 
            .I1(n2727), .I2(VCC_net), .I3(n43804), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_9 (.CI(n43804), 
            .I0(n2727), .I1(VCC_net), .CO(n43805));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_8_lut (.I0(GND_net), 
            .I1(n2728), .I2(VCC_net), .I3(n43803), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_8 (.CI(n43803), 
            .I0(n2728), .I1(VCC_net), .CO(n43804));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_7_lut (.I0(GND_net), 
            .I1(n2729), .I2(GND_net), .I3(n43802), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_13_lut (.I0(GND_net), .I1(n4893), .I2(n4918), .I3(n43328), 
            .O(n430)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_7 (.CI(n43802), 
            .I0(n2729), .I1(GND_net), .CO(n43803));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_6_lut (.I0(GND_net), 
            .I1(n2730), .I2(GND_net), .I3(n43801), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_6 (.CI(n43801), 
            .I0(n2730), .I1(GND_net), .CO(n43802));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_10_lut (.I0(GND_net), 
            .I1(n1326), .I2(VCC_net), .I3(n43560), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_10 (.CI(n43560), 
            .I0(n1326), .I1(VCC_net), .CO(n43561));
    SB_CARRY add_1039_13 (.CI(n43328), .I0(n4893), .I1(n4918), .CO(n43329));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_9_lut (.I0(GND_net), 
            .I1(n1327), .I2(VCC_net), .I3(n43559), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_5_lut (.I0(GND_net), 
            .I1(n2731), .I2(VCC_net), .I3(n43800), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_12_lut (.I0(GND_net), .I1(n4894), .I2(n4919), .I3(n43327), 
            .O(n431)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_9 (.CI(n43559), 
            .I0(n1327), .I1(VCC_net), .CO(n43560));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_5 (.CI(n43800), 
            .I0(n2731), .I1(VCC_net), .CO(n43801));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_4_lut (.I0(GND_net), 
            .I1(n2732), .I2(GND_net), .I3(n43799), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_12 (.CI(n43327), .I0(n4894), .I1(n4919), .CO(n43328));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_4 (.CI(n43799), 
            .I0(n2732), .I1(GND_net), .CO(n43800));
    SB_LUT4 add_1039_11_lut (.I0(GND_net), .I1(n4895), .I2(n4920), .I3(n43326), 
            .O(n432)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_8_lut (.I0(GND_net), 
            .I1(n1328), .I2(VCC_net), .I3(n43558), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_11 (.CI(n43326), .I0(n4895), .I1(n4920), .CO(n43327));
    SB_LUT4 add_1039_10_lut (.I0(GND_net), .I1(n4896), .I2(n4921), .I3(n43325), 
            .O(n433)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_3_lut (.I0(GND_net), 
            .I1(n2733), .I2(VCC_net), .I3(n43798), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_8 (.CI(n43558), 
            .I0(n1328), .I1(VCC_net), .CO(n43559));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_7_lut (.I0(GND_net), 
            .I1(n1329), .I2(GND_net), .I3(n43557), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_7 (.CI(n43557), 
            .I0(n1329), .I1(GND_net), .CO(n43558));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_6_lut (.I0(GND_net), 
            .I1(n1330), .I2(GND_net), .I3(n43556), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_6 (.CI(n43556), 
            .I0(n1330), .I1(GND_net), .CO(n43557));
    SB_CARRY add_1039_10 (.CI(n43325), .I0(n4896), .I1(n4921), .CO(n43326));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_3 (.CI(n43798), 
            .I0(n2733), .I1(VCC_net), .CO(n43799));
    SB_LUT4 add_1039_9_lut (.I0(GND_net), .I1(n4897), .I2(n4922), .I3(n43324), 
            .O(n434)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_2_lut (.I0(GND_net), 
            .I1(n538), .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_9 (.CI(n43324), .I0(n4897), .I1(n4922), .CO(n43325));
    SB_LUT4 add_1039_8_lut (.I0(GND_net), .I1(n4898), .I2(n4923), .I3(n43323), 
            .O(n435)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_2 (.CI(VCC_net), 
            .I0(n538), .I1(GND_net), .CO(n43798));
    SB_CARRY add_1039_8 (.CI(n43323), .I0(n4898), .I1(n4923), .CO(n43324));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_5_lut (.I0(GND_net), 
            .I1(n1331), .I2(VCC_net), .I3(n43555), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_7_lut (.I0(GND_net), .I1(n4899), .I2(n4924), .I3(n43322), 
            .O(n436)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n43181), .O(n1537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_26_lut (.I0(n55879), 
            .I1(n2610), .I2(VCC_net), .I3(n43797), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_25_lut (.I0(GND_net), 
            .I1(n2611), .I2(VCC_net), .I3(n43796), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_25 (.CI(n43796), 
            .I0(n2611), .I1(VCC_net), .CO(n43797));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_5 (.CI(n43555), 
            .I0(n1331), .I1(VCC_net), .CO(n43556));
    SB_CARRY add_1039_7 (.CI(n43322), .I0(n4899), .I1(n4924), .CO(n43323));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_24_lut (.I0(GND_net), 
            .I1(n2612), .I2(VCC_net), .I3(n43795), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_6_lut (.I0(GND_net), .I1(n4900), .I2(n4925), .I3(n43321), 
            .O(n437)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_4_lut (.I0(GND_net), 
            .I1(n1332), .I2(GND_net), .I3(n43554), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_28 (.CI(n43181), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n43182));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_24 (.CI(n43795), 
            .I0(n2612), .I1(VCC_net), .CO(n43796));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_23_lut (.I0(GND_net), 
            .I1(n2613), .I2(VCC_net), .I3(n43794), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_23 (.CI(n43794), 
            .I0(n2613), .I1(VCC_net), .CO(n43795));
    SB_CARRY add_1039_6 (.CI(n43321), .I0(n4900), .I1(n4925), .CO(n43322));
    SB_LUT4 add_1039_5_lut (.I0(GND_net), .I1(n4901), .I2(n4926), .I3(n43320), 
            .O(n438)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_4 (.CI(n43554), 
            .I0(n1332), .I1(GND_net), .CO(n43555));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_3_lut (.I0(GND_net), 
            .I1(n1333), .I2(VCC_net), .I3(n43553), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_22_lut (.I0(GND_net), 
            .I1(n2614), .I2(VCC_net), .I3(n43793), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_22 (.CI(n43793), 
            .I0(n2614), .I1(VCC_net), .CO(n43794));
    SB_LUT4 add_175_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n43180), .O(n1538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_5 (.CI(n43320), .I0(n4901), .I1(n4926), .CO(n43321));
    SB_LUT4 add_1039_4_lut (.I0(GND_net), .I1(n4902), .I2(n4927), .I3(n43319), 
            .O(n439)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_21_lut (.I0(GND_net), 
            .I1(n2615), .I2(VCC_net), .I3(n43792), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_21 (.CI(n43792), 
            .I0(n2615), .I1(VCC_net), .CO(n43793));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_20_lut (.I0(GND_net), 
            .I1(n2616), .I2(VCC_net), .I3(n43791), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_20 (.CI(n43791), 
            .I0(n2616), .I1(VCC_net), .CO(n43792));
    SB_CARRY add_175_27 (.CI(n43180), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n43181));
    SB_CARRY add_1039_4 (.CI(n43319), .I0(n4902), .I1(n4927), .CO(n43320));
    SB_LUT4 add_175_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n43179), .O(n1539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_3 (.CI(n43553), 
            .I0(n1333), .I1(VCC_net), .CO(n43554));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_19_lut (.I0(GND_net), 
            .I1(n2617), .I2(VCC_net), .I3(n43790), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_16 (.CI(n43117), .I0(duty[17]), .I1(n56288), .CO(n43118));
    SB_CARRY add_175_26 (.CI(n43179), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n43180));
    SB_LUT4 add_1039_3_lut (.I0(GND_net), .I1(n4903), .I2(n4928), .I3(n43318), 
            .O(n440)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_900_2_lut (.I0(GND_net), 
            .I1(n524), .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n43178), .O(n1540)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_19 (.CI(n43790), 
            .I0(n2617), .I1(VCC_net), .CO(n43791));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_900_2 (.CI(VCC_net), 
            .I0(n524), .I1(GND_net), .CO(n43553));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_18_lut (.I0(GND_net), 
            .I1(n2618), .I2(VCC_net), .I3(n43789), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_15_lut (.I0(current[15]), .I1(duty[16]), .I2(n56288), 
            .I3(n43116), .O(n257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_15_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 unary_minus_18_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15299_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n50602), 
            .I3(GND_net), .O(n29375));   // verilog/coms.v(128[12] 303[6])
    defparam i15299_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15300_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n50602), 
            .I3(GND_net), .O(n29376));   // verilog/coms.v(128[12] 303[6])
    defparam i15300_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i11_3_lut (.I0(encoder0_position_scaled_23__N_327[10]), 
            .I1(n23_adj_5488), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1593_3_lut (.I0(n534), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1660_3_lut (.I0(n2433), 
            .I1(n2500), .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i12_3_lut (.I0(encoder0_position_scaled_23__N_327[11]), 
            .I1(n22_adj_5489), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n533));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1525_rep_44_3_lut (.I0(n533), 
            .I1(n2301), .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1525_rep_44_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n7593), 
            .D(n1562), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n7593), 
            .D(n1561), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n7593), 
            .D(n1560), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1592_3_lut (.I0(n2333), 
            .I1(n2400), .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n7593), 
            .D(n1559), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1659_3_lut (.I0(n2432), 
            .I1(n2499), .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n7593), 
            .D(n1558), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n7593), 
            .D(n1557), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n7593), 
            .D(n1556), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n7593), 
            .D(n1555), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n7593), 
            .D(n1554), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n7593), .D(n1553), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n7593), .D(n1552), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n7593), .D(n1551), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n7593), .D(n1550), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n7593), .D(n1549), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n7593), .D(n1548), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(clk16MHz), 
            .E(n7593), .D(n1547), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(clk16MHz), 
            .E(n7593), .D(n1546), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i15301_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n50602), 
            .I3(GND_net), .O(n29377));   // verilog/coms.v(128[12] 303[6])
    defparam i15301_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15302_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n50602), 
            .I3(GND_net), .O(n29378));   // verilog/coms.v(128[12] 303[6])
    defparam i15302_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_18 (.CI(n43789), 
            .I0(n2618), .I1(VCC_net), .CO(n43790));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_17_lut (.I0(GND_net), 
            .I1(n2619), .I2(VCC_net), .I3(n43788), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_17 (.CI(n43788), 
            .I0(n2619), .I1(VCC_net), .CO(n43789));
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(clk16MHz), 
            .E(n7593), .D(n1545), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(clk16MHz), 
            .E(n7593), .D(n1544), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(clk16MHz), 
            .E(n7593), .D(n1543), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(clk16MHz), 
            .E(n7593), .D(n1542), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(clk16MHz), 
            .E(n7593), .D(n1541), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(clk16MHz), 
            .E(n7593), .D(n1540), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_16_lut (.I0(GND_net), 
            .I1(n2620), .I2(VCC_net), .I3(n43787), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n51212));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(clk16MHz), 
            .E(n7593), .D(n1539), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(clk16MHz), 
            .E(n7593), .D(n1538), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(clk16MHz), 
            .E(n7593), .D(n1537), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(clk16MHz), 
            .E(n7593), .D(n1536), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(clk16MHz), 
            .E(n7593), .D(n1535), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(clk16MHz), 
            .E(n7593), .D(n1534), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(clk16MHz), 
            .E(n7593), .D(n1533), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(clk16MHz), 
            .E(n7593), .D(n1532), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 i1_4_lut_adj_1731 (.I0(n7974), .I1(n20976), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n49436));
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'heaee;
    SB_LUT4 i2_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(n35728), .I2(\ID_READOUT_FSM.state [1]), 
            .I3(n49436), .O(n28795));
    defparam i2_4_lut.LUT_INIT = 16'h4c00;
    SB_LUT4 i12_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n7974), .I2(n28795), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n47754));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15308_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n50602), 
            .I3(GND_net), .O(n29384));   // verilog/coms.v(128[12] 303[6])
    defparam i15308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15309_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n50602), 
            .I3(GND_net), .O(n29385));   // verilog/coms.v(128[12] 303[6])
    defparam i15309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15310_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n50602), 
            .I3(GND_net), .O(n29386));   // verilog/coms.v(128[12] 303[6])
    defparam i15310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15311_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n50602), 
            .I3(GND_net), .O(n29387));   // verilog/coms.v(128[12] 303[6])
    defparam i15311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15312_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n50602), 
            .I3(GND_net), .O(n29388));   // verilog/coms.v(128[12] 303[6])
    defparam i15312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15313_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n50602), 
            .I3(GND_net), .O(n29389));   // verilog/coms.v(128[12] 303[6])
    defparam i15313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39931_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55724));
    defparam i39931_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15314_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n50602), 
            .I3(GND_net), .O(n29390));   // verilog/coms.v(128[12] 303[6])
    defparam i15314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15315_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n50602), 
            .I3(GND_net), .O(n29391));   // verilog/coms.v(128[12] 303[6])
    defparam i15315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15758_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29834));   // verilog/coms.v(128[12] 303[6])
    defparam i15758_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15759_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29835));   // verilog/coms.v(128[12] 303[6])
    defparam i15759_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15739_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29815));   // verilog/coms.v(128[12] 303[6])
    defparam i15739_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5512));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut (.I0(duty[0]), .I1(duty[23]), .I2(duty[1]), .I3(duty[2]), 
            .O(n211));   // verilog/TinyFPGA_B.v(111[25:31])
    defparam i14_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i15318_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n50602), 
            .I3(GND_net), .O(n29394));   // verilog/coms.v(128[12] 303[6])
    defparam i15318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15740_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29816));   // verilog/coms.v(128[12] 303[6])
    defparam i15740_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15741_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29817));   // verilog/coms.v(128[12] 303[6])
    defparam i15741_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15319_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n50602), 
            .I3(GND_net), .O(n29395));   // verilog/coms.v(128[12] 303[6])
    defparam i15319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15742_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29818));   // verilog/coms.v(128[12] 303[6])
    defparam i15742_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5513));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15743_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29819));   // verilog/coms.v(128[12] 303[6])
    defparam i15743_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1444_3_lut (.I0(n2121), 
            .I1(n2188), .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15185_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n35837), 
            .I3(n27227), .O(n29261));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15185_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15180_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position_scaled[11]), 
            .I2(n24373), .I3(GND_net), .O(n29256));   // verilog/coms.v(128[12] 303[6])
    defparam i15180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40303_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56096));
    defparam i40303_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1103_3_lut (.I0(n1620), 
            .I1(n1687), .I2(n1653), .I3(GND_net), .O(n1719));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15760_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29836));   // verilog/coms.v(128[12] 303[6])
    defparam i15760_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15320_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n50602), 
            .I3(GND_net), .O(n29396));   // verilog/coms.v(128[12] 303[6])
    defparam i15320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33803_4_lut (.I0(n26_adj_5594), .I1(state_adj_5716[0]), .I2(n6_adj_5650), 
            .I3(state_adj_5747[0]), .O(n49533));
    defparam i33803_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_3_lut_adj_1732 (.I0(state_adj_5716[1]), .I1(read), .I2(n49611), 
            .I3(GND_net), .O(n12_adj_5510));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_3_lut_adj_1732.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_4_lut_adj_1733 (.I0(n36101), .I1(n12_adj_5510), .I2(state_adj_5716[0]), 
            .I3(n49611), .O(n48226));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1733.LUT_INIT = 16'h88a8;
    SB_CARRY add_1039_3 (.CI(n43318), .I0(n4903), .I1(n4928), .CO(n43319));
    SB_LUT4 i15761_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29837));   // verilog/coms.v(128[12] 303[6])
    defparam i15761_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1039_2_lut (.I0(GND_net), .I1(n4904), .I2(n4929), .I3(GND_net), 
            .O(n441)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15762_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29838));   // verilog/coms.v(128[12] 303[6])
    defparam i15762_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15324_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n50602), 
            .I3(GND_net), .O(n29400));   // verilog/coms.v(128[12] 303[6])
    defparam i15324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5514));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15325_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n50602), 
            .I3(GND_net), .O(n29401));   // verilog/coms.v(128[12] 303[6])
    defparam i15325_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15763_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29839));   // verilog/coms.v(128[12] 303[6])
    defparam i15763_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15326_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n50602), 
            .I3(GND_net), .O(n29402));   // verilog/coms.v(128[12] 303[6])
    defparam i15326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15327_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n50602), 
            .I3(GND_net), .O(n29403));   // verilog/coms.v(128[12] 303[6])
    defparam i15327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15328_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n50602), 
            .I3(GND_net), .O(n29404));   // verilog/coms.v(128[12] 303[6])
    defparam i15328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15329_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n50602), 
            .I3(GND_net), .O(n29405));   // verilog/coms.v(128[12] 303[6])
    defparam i15329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15330_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n50602), 
            .I3(GND_net), .O(n29406));   // verilog/coms.v(128[12] 303[6])
    defparam i15330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15187_4_lut (.I0(state_7__N_4306[3]), .I1(data[1]), .I2(n10_adj_5617), 
            .I3(n27267), .O(n29263));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15187_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15188_4_lut (.I0(state_7__N_4306[3]), .I1(data[2]), .I2(n4), 
            .I3(n27262), .O(n29264));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15188_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15189_4_lut (.I0(state_7__N_4306[3]), .I1(data[3]), .I2(n4), 
            .I3(n27267), .O(n29265));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15189_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15331_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n50602), 
            .I3(GND_net), .O(n29407));   // verilog/coms.v(128[12] 303[6])
    defparam i15331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15190_4_lut (.I0(state_7__N_4306[3]), .I1(data[4]), .I2(n4_adj_5459), 
            .I3(n27262), .O(n29266));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15190_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15332_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n50602), 
            .I3(GND_net), .O(n29408));   // verilog/coms.v(128[12] 303[6])
    defparam i15332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15191_4_lut (.I0(state_7__N_4306[3]), .I1(data[5]), .I2(n4_adj_5459), 
            .I3(n27267), .O(n29267));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15191_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15192_4_lut (.I0(state_7__N_4306[3]), .I1(data[6]), .I2(n35819), 
            .I3(n27262), .O(n29268));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15192_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15193_4_lut (.I0(state_7__N_4306[3]), .I1(data[7]), .I2(n35819), 
            .I3(n27267), .O(n29269));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15193_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15333_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n50602), 
            .I3(GND_net), .O(n29409));   // verilog/coms.v(128[12] 303[6])
    defparam i15333_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15197_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position_scaled[9]), 
            .I2(n24373), .I3(GND_net), .O(n29273));   // verilog/coms.v(128[12] 303[6])
    defparam i15197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15198_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position_scaled[8]), 
            .I2(n24373), .I3(GND_net), .O(n29274));   // verilog/coms.v(128[12] 303[6])
    defparam i15198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15199_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position_scaled[23]), 
            .I2(n24373), .I3(GND_net), .O(n29275));   // verilog/coms.v(128[12] 303[6])
    defparam i15199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15200_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29276));   // verilog/coms.v(128[12] 303[6])
    defparam i15200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15201_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n50602), 
            .I3(GND_net), .O(n29277));   // verilog/coms.v(128[12] 303[6])
    defparam i15201_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15202_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n50602), 
            .I3(GND_net), .O(n29278));   // verilog/coms.v(128[12] 303[6])
    defparam i15202_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15203_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29279));   // verilog/coms.v(128[12] 303[6])
    defparam i15203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15334_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n50602), 
            .I3(GND_net), .O(n29410));   // verilog/coms.v(128[12] 303[6])
    defparam i15334_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15204_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n50620), .I3(GND_net), .O(n29280));   // verilog/coms.v(128[12] 303[6])
    defparam i15204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40402_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56195));
    defparam i40402_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15206_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29282));   // verilog/coms.v(128[12] 303[6])
    defparam i15206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15207_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29283));   // verilog/coms.v(128[12] 303[6])
    defparam i15207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15208_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29284));   // verilog/coms.v(128[12] 303[6])
    defparam i15208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1179_3_lut (.I0(n1728), 
            .I1(n1795), .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15335_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n50602), 
            .I3(GND_net), .O(n29411));   // verilog/coms.v(128[12] 303[6])
    defparam i15335_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n51220));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i15181_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n51220), .I3(GND_net), 
            .O(n29257));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40282_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56075));
    defparam i40282_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40090_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55883));
    defparam i40090_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1639_3_lut (.I0(n2412), 
            .I1(n2479), .I2(n2445), .I3(GND_net), .O(n2511));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1639_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n544));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40444_1_lut (.I0(n36808), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56237));
    defparam i40444_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2196_3_lut (.I0(n3225), 
            .I1(n3292), .I2(n3237), .I3(GND_net), .O(n21_adj_5653));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2192_3_lut (.I0(n3221), 
            .I1(n3288), .I2(n3237), .I3(GND_net), .O(n29_adj_5655));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2189_3_lut (.I0(n3218), 
            .I1(n3285), .I2(n3237), .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2190_3_lut (.I0(n3219), 
            .I1(n3286), .I2(n3237), .I3(GND_net), .O(n33_adj_5656));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2193_3_lut (.I0(n3222), 
            .I1(n3289), .I2(n3237), .I3(GND_net), .O(n27_adj_5654));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2200_3_lut (.I0(n3229), 
            .I1(n3296), .I2(n3237), .I3(GND_net), .O(n13_adj_5651));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5464));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1734 (.I0(n3220), .I1(n21_adj_5653), .I2(n3287), 
            .I3(n3237), .O(n51472));
    defparam i1_4_lut_adj_1734.LUT_INIT = 16'heefc;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(260[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1735 (.I0(n3227), .I1(n29_adj_5655), .I2(n3294), 
            .I3(n3237), .O(n51482));
    defparam i1_4_lut_adj_1735.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2199_3_lut (.I0(n3228), 
            .I1(n3295), .I2(n3237), .I3(GND_net), .O(n15_adj_5652));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(n3223), .I1(n33_adj_5656), .I2(n3290), 
            .I3(n3237), .O(n51478));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n3224), .I1(n35), .I2(n3291), .I3(n3237), 
            .O(n51476));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1738 (.I0(n51478), .I1(n3217), .I2(n3284), .I3(n3237), 
            .O(n51484));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'heefa;
    SB_LUT4 i1_4_lut_adj_1739 (.I0(n15_adj_5652), .I1(n51482), .I2(n51472), 
            .I3(n13_adj_5651), .O(n51490));
    defparam i1_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1740 (.I0(n3226), .I1(n27_adj_5654), .I2(n3293), 
            .I3(n3237), .O(n51474));
    defparam i1_4_lut_adj_1740.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1741 (.I0(n51474), .I1(n51490), .I2(n51484), 
            .I3(n51476), .O(n51494));
    defparam i1_4_lut_adj_1741.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1742 (.I0(n51494), .I1(n3216), .I2(n3283), .I3(n3237), 
            .O(n51496));
    defparam i1_4_lut_adj_1742.LUT_INIT = 16'heefa;
    SB_LUT4 i22446_4_lut (.I0(n544), .I1(n543), .I2(n3301), .I3(n3237), 
            .O(n36510));
    defparam i22446_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i22556_4_lut (.I0(n36510), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n36626));
    defparam i22556_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5649));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n54294), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5614));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.i_31__N_2843 ), .I1(n3303), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5607));   // verilog/coms.v(128[12] 303[6])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1743 (.I0(n3215), .I1(n51496), .I2(n3282), .I3(n3237), 
            .O(n51498));
    defparam i1_4_lut_adj_1743.LUT_INIT = 16'heefc;
    SB_LUT4 i22622_4_lut (.I0(n36626), .I1(n3232), .I2(n3299), .I3(n3237), 
            .O(n36692));
    defparam i22622_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2185_3_lut (.I0(n3214), 
            .I1(n3281), .I2(n3237), .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(n43), .I1(n36692), .I2(n51498), .I3(n5_adj_5614), 
            .O(n51502));
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1745 (.I0(n3213), .I1(n51502), .I2(n3280), .I3(n3237), 
            .O(n51504));
    defparam i1_4_lut_adj_1745.LUT_INIT = 16'heefc;
    SB_LUT4 i3_4_lut_adj_1746 (.I0(n48616), .I1(n4_adj_5606), .I2(n48672), 
            .I3(n9_adj_5607), .O(n51036));   // verilog/coms.v(128[12] 303[6])
    defparam i3_4_lut_adj_1746.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1747 (.I0(n3212), .I1(n51504), .I2(n3279), .I3(n3237), 
            .O(n51506));
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1748 (.I0(n63), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n51036), .I3(n22902), .O(n48016));   // verilog/coms.v(128[12] 303[6])
    defparam i1_4_lut_adj_1748.LUT_INIT = 16'hd5f5;
    SB_LUT4 i15210_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position_scaled[22]), 
            .I2(n24373), .I3(GND_net), .O(n29286));   // verilog/coms.v(128[12] 303[6])
    defparam i15210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1749 (.I0(n3211), .I1(n51506), .I2(n3278), .I3(n3237), 
            .O(n51508));
    defparam i1_4_lut_adj_1749.LUT_INIT = 16'heefc;
    SB_LUT4 i15211_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position_scaled[21]), 
            .I2(n24373), .I3(GND_net), .O(n29287));   // verilog/coms.v(128[12] 303[6])
    defparam i15211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15212_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position_scaled[20]), 
            .I2(n24373), .I3(GND_net), .O(n29288));   // verilog/coms.v(128[12] 303[6])
    defparam i15212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1750 (.I0(n3210), .I1(n51508), .I2(n3277), .I3(n3237), 
            .O(n51510));
    defparam i1_4_lut_adj_1750.LUT_INIT = 16'heefc;
    SB_LUT4 i15213_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(control_update), .I3(GND_net), .O(n29289));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1751 (.I0(n3209), .I1(n51510), .I2(n3276), .I3(n3237), 
            .O(n51512));
    defparam i1_4_lut_adj_1751.LUT_INIT = 16'heefc;
    SB_LUT4 i15214_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position_scaled[19]), 
            .I2(n24373), .I3(GND_net), .O(n29290));   // verilog/coms.v(128[12] 303[6])
    defparam i15214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1752 (.I0(n3208), .I1(n51512), .I2(n3275), .I3(n3237), 
            .O(n51514));
    defparam i1_4_lut_adj_1752.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(n3207), .I1(n51514), .I2(n3274), .I3(n3237), 
            .O(n51516));
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n3206), .I1(n51516), .I2(n3273), .I3(n3237), 
            .O(n51518));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'heefc;
    SB_LUT4 i15215_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position_scaled[18]), 
            .I2(n24373), .I3(GND_net), .O(n29291));   // verilog/coms.v(128[12] 303[6])
    defparam i15215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5515));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(n3205), .I1(n51518), .I2(n3272), .I3(n3237), 
            .O(n51520));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'heefc;
    SB_LUT4 i40447_4_lut (.I0(n51520), .I1(n3204), .I2(n3271), .I3(n3237), 
            .O(n36808));
    defparam i40447_4_lut.LUT_INIT = 16'h1105;
    SB_LUT4 i15216_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position_scaled[17]), 
            .I2(n24373), .I3(GND_net), .O(n29292));   // verilog/coms.v(128[12] 303[6])
    defparam i15216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2110_3_lut (.I0(n3107), 
            .I1(n3174), .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2116_3_lut (.I0(n3113), 
            .I1(n3180), .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2109_3_lut (.I0(n3106), 
            .I1(n3173), .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15764_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29840));   // verilog/coms.v(128[12] 303[6])
    defparam i15764_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40026_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55819));
    defparam i40026_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2123_3_lut (.I0(n3120), 
            .I1(n3187), .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15765_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29841));   // verilog/coms.v(128[12] 303[6])
    defparam i15765_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2122_3_lut (.I0(n3119), 
            .I1(n3186), .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15766_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29842));   // verilog/coms.v(128[12] 303[6])
    defparam i15766_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2120_3_lut (.I0(n3117), 
            .I1(n3184), .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15767_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29843));   // verilog/coms.v(128[12] 303[6])
    defparam i15767_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2113_3_lut (.I0(n3110), 
            .I1(n3177), .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15217_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position_scaled[16]), 
            .I2(n24373), .I3(GND_net), .O(n29293));   // verilog/coms.v(128[12] 303[6])
    defparam i15217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15768_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29844));   // verilog/coms.v(128[12] 303[6])
    defparam i15768_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2112_3_lut (.I0(n3109), 
            .I1(n3176), .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2111_3_lut (.I0(n3108), 
            .I1(n3175), .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2117_3_lut (.I0(n3114), 
            .I1(n3181), .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2115_3_lut (.I0(n3112), 
            .I1(n3179), .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2114_3_lut (.I0(n3111), 
            .I1(n3178), .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2134_3_lut (.I0(n3131), 
            .I1(n3198), .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2133_3_lut (.I0(n3130), 
            .I1(n3197), .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position_scaled_23__N_327[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5648));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2121_3_lut (.I0(n3118), 
            .I1(n3185), .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15218_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n24373), .I3(GND_net), .O(n29294));   // verilog/coms.v(128[12] 303[6])
    defparam i15218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15769_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29845));   // verilog/coms.v(128[12] 303[6])
    defparam i15769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2119_3_lut (.I0(n3116), 
            .I1(n3183), .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15770_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29846));   // verilog/coms.v(128[12] 303[6])
    defparam i15770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2118_3_lut (.I0(n3115), 
            .I1(n3182), .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2132_3_lut (.I0(n3129), 
            .I1(n3196), .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15771_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29847));   // verilog/coms.v(128[12] 303[6])
    defparam i15771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15772_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29848));   // verilog/coms.v(128[12] 303[6])
    defparam i15772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2127_3_lut (.I0(n3124), 
            .I1(n3191), .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2131_3_lut (.I0(n3128), 
            .I1(n3195), .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15773_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29849));   // verilog/coms.v(128[12] 303[6])
    defparam i15773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2126_3_lut (.I0(n3123), 
            .I1(n3190), .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15774_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29850));   // verilog/coms.v(128[12] 303[6])
    defparam i15774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2128_3_lut (.I0(n3125), 
            .I1(n3192), .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2130_3_lut (.I0(n3127), 
            .I1(n3194), .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15219_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n24373), .I3(GND_net), .O(n29295));   // verilog/coms.v(128[12] 303[6])
    defparam i15219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15775_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29851));   // verilog/coms.v(128[12] 303[6])
    defparam i15775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2124_3_lut (.I0(n3121), 
            .I1(n3188), .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15776_3_lut (.I0(\data_in_frame[23] [7]), .I1(rx_data[7]), 
            .I2(n48638), .I3(GND_net), .O(n29852));   // verilog/coms.v(128[12] 303[6])
    defparam i15776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1722_3_lut (.I0(n2527), 
            .I1(n2594), .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15339_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n50602), 
            .I3(GND_net), .O(n29415));   // verilog/coms.v(128[12] 303[6])
    defparam i15339_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_16 (.CI(n43787), 
            .I0(n2620), .I1(VCC_net), .CO(n43788));
    SB_CARRY add_1039_2 (.CI(GND_net), .I0(n4904), .I1(n4929), .CO(n43318));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_12_lut (.I0(n56181), 
            .I1(n1224), .I2(VCC_net), .I3(n43552), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_175_25 (.CI(n43178), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n43179));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_15_lut (.I0(GND_net), 
            .I1(n2621), .I2(VCC_net), .I3(n43786), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_15 (.CI(n43786), 
            .I0(n2621), .I1(VCC_net), .CO(n43787));
    SB_LUT4 add_175_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n43177), .O(n1541)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_11_lut (.I0(GND_net), 
            .I1(n1225), .I2(VCC_net), .I3(n43551), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_14_lut (.I0(GND_net), 
            .I1(n2622), .I2(VCC_net), .I3(n43785), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_24 (.CI(n43177), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n43178));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_11 (.CI(n43551), 
            .I0(n1225), .I1(VCC_net), .CO(n43552));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_14 (.CI(n43785), 
            .I0(n2622), .I1(VCC_net), .CO(n43786));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_10_lut (.I0(GND_net), 
            .I1(n1226), .I2(VCC_net), .I3(n43550), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_13_lut (.I0(GND_net), 
            .I1(n2623), .I2(VCC_net), .I3(n43784), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n43176), .O(n1542)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_23 (.CI(n43176), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n43177));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_13 (.CI(n43784), 
            .I0(n2623), .I1(VCC_net), .CO(n43785));
    SB_LUT4 add_263_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n43083), .O(encoder1_position_scaled_23__N_75[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_12_lut (.I0(GND_net), 
            .I1(n2624), .I2(VCC_net), .I3(n43783), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_12 (.CI(n43783), 
            .I0(n2624), .I1(VCC_net), .CO(n43784));
    SB_CARRY add_261_15 (.CI(n43116), .I0(duty[16]), .I1(n56288), .CO(n43117));
    SB_LUT4 add_261_14_lut (.I0(current[15]), .I1(duty[15]), .I2(n56288), 
            .I3(n43115), .O(n258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_14_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_10 (.CI(n43550), 
            .I0(n1226), .I1(VCC_net), .CO(n43551));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_9_lut (.I0(GND_net), 
            .I1(n1227), .I2(VCC_net), .I3(n43549), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2125_3_lut (.I0(n3122), 
            .I1(n3189), .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_263_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n43091), .O(encoder1_position_scaled_23__N_75[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n43175), .O(n1543)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2129_3_lut (.I0(n3126), 
            .I1(n3193), .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2137_3_lut (.I0(n542), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15777_3_lut (.I0(\data_in_frame[23] [6]), .I1(rx_data[6]), 
            .I2(n48638), .I3(GND_net), .O(n29853));   // verilog/coms.v(128[12] 303[6])
    defparam i15777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15778_3_lut (.I0(\data_in_frame[23] [5]), .I1(rx_data[5]), 
            .I2(n48638), .I3(GND_net), .O(n29854));   // verilog/coms.v(128[12] 303[6])
    defparam i15778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2136_3_lut (.I0(n3133), 
            .I1(n3200), .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15779_3_lut (.I0(\data_in_frame[23] [4]), .I1(rx_data[4]), 
            .I2(n48638), .I3(GND_net), .O(n29855));   // verilog/coms.v(128[12] 303[6])
    defparam i15779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2135_3_lut (.I0(n3132), 
            .I1(n3199), .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_11_lut (.I0(GND_net), 
            .I1(n2625), .I2(VCC_net), .I3(n43782), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_14 (.CI(n43115), .I0(duty[15]), .I1(n56288), .CO(n43116));
    SB_CARRY add_175_22 (.CI(n43175), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n43176));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position_scaled_23__N_327[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5647));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15780_3_lut (.I0(\data_in_frame[23] [3]), .I1(rx_data[3]), 
            .I2(n48638), .I3(GND_net), .O(n29856));   // verilog/coms.v(128[12] 303[6])
    defparam i15780_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_263_5 (.CI(n43083), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n43084));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i2_3_lut (.I0(encoder0_position_scaled_23__N_327[1]), 
            .I1(n32), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n543));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_11 (.CI(n43782), 
            .I0(n2625), .I1(VCC_net), .CO(n43783));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_10_lut (.I0(GND_net), 
            .I1(n2626), .I2(VCC_net), .I3(n43781), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1511_3_lut (.I0(n2220), 
            .I1(n2287), .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_10 (.CI(n43781), 
            .I0(n2626), .I1(VCC_net), .CO(n43782));
    SB_LUT4 add_175_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n43174), .O(n1544)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40477_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56270));
    defparam i40477_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_9_lut (.I0(GND_net), 
            .I1(n2627), .I2(VCC_net), .I3(n43780), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_9 (.CI(n43780), 
            .I0(n2627), .I1(VCC_net), .CO(n43781));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_8_lut (.I0(GND_net), 
            .I1(n2628), .I2(VCC_net), .I3(n43779), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_9 (.CI(n43549), 
            .I0(n1227), .I1(VCC_net), .CO(n43550));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_8_lut (.I0(GND_net), 
            .I1(n1228), .I2(VCC_net), .I3(n43548), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_8 (.CI(n43548), 
            .I0(n1228), .I1(VCC_net), .CO(n43549));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_8 (.CI(n43779), 
            .I0(n2628), .I1(VCC_net), .CO(n43780));
    SB_LUT4 i22624_4_lut (.I0(n543), .I1(n3231), .I2(n3232), .I3(n3233), 
            .O(n36694));
    defparam i22624_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_7_lut (.I0(GND_net), 
            .I1(n2629), .I2(GND_net), .I3(n43778), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_7 (.CI(n43778), 
            .I0(n2629), .I1(GND_net), .CO(n43779));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_6_lut (.I0(GND_net), 
            .I1(n2630), .I2(GND_net), .I3(n43777), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1756 (.I0(n3225), .I1(n3221), .I2(n3220), .I3(GND_net), 
            .O(n51948));
    defparam i1_3_lut_adj_1756.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1757 (.I0(n3226), .I1(n3224), .I2(n3222), .I3(n3227), 
            .O(n51962));
    defparam i1_4_lut_adj_1757.LUT_INIT = 16'hfffe;
    SB_LUT4 i15781_3_lut (.I0(\data_in_frame[23] [2]), .I1(rx_data[2]), 
            .I2(n48638), .I3(GND_net), .O(n29857));   // verilog/coms.v(128[12] 303[6])
    defparam i15781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1758 (.I0(n51962), .I1(n3223), .I2(n3228), .I3(GND_net), 
            .O(n51964));
    defparam i1_3_lut_adj_1758.LUT_INIT = 16'hfefe;
    SB_CARRY add_175_21 (.CI(n43174), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n43175));
    SB_LUT4 i1_4_lut_adj_1759 (.I0(n3214), .I1(n3215), .I2(n3217), .I3(n51964), 
            .O(n51970));
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 i15782_3_lut (.I0(\data_in_frame[23] [1]), .I1(rx_data[1]), 
            .I2(n48638), .I3(GND_net), .O(n29858));   // verilog/coms.v(128[12] 303[6])
    defparam i15782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(n3210), .I1(n3211), .I2(n3213), .I3(n51970), 
            .O(n51976));
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 i15567_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n50620), .I3(GND_net), .O(n29643));   // verilog/coms.v(128[12] 303[6])
    defparam i15567_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15568_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n50620), .I3(GND_net), .O(n29644));   // verilog/coms.v(128[12] 303[6])
    defparam i15568_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_6 (.CI(n43777), 
            .I0(n2630), .I1(GND_net), .CO(n43778));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_5_lut (.I0(GND_net), 
            .I1(n2631), .I2(VCC_net), .I3(n43776), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n43173), .O(n1545)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_5 (.CI(n43776), 
            .I0(n2631), .I1(VCC_net), .CO(n43777));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_4_lut (.I0(GND_net), 
            .I1(n2632), .I2(GND_net), .I3(n43775), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_4 (.CI(n43775), 
            .I0(n2632), .I1(GND_net), .CO(n43776));
    SB_LUT4 i40419_4_lut (.I0(n1026), .I1(n49689), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i40419_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15340_3_lut (.I0(deadband[23]), .I1(\data_in_frame[14] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29416));   // verilog/coms.v(128[12] 303[6])
    defparam i15340_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15569_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n50620), .I3(GND_net), .O(n29645));   // verilog/coms.v(128[12] 303[6])
    defparam i15569_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_3_lut (.I0(GND_net), 
            .I1(n2633), .I2(VCC_net), .I3(n43774), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15570_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n50620), .I3(GND_net), .O(n29646));   // verilog/coms.v(128[12] 303[6])
    defparam i15570_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15571_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[15]), .I2(n35803), 
            .I3(n27287), .O(n29647));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15571_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_7_lut (.I0(GND_net), 
            .I1(n1229), .I2(GND_net), .I3(n43547), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_7 (.CI(n43547), 
            .I0(n1229), .I1(GND_net), .CO(n43548));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_3 (.CI(n43774), 
            .I0(n2633), .I1(VCC_net), .CO(n43775));
    SB_CARRY add_175_20 (.CI(n43173), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n43174));
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n3229), .I1(n51948), .I2(n36694), .I3(n3230), 
            .O(n51950));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'heccc;
    SB_LUT4 i15572_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n50620), .I3(GND_net), .O(n29648));   // verilog/coms.v(128[12] 303[6])
    defparam i15572_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_6_lut (.I0(GND_net), 
            .I1(n1230), .I2(GND_net), .I3(n43546), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15783_3_lut (.I0(\data_in_frame[23] [0]), .I1(rx_data[0]), 
            .I2(n48638), .I3(GND_net), .O(n29859));   // verilog/coms.v(128[12] 303[6])
    defparam i15783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position_scaled_23__N_327[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5646));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15573_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n50620), .I3(GND_net), .O(n29649));   // verilog/coms.v(128[12] 303[6])
    defparam i15573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1762 (.I0(n3216), .I1(n3218), .I2(n3219), .I3(GND_net), 
            .O(n52004));
    defparam i1_3_lut_adj_1762.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1771_2_lut (.I0(GND_net), 
            .I1(n537), .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i641_3_lut (.I0(n520), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1578_3_lut (.I0(n2319), 
            .I1(n2386), .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n51976), 
            .O(n51982));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'hfffe;
    SB_LUT4 i22666_4_lut (.I0(n522), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n36736));
    defparam i22666_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1645_3_lut (.I0(n2418), 
            .I1(n2485), .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15574_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n50620), .I3(GND_net), .O(n29650));   // verilog/coms.v(128[12] 303[6])
    defparam i15574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n3205), .I1(n52004), .I2(n51950), .I3(n3212), 
            .O(n51954));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hfffe;
    SB_LUT4 i15575_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n50620), .I3(GND_net), .O(n29651));   // verilog/coms.v(128[12] 303[6])
    defparam i15575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40481_4_lut (.I0(n3206), .I1(n51954), .I2(n51982), .I3(n3204), 
            .O(n3237));
    defparam i40481_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15576_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n50620), .I3(GND_net), .O(n29652));   // verilog/coms.v(128[12] 303[6])
    defparam i15576_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1771_2 (.CI(VCC_net), 
            .I0(n537), .I1(GND_net), .CO(n43774));
    SB_LUT4 add_175_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n43172), .O(n1546)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2045_3_lut (.I0(n3010), 
            .I1(n3077), .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i13_3_lut (.I0(encoder0_position_scaled_23__N_327[12]), 
            .I1(n21_adj_5490), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n532));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_6 (.CI(n43546), 
            .I0(n1230), .I1(GND_net), .CO(n43547));
    SB_LUT4 i40388_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56181));
    defparam i40388_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15577_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n50620), .I3(GND_net), .O(n29653));   // verilog/coms.v(128[12] 303[6])
    defparam i15577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_5_lut (.I0(GND_net), 
            .I1(n1231), .I2(VCC_net), .I3(n43545), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_5 (.CI(n43545), 
            .I0(n1231), .I1(VCC_net), .CO(n43546));
    SB_LUT4 i15578_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n50620), .I3(GND_net), .O(n29654));   // verilog/coms.v(128[12] 303[6])
    defparam i15578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_25_lut (.I0(n55883), 
            .I1(n2511), .I2(VCC_net), .I3(n43773), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_4_lut (.I0(GND_net), 
            .I1(n1232), .I2(GND_net), .I3(n43544), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2044_3_lut (.I0(n3009), 
            .I1(n3076), .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_19 (.CI(n43172), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n43173));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2043_3_lut (.I0(n3008), 
            .I1(n3075), .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15579_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n50620), .I3(GND_net), .O(n29655));   // verilog/coms.v(128[12] 303[6])
    defparam i15579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_24_lut (.I0(GND_net), 
            .I1(n2512), .I2(VCC_net), .I3(n43772), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_24 (.CI(n43772), 
            .I0(n2512), .I1(VCC_net), .CO(n43773));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_23_lut (.I0(GND_net), 
            .I1(n2513), .I2(VCC_net), .I3(n43771), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_4 (.CI(n43544), 
            .I0(n1232), .I1(GND_net), .CO(n43545));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_3_lut (.I0(GND_net), 
            .I1(n1233), .I2(VCC_net), .I3(n43543), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_3 (.CI(n43543), 
            .I0(n1233), .I1(VCC_net), .CO(n43544));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_833_2_lut (.I0(GND_net), 
            .I1(n523), .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position_scaled_23__N_327[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5645));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15580_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n50620), .I3(GND_net), .O(n29656));   // verilog/coms.v(128[12] 303[6])
    defparam i15580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2041_3_lut (.I0(n3006), 
            .I1(n3073), .I2(n3039), .I3(GND_net), .O(n3105));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15581_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n50620), .I3(GND_net), .O(n29657));   // verilog/coms.v(128[12] 303[6])
    defparam i15581_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_23 (.CI(n43771), 
            .I0(n2513), .I1(VCC_net), .CO(n43772));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2042_rep_35_3_lut (.I0(n3007), 
            .I1(n3074), .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2042_rep_35_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_22_lut (.I0(GND_net), 
            .I1(n2514), .I2(VCC_net), .I3(n43770), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_22 (.CI(n43770), 
            .I0(n2514), .I1(VCC_net), .CO(n43771));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2049_3_lut (.I0(n3014), 
            .I1(n3081), .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15582_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n50620), .I3(GND_net), .O(n29658));   // verilog/coms.v(128[12] 303[6])
    defparam i15582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_175_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n43171), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2048_3_lut (.I0(n3013), 
            .I1(n3080), .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_21_lut (.I0(GND_net), 
            .I1(n2515), .I2(VCC_net), .I3(n43769), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2046_rep_53_3_lut (.I0(n3011), 
            .I1(n3078), .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2046_rep_53_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15583_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n50620), .I3(GND_net), .O(n29659));   // verilog/coms.v(128[12] 303[6])
    defparam i15583_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_21 (.CI(n43769), 
            .I0(n2515), .I1(VCC_net), .CO(n43770));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_20_lut (.I0(GND_net), 
            .I1(n2516), .I2(VCC_net), .I3(n43768), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_20 (.CI(n43768), 
            .I0(n2516), .I1(VCC_net), .CO(n43769));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_19_lut (.I0(GND_net), 
            .I1(n2517), .I2(VCC_net), .I3(n43767), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_19 (.CI(n43767), 
            .I0(n2517), .I1(VCC_net), .CO(n43768));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_18_lut (.I0(GND_net), 
            .I1(n2518), .I2(VCC_net), .I3(n43766), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15584_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n50620), .I3(GND_net), .O(n29660));   // verilog/coms.v(128[12] 303[6])
    defparam i15584_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_833_2 (.CI(VCC_net), 
            .I0(n523), .I1(GND_net), .CO(n43543));
    SB_LUT4 add_261_13_lut (.I0(current[11]), .I1(duty[14]), .I2(n56288), 
            .I3(n43114), .O(n259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_13_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_3_lut_adj_1765 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n51394));
    defparam i1_3_lut_adj_1765.LUT_INIT = 16'hfefe;
    SB_LUT4 i15585_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n50620), .I3(GND_net), .O(n29661));   // verilog/coms.v(128[12] 303[6])
    defparam i15585_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_18 (.CI(n43171), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n43172));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_18 (.CI(n43766), 
            .I0(n2518), .I1(VCC_net), .CO(n43767));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2047_3_lut (.I0(n3012), 
            .I1(n3079), .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15586_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n50620), .I3(GND_net), .O(n29662));   // verilog/coms.v(128[12] 303[6])
    defparam i15586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1457_3_lut (.I0(n532), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233_adj_5612));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_17_lut (.I0(GND_net), 
            .I1(n2519), .I2(VCC_net), .I3(n43765), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2051_3_lut (.I0(n3016), 
            .I1(n3083), .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1766 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n51644));
    defparam i1_2_lut_adj_1766.LUT_INIT = 16'h8888;
    SB_LUT4 add_261_16_lut (.I0(current[15]), .I1(duty[17]), .I2(n56288), 
            .I3(n43117), .O(n256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_16_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_175_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n43170), .O(n1548)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15587_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n50620), .I3(GND_net), .O(n29663));   // verilog/coms.v(128[12] 303[6])
    defparam i15587_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_17 (.CI(n43170), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n43171));
    SB_LUT4 i15588_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n50620), .I3(GND_net), .O(n29664));   // verilog/coms.v(128[12] 303[6])
    defparam i15588_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_17 (.CI(n43765), 
            .I0(n2519), .I1(VCC_net), .CO(n43766));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_16_lut (.I0(GND_net), 
            .I1(n2520), .I2(VCC_net), .I3(n43764), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i40406_4_lut (.I0(n51644), .I1(n1125), .I2(n51394), .I3(n36736), 
            .O(n1158));
    defparam i40406_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 add_175_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n43169), .O(n1549)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_11_lut (.I0(n56195), 
            .I1(n1125), .I2(VCC_net), .I3(n43542), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2052_3_lut (.I0(n3017), 
            .I1(n3084), .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2050_3_lut (.I0(n3015), 
            .I1(n3082), .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_263_13 (.CI(n43091), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n43092));
    SB_LUT4 i15589_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n50620), .I3(GND_net), .O(n29665));   // verilog/coms.v(128[12] 303[6])
    defparam i15589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2059_3_lut (.I0(n3024), 
            .I1(n3091), .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2062_3_lut (.I0(n3027), 
            .I1(n3094), .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_16 (.CI(n43764), 
            .I0(n2520), .I1(VCC_net), .CO(n43765));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_15_lut (.I0(GND_net), 
            .I1(n2521), .I2(VCC_net), .I3(n43763), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15590_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n50620), .I3(GND_net), .O(n29666));   // verilog/coms.v(128[12] 303[6])
    defparam i15590_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_15 (.CI(n43763), 
            .I0(n2521), .I1(VCC_net), .CO(n43764));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_14_lut (.I0(GND_net), 
            .I1(n2522), .I2(VCC_net), .I3(n43762), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2061_3_lut (.I0(n3026), 
            .I1(n3093), .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_261_13 (.CI(n43114), .I0(duty[14]), .I1(n56288), .CO(n43115));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2069_3_lut (.I0(n541), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15791_3_lut (.I0(\data_out_frame[21] [6]), .I1(current[15]), 
            .I2(n24373), .I3(GND_net), .O(n29867));   // verilog/coms.v(128[12] 303[6])
    defparam i15791_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_175_16 (.CI(n43169), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n43170));
    SB_LUT4 i15591_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n49594), .I3(GND_net), .O(n29667));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_263_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n43082), .O(encoder1_position_scaled_23__N_75[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2068_3_lut (.I0(n3033), 
            .I1(n3100), .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position_scaled_23__N_327[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5644));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15592_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n49594), .I3(GND_net), .O(n29668));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i3_3_lut (.I0(encoder0_position_scaled_23__N_327[2]), 
            .I1(n31), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n542));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2060_3_lut (.I0(n3025), 
            .I1(n3092), .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2054_3_lut (.I0(n3019), 
            .I1(n3086), .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15593_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n49594), .I3(GND_net), .O(n29669));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15593_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_14 (.CI(n43762), 
            .I0(n2522), .I1(VCC_net), .CO(n43763));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2053_3_lut (.I0(n3018), 
            .I1(n3085), .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15792_3_lut (.I0(\data_out_frame[21] [5]), .I1(current[15]), 
            .I2(n24373), .I3(GND_net), .O(n29868));   // verilog/coms.v(128[12] 303[6])
    defparam i15792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15594_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n49594), .I3(GND_net), .O(n29670));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15594_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15793_3_lut (.I0(\data_out_frame[21] [4]), .I1(current[15]), 
            .I2(n24373), .I3(GND_net), .O(n29869));   // verilog/coms.v(128[12] 303[6])
    defparam i15793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_13_lut (.I0(GND_net), 
            .I1(n2523), .I2(VCC_net), .I3(n43761), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2067_3_lut (.I0(n3032), 
            .I1(n3099), .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22598_3_lut (.I0(n523), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n36668));
    defparam i22598_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2066_3_lut (.I0(n3031), 
            .I1(n3098), .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15595_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n49594), .I3(GND_net), .O(n29671));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15595_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_13 (.CI(n43761), 
            .I0(n2523), .I1(VCC_net), .CO(n43762));
    SB_LUT4 i15794_3_lut (.I0(\data_out_frame[21] [3]), .I1(current[11]), 
            .I2(n24373), .I3(GND_net), .O(n29870));   // verilog/coms.v(128[12] 303[6])
    defparam i15794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15596_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n49594), .I3(GND_net), .O(n29672));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15596_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15597_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n49594), .I3(GND_net), .O(n29673));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15597_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15598_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n49594), .I3(GND_net), .O(n29674));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15598_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2065_3_lut (.I0(n3030), 
            .I1(n3097), .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5516));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15795_3_lut (.I0(\data_out_frame[21] [2]), .I1(current[10]), 
            .I2(n24373), .I3(GND_net), .O(n29871));   // verilog/coms.v(128[12] 303[6])
    defparam i15795_3_lut.LUT_INIT = 16'hcaca;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2055_3_lut (.I0(n3020), 
            .I1(n3087), .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2056_3_lut (.I0(n3021), 
            .I1(n3088), .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_263_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n43090), .O(encoder1_position_scaled_23__N_75[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position_scaled_23__N_327[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5643));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15599_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n49594), .I3(GND_net), .O(n29675));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15599_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_10_lut (.I0(GND_net), 
            .I1(n1126), .I2(VCC_net), .I3(n43541), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15600_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n49594), .I3(GND_net), .O(n29676));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15600_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_12_lut (.I0(GND_net), 
            .I1(n2524), .I2(VCC_net), .I3(n43760), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2063_3_lut (.I0(n3028), 
            .I1(n3095), .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15796_3_lut (.I0(\data_out_frame[21] [1]), .I1(current[9]), 
            .I2(n24373), .I3(GND_net), .O(n29872));   // verilog/coms.v(128[12] 303[6])
    defparam i15796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15797_3_lut (.I0(\data_out_frame[21] [0]), .I1(current[8]), 
            .I2(n24373), .I3(GND_net), .O(n29873));   // verilog/coms.v(128[12] 303[6])
    defparam i15797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2058_3_lut (.I0(n3023), 
            .I1(n3090), .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1767 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n51662));
    defparam i1_3_lut_adj_1767.LUT_INIT = 16'hfefe;
    SB_LUT4 i15601_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n49594), .I3(GND_net), .O(n29677));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15601_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_10 (.CI(n43541), 
            .I0(n1126), .I1(VCC_net), .CO(n43542));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_12 (.CI(n43760), 
            .I0(n2524), .I1(VCC_net), .CO(n43761));
    SB_LUT4 i15602_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n49594), .I3(GND_net), .O(n29678));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15602_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_11_lut (.I0(GND_net), 
            .I1(n2525), .I2(VCC_net), .I3(n43759), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15603_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n49594), .I3(GND_net), .O(n29679));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15603_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_11 (.CI(n43759), 
            .I0(n2525), .I1(VCC_net), .CO(n43760));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_10_lut (.I0(GND_net), 
            .I1(n2526), .I2(VCC_net), .I3(n43758), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n47754));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF read_221 (.Q(read), .C(clk16MHz), .D(n51212));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_9_lut (.I0(GND_net), 
            .I1(n1127), .I2(VCC_net), .I3(n43540), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_10 (.CI(n43758), 
            .I0(n2526), .I1(VCC_net), .CO(n43759));
    SB_LUT4 i1_4_lut_adj_1768 (.I0(n1229), .I1(n36668), .I2(n1230), .I3(n1231), 
            .O(n49684));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_9_lut (.I0(GND_net), 
            .I1(n2527), .I2(VCC_net), .I3(n43757), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2064_3_lut (.I0(n3029), 
            .I1(n3096), .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1524_3_lut (.I0(n2233_adj_5612), 
            .I1(n2300), .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_9 (.CI(n43757), 
            .I0(n2527), .I1(VCC_net), .CO(n43758));
    SB_LUT4 i15798_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n24373), .I3(GND_net), .O(n29874));   // verilog/coms.v(128[12] 303[6])
    defparam i15798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15604_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n49594), .I3(GND_net), .O(n29680));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15604_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2057_3_lut (.I0(n3022), 
            .I1(n3089), .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_8_lut (.I0(GND_net), 
            .I1(n2528), .I2(VCC_net), .I3(n43756), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_8 (.CI(n43756), 
            .I0(n2528), .I1(VCC_net), .CO(n43757));
    SB_LUT4 i15799_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n24373), .I3(GND_net), .O(n29875));   // verilog/coms.v(128[12] 303[6])
    defparam i15799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15605_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n49594), .I3(GND_net), .O(n29681));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15605_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15341_3_lut (.I0(deadband[22]), .I1(\data_in_frame[14] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29417));   // verilog/coms.v(128[12] 303[6])
    defparam i15341_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15606_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n49594), .I3(GND_net), .O(n29682));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15606_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15800_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n24373), .I3(GND_net), .O(n29876));   // verilog/coms.v(128[12] 303[6])
    defparam i15800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1037_i1_4_lut (.I0(n54231), .I1(duty[0]), .I2(n296), .I3(n356), 
            .O(n4929));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam mux_1037_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position_scaled_23__N_327[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5642));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15801_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n24373), .I3(GND_net), .O(n29877));   // verilog/coms.v(128[12] 303[6])
    defparam i15801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n3121), .I1(n3128), .I2(n3122), .I3(n3127), 
            .O(n51334));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_LUT4 i15607_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n49594), .I3(GND_net), .O(n29683));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15607_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15608_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n49594), .I3(GND_net), .O(n29684));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15608_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15802_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n24373), .I3(GND_net), .O(n29878));   // verilog/coms.v(128[12] 303[6])
    defparam i15802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15342_3_lut (.I0(deadband[21]), .I1(\data_in_frame[14] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29418));   // verilog/coms.v(128[12] 303[6])
    defparam i15342_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15609_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n24373), .I3(GND_net), .O(n29685));   // verilog/coms.v(128[12] 303[6])
    defparam i15609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22560_3_lut (.I0(n542), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n36630));
    defparam i22560_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15610_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n24373), .I3(GND_net), .O(n29686));   // verilog/coms.v(128[12] 303[6])
    defparam i15610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15611_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n24373), .I3(GND_net), .O(n29687));   // verilog/coms.v(128[12] 303[6])
    defparam i15611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1770 (.I0(n3120), .I1(n3119), .I2(GND_net), .I3(GND_net), 
            .O(n51708));
    defparam i1_2_lut_adj_1770.LUT_INIT = 16'heeee;
    SB_LUT4 i40392_4_lut (.I0(n1225), .I1(n1224), .I2(n49684), .I3(n51662), 
            .O(n1257));
    defparam i40392_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15803_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n24373), .I3(GND_net), .O(n29879));   // verilog/coms.v(128[12] 303[6])
    defparam i15803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1591_3_lut (.I0(n2332), 
            .I1(n2399), .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15612_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n49594), .I3(GND_net), .O(n29688));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15612_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15804_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n24373), .I3(GND_net), .O(n29880));   // verilog/coms.v(128[12] 303[6])
    defparam i15804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15613_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n49594), .I3(GND_net), .O(n29689));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15613_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(n3129), .I1(n36630), .I2(n3130), .I3(n3131), 
            .O(n49790));
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'ha080;
    SB_LUT4 i15805_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n24373), .I3(GND_net), .O(n29881));   // verilog/coms.v(128[12] 303[6])
    defparam i15805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n3117), .I1(n51334), .I2(n3118), .I3(n3124), 
            .O(n51338));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1773 (.I0(n3125), .I1(n3126), .I2(n3123), .I3(GND_net), 
            .O(n51988));
    defparam i1_3_lut_adj_1773.LUT_INIT = 16'hfefe;
    SB_LUT4 i15614_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n49594), .I3(GND_net), .O(n29690));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15614_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14967_2_lut (.I0(n28583), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n29049));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i14967_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39783_4_lut (.I0(commutation_state[1]), .I1(n24565), .I2(dti), 
            .I3(commutation_state[2]), .O(n28583));
    defparam i39783_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i15615_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n49594), .I3(GND_net), .O(n29691));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15615_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15616_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n49594), .I3(GND_net), .O(n29692));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15616_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n3114), .I1(n51988), .I2(n51338), .I3(n3116), 
            .O(n51342));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'hfffe;
    SB_LUT4 i15220_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n24373), .I3(GND_net), .O(n29296));   // verilog/coms.v(128[12] 303[6])
    defparam i15220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15617_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n49594), .I3(GND_net), .O(n29693));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15617_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(n3115), .I1(n3111), .I2(n49790), .I3(n51708), 
            .O(n50867));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n3110), .I1(n3112), .I2(n3113), .I3(n51342), 
            .O(n51348));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'hfffe;
    SB_LUT4 i15221_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n24373), .I3(GND_net), .O(n29297));   // verilog/coms.v(128[12] 303[6])
    defparam i15221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15222_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n24373), .I3(GND_net), .O(n29298));   // verilog/coms.v(128[12] 303[6])
    defparam i15222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15618_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n49594), .I3(GND_net), .O(n29694));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15618_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15223_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n24373), .I3(GND_net), .O(n29299));   // verilog/coms.v(128[12] 303[6])
    defparam i15223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n3108), .I1(n3109), .I2(n51348), .I3(n50867), 
            .O(n51354));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_LUT4 i15619_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n49594), .I3(GND_net), .O(n29695));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15619_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15224_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n24373), .I3(GND_net), .O(n29300));   // verilog/coms.v(128[12] 303[6])
    defparam i15224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15225_3_lut (.I0(current[0]), .I1(data_adj_5722[0]), .I2(n28640), 
            .I3(GND_net), .O(n29301));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39934_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n51354), 
            .O(n3138));
    defparam i39934_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1778 (.I0(enable_slow_N_4393), .I1(data_ready), 
            .I2(state_adj_5716[1]), .I3(state_adj_5716[0]), .O(n48368));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hccd0;
    SB_LUT4 i15620_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n49594), .I3(GND_net), .O(n29696));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15620_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15227_4_lut (.I0(rw), .I1(state_adj_5716[0]), .I2(state_adj_5716[1]), 
            .I3(n6272), .O(n29303));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15227_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i15621_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n49594), .I3(GND_net), .O(n29697));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15621_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1980_3_lut (.I0(n2913), 
            .I1(n2980), .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15228_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n24373), .I3(GND_net), .O(n29304));   // verilog/coms.v(128[12] 303[6])
    defparam i15228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1979_3_lut (.I0(n2912), 
            .I1(n2979), .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15229_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n24373), .I3(GND_net), .O(n29305));   // verilog/coms.v(128[12] 303[6])
    defparam i15229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15230_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n24373), .I3(GND_net), .O(n29306));   // verilog/coms.v(128[12] 303[6])
    defparam i15230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15231_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n24373), .I3(GND_net), .O(n29307));   // verilog/coms.v(128[12] 303[6])
    defparam i15231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15232_3_lut (.I0(CS_c), .I1(state_adj_5724[0]), .I2(state_adj_5724[1]), 
            .I3(GND_net), .O(n29308));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15232_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1977_3_lut (.I0(n2910), 
            .I1(n2977), .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40490_4_lut (.I0(n15_adj_5481), .I1(clk_out), .I2(state_adj_5724[0]), 
            .I3(state_adj_5724[1]), .O(n9_adj_5511));   // verilog/tli4970.v(35[10] 68[6])
    defparam i40490_4_lut.LUT_INIT = 16'hc8fc;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_7_lut (.I0(GND_net), 
            .I1(n2529), .I2(GND_net), .I3(n43755), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15622_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n49594), .I3(GND_net), .O(n29698));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15622_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1975_3_lut (.I0(n2908), 
            .I1(n2975), .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15623_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n49594), .I3(GND_net), .O(n29699));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15623_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1994_3_lut (.I0(n2927), 
            .I1(n2994), .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15234_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n24373), .I3(GND_net), .O(n29310));   // verilog/coms.v(128[12] 303[6])
    defparam i15234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1986_3_lut (.I0(n2919), 
            .I1(n2986), .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15235_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n24373), .I3(GND_net), .O(n29311));   // verilog/coms.v(128[12] 303[6])
    defparam i15235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15624_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n49594), .I3(GND_net), .O(n29700));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15624_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15236_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n24373), .I3(GND_net), .O(n29312));   // verilog/coms.v(128[12] 303[6])
    defparam i15236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15237_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n24373), .I3(GND_net), .O(n29313));   // verilog/coms.v(128[12] 303[6])
    defparam i15237_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_9 (.CI(n43540), 
            .I0(n1127), .I1(VCC_net), .CO(n43541));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_8_lut (.I0(GND_net), 
            .I1(n1128), .I2(VCC_net), .I3(n43539), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_7 (.CI(n43755), 
            .I0(n2529), .I1(GND_net), .CO(n43756));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_8 (.CI(n43539), 
            .I0(n1128), .I1(VCC_net), .CO(n43540));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_7_lut (.I0(GND_net), 
            .I1(n1129), .I2(GND_net), .I3(n43538), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15238_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n24373), .I3(GND_net), .O(n29314));   // verilog/coms.v(128[12] 303[6])
    defparam i15238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_175_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n43168), .O(n1550)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_6_lut (.I0(GND_net), 
            .I1(n2530), .I2(GND_net), .I3(n43754), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_15 (.CI(n43168), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n43169));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1985_3_lut (.I0(n2918), 
            .I1(n2985), .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15239_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n24373), .I3(GND_net), .O(n29315));   // verilog/coms.v(128[12] 303[6])
    defparam i15239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15625_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n24373), .I3(GND_net), .O(n29701));   // verilog/coms.v(128[12] 303[6])
    defparam i15625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1984_3_lut (.I0(n2917), 
            .I1(n2984), .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15626_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n24373), .I3(GND_net), .O(n29702));   // verilog/coms.v(128[12] 303[6])
    defparam i15626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1982_3_lut (.I0(n2915), 
            .I1(n2982), .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15240_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n24373), .I3(GND_net), .O(n29316));   // verilog/coms.v(128[12] 303[6])
    defparam i15240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15627_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n24373), .I3(GND_net), .O(n29703));   // verilog/coms.v(128[12] 303[6])
    defparam i15627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15241_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[11]), .I2(n35841), 
            .I3(n27222), .O(n29317));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15241_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_6 (.CI(n43754), 
            .I0(n2530), .I1(GND_net), .CO(n43755));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1978_3_lut (.I0(n2911), 
            .I1(n2978), .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15628_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n24373), .I3(GND_net), .O(n29704));   // verilog/coms.v(128[12] 303[6])
    defparam i15628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15242_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n24373), .I3(GND_net), .O(n29318));   // verilog/coms.v(128[12] 303[6])
    defparam i15242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15243_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n24373), .I3(GND_net), .O(n29319));   // verilog/coms.v(128[12] 303[6])
    defparam i15243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15629_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n24373), .I3(GND_net), .O(n29705));   // verilog/coms.v(128[12] 303[6])
    defparam i15629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1976_3_lut (.I0(n2909), 
            .I1(n2976), .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15630_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n24373), .I3(GND_net), .O(n29706));   // verilog/coms.v(128[12] 303[6])
    defparam i15630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15631_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n24373), .I3(GND_net), .O(n29707));   // verilog/coms.v(128[12] 303[6])
    defparam i15631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1983_3_lut (.I0(n2916), 
            .I1(n2983), .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1981_3_lut (.I0(n2914), 
            .I1(n2981), .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_261_12_lut (.I0(current[10]), .I1(duty[13]), .I2(n56288), 
            .I3(n43113), .O(n260)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_12_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i15632_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n51220), .I3(GND_net), 
            .O(n29708));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15632_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1988_3_lut (.I0(n2921), 
            .I1(n2988), .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1992_3_lut (.I0(n2925), 
            .I1(n2992), .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15633_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n51220), .I3(GND_net), 
            .O(n29709));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15633_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_5_lut (.I0(GND_net), 
            .I1(n2531), .I2(VCC_net), .I3(n43753), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1996_3_lut (.I0(n2929), 
            .I1(n2996), .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15634_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n51220), .I3(GND_net), 
            .O(n29710));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2001_3_lut (.I0(n540), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15635_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n51220), .I3(GND_net), 
            .O(n29711));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15635_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_5 (.CI(n43753), 
            .I0(n2531), .I1(VCC_net), .CO(n43754));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_4_lut (.I0(GND_net), 
            .I1(n2532), .I2(GND_net), .I3(n43752), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1658_3_lut (.I0(n2431), 
            .I1(n2498), .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15636_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n51220), .I3(GND_net), 
            .O(n29712));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15636_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_4 (.CI(n43752), 
            .I0(n2532), .I1(GND_net), .CO(n43753));
    SB_CARRY add_261_12 (.CI(n43113), .I0(duty[13]), .I1(n56288), .CO(n43114));
    SB_LUT4 i33748_3_lut (.I0(n6_adj_5505), .I1(n8588), .I2(n49468), .I3(GND_net), 
            .O(n49475));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_261_11_lut (.I0(current[9]), .I1(duty[12]), .I2(n56288), 
            .I3(n43112), .O(n261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_11_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_7 (.CI(n43538), 
            .I0(n1129), .I1(GND_net), .CO(n43539));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_3_lut (.I0(GND_net), 
            .I1(n2533), .I2(VCC_net), .I3(n43751), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_6_lut (.I0(GND_net), 
            .I1(n1130), .I2(GND_net), .I3(n43537), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15637_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n51220), .I3(GND_net), 
            .O(n29713));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15638_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n51220), .I3(GND_net), 
            .O(n29714));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15638_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22596_3_lut (.I0(n524), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n36666));
    defparam i22596_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i2000_3_lut (.I0(n2933), 
            .I1(n3000), .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i4_3_lut (.I0(encoder0_position_scaled_23__N_327[3]), 
            .I1(n30), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n541));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15640_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n24373), .I3(GND_net), .O(n29716));   // verilog/coms.v(128[12] 303[6])
    defparam i15640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15641_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n24373), .I3(GND_net), .O(n29717));   // verilog/coms.v(128[12] 303[6])
    defparam i15641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15642_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n24373), .I3(GND_net), .O(n29718));   // verilog/coms.v(128[12] 303[6])
    defparam i15642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15643_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n24373), .I3(GND_net), .O(n29719));   // verilog/coms.v(128[12] 303[6])
    defparam i15643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15644_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n24373), .I3(GND_net), .O(n29720));   // verilog/coms.v(128[12] 303[6])
    defparam i15644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15645_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n24373), .I3(GND_net), .O(n29721));   // verilog/coms.v(128[12] 303[6])
    defparam i15645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15646_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n24373), .I3(GND_net), .O(n29722));   // verilog/coms.v(128[12] 303[6])
    defparam i15646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1999_3_lut (.I0(n2932), 
            .I1(n2999), .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15647_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n24373), .I3(GND_net), .O(n29723));   // verilog/coms.v(128[12] 303[6])
    defparam i15647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15648_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n24373), .I3(GND_net), .O(n29724));   // verilog/coms.v(128[12] 303[6])
    defparam i15648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15649_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n24373), .I3(GND_net), .O(n29725));   // verilog/coms.v(128[12] 303[6])
    defparam i15649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1998_3_lut (.I0(n2931), 
            .I1(n2998), .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15650_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n24373), .I3(GND_net), .O(n29726));   // verilog/coms.v(128[12] 303[6])
    defparam i15650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15651_4_lut (.I0(state_7__N_4306[3]), .I1(data[0]), .I2(n10_adj_5617), 
            .I3(n27262), .O(n29727));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15651_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_3 (.CI(n43751), 
            .I0(n2533), .I1(VCC_net), .CO(n43752));
    SB_LUT4 i15660_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[1]), .I2(n6_adj_5571), 
            .I3(n27294), .O(n29736));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15660_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15664_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_5595), 
            .I3(n27232), .O(n29740));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15664_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15665_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[0]), .I2(n7_adj_5597), 
            .I3(state_7__N_4499), .O(n29741));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15665_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_18_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1997_3_lut (.I0(n2930), 
            .I1(n2997), .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15672_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_5478), 
            .I3(n27227), .O(n29748));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15672_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15673_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n35837), 
            .I3(n27232), .O(n29749));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15673_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1993_3_lut (.I0(n2926), 
            .I1(n2993), .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15674_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[2]), .I2(n6_adj_5571), 
            .I3(n27281), .O(n29750));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15674_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1990_3_lut (.I0(n2923), 
            .I1(n2990), .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15675_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n24373), .I3(GND_net), .O(n29751));   // verilog/coms.v(128[12] 303[6])
    defparam i15675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1987_3_lut (.I0(n2920), 
            .I1(n2987), .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1704_2_lut (.I0(GND_net), 
            .I1(n536), .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1989_3_lut (.I0(n2922), 
            .I1(n2989), .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1704_2 (.CI(VCC_net), 
            .I0(n536), .I1(GND_net), .CO(n43751));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1991_3_lut (.I0(n2924), 
            .I1(n2991), .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_24_lut (.I0(GND_net), 
            .I1(n2412), .I2(VCC_net), .I3(n43750), .O(n2479)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_6 (.CI(n43537), 
            .I0(n1130), .I1(GND_net), .CO(n43538));
    SB_LUT4 i15676_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n24373), .I3(GND_net), .O(n29752));   // verilog/coms.v(128[12] 303[6])
    defparam i15676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1995_3_lut (.I0(n2928), 
            .I1(n2995), .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_23_lut (.I0(GND_net), 
            .I1(n2413), .I2(VCC_net), .I3(n43749), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_23 (.CI(n43749), 
            .I0(n2413), .I1(VCC_net), .CO(n43750));
    SB_LUT4 i15244_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[12]), .I2(n35803), 
            .I3(n27256), .O(n29320));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15244_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_5_lut (.I0(GND_net), 
            .I1(n1131), .I2(VCC_net), .I3(n43536), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15677_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n24373), .I3(GND_net), .O(n29753));   // verilog/coms.v(128[12] 303[6])
    defparam i15677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39963_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55756));
    defparam i39963_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15678_3_lut (.I0(\data_out_frame[22] [7]), .I1(current[7]), 
            .I2(n24373), .I3(GND_net), .O(n29754));   // verilog/coms.v(128[12] 303[6])
    defparam i15678_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_5 (.CI(n43536), 
            .I0(n1131), .I1(VCC_net), .CO(n43537));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_22_lut (.I0(GND_net), 
            .I1(n2414), .I2(VCC_net), .I3(n43748), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_22 (.CI(n43748), 
            .I0(n2414), .I1(VCC_net), .CO(n43749));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_21_lut (.I0(GND_net), 
            .I1(n2415), .I2(VCC_net), .I3(n43747), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33749_3_lut (.I0(encoder0_position_scaled_23__N_327[27]), .I1(n49475), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22562_3_lut (.I0(n541), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n36632));
    defparam i22562_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_21 (.CI(n43747), 
            .I0(n2415), .I1(VCC_net), .CO(n43748));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_20_lut (.I0(GND_net), 
            .I1(n2416), .I2(VCC_net), .I3(n43746), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n1324), .I1(n1323), .I2(n1327), .I3(n1328), 
            .O(n50654));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_20 (.CI(n43746), 
            .I0(n2416), .I1(VCC_net), .CO(n43747));
    SB_LUT4 add_175_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n43167), .O(n1551)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_19_lut (.I0(GND_net), 
            .I1(n2417), .I2(VCC_net), .I3(n43745), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15679_3_lut (.I0(\data_out_frame[22] [6]), .I1(current[6]), 
            .I2(n24373), .I3(GND_net), .O(n29755));   // verilog/coms.v(128[12] 303[6])
    defparam i15679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1780 (.I0(n1329), .I1(n36666), .I2(n1330), .I3(n1331), 
            .O(n49681));
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_19 (.CI(n43745), 
            .I0(n2417), .I1(VCC_net), .CO(n43746));
    SB_LUT4 i40377_4_lut (.I0(n49681), .I1(n50654), .I2(n1325), .I3(n1326), 
            .O(n1356));
    defparam i40377_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15680_3_lut (.I0(\data_out_frame[22] [5]), .I1(current[5]), 
            .I2(n24373), .I3(GND_net), .O(n29756));   // verilog/coms.v(128[12] 303[6])
    defparam i15680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_18_lut (.I0(GND_net), 
            .I1(n2418), .I2(VCC_net), .I3(n43744), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1781 (.I0(n3027), .I1(n3023), .I2(n3021), .I3(n3019), 
            .O(n51908));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1782 (.I0(n3028), .I1(n3024), .I2(n3020), .I3(GND_net), 
            .O(n51906));
    defparam i1_3_lut_adj_1782.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15681_3_lut (.I0(\data_out_frame[22] [4]), .I1(current[4]), 
            .I2(n24373), .I3(GND_net), .O(n29757));   // verilog/coms.v(128[12] 303[6])
    defparam i15681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1783 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n51672));
    defparam i1_2_lut_adj_1783.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_18 (.CI(n43744), 
            .I0(n2418), .I1(VCC_net), .CO(n43745));
    SB_CARRY add_175_14 (.CI(n43167), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n43168));
    SB_LUT4 i1_4_lut_adj_1784 (.I0(n51906), .I1(n51908), .I2(n3022), .I3(n3025), 
            .O(n51912));
    defparam i1_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_4_lut (.I0(GND_net), 
            .I1(n1132), .I2(GND_net), .I3(n43535), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_17_lut (.I0(GND_net), 
            .I1(n2419), .I2(VCC_net), .I3(n43743), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_17 (.CI(n43743), 
            .I0(n2419), .I1(VCC_net), .CO(n43744));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_4 (.CI(n43535), 
            .I0(n1132), .I1(GND_net), .CO(n43536));
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n3029), .I1(n36632), .I2(n3030), .I3(n3031), 
            .O(n49830));
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'ha080;
    SB_LUT4 i15682_3_lut (.I0(\data_out_frame[22] [3]), .I1(current[3]), 
            .I2(n24373), .I3(GND_net), .O(n29758));   // verilog/coms.v(128[12] 303[6])
    defparam i15682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_16_lut (.I0(GND_net), 
            .I1(n2420), .I2(VCC_net), .I3(n43742), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15683_3_lut (.I0(\data_out_frame[22] [2]), .I1(current[2]), 
            .I2(n24373), .I3(GND_net), .O(n29759));   // verilog/coms.v(128[12] 303[6])
    defparam i15683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15684_3_lut (.I0(\data_out_frame[22] [1]), .I1(current[1]), 
            .I2(n24373), .I3(GND_net), .O(n29760));   // verilog/coms.v(128[12] 303[6])
    defparam i15684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position_scaled_23__N_327[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5641));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n3013), .I1(n3015), .I2(n49830), .I3(n51912), 
            .O(n51918));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'hfffe;
    SB_LUT4 i15685_3_lut (.I0(\data_out_frame[22] [0]), .I1(current[0]), 
            .I2(n24373), .I3(GND_net), .O(n29761));   // verilog/coms.v(128[12] 303[6])
    defparam i15685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15686_3_lut (.I0(\data_out_frame[21] [7]), .I1(current[15]), 
            .I2(n24373), .I3(GND_net), .O(n29762));   // verilog/coms.v(128[12] 303[6])
    defparam i15686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15687_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[3]), .I2(n6_adj_5571), 
            .I3(n27287), .O(n29763));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15687_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(n3016), .I1(n3017), .I2(n3018), .I3(n3026), 
            .O(n51932));
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_16 (.CI(n43742), 
            .I0(n2420), .I1(VCC_net), .CO(n43743));
    SB_LUT4 i1_4_lut_adj_1788 (.I0(hall3), .I1(commutation_state[1]), .I2(hall2), 
            .I3(hall1), .O(n48472));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'hd054;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_3_lut (.I0(GND_net), 
            .I1(n1133), .I2(VCC_net), .I3(n43534), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_15_lut (.I0(GND_net), 
            .I1(n2421), .I2(VCC_net), .I3(n43741), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i15690_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_5595), 
            .I3(n27227), .O(n29766));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15690_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i22594_3_lut (.I0(n525), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n36664));
    defparam i22594_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_15 (.CI(n43741), 
            .I0(n2421), .I1(VCC_net), .CO(n43742));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_14_lut (.I0(GND_net), 
            .I1(n2422), .I2(VCC_net), .I3(n43740), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_14 (.CI(n43740), 
            .I0(n2422), .I1(VCC_net), .CO(n43741));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_13_lut (.I0(GND_net), 
            .I1(n2423), .I2(VCC_net), .I3(n43739), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_13 (.CI(n43739), 
            .I0(n2423), .I1(VCC_net), .CO(n43740));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i839_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_3 (.CI(n43534), 
            .I0(n1133), .I1(VCC_net), .CO(n43535));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_12_lut (.I0(GND_net), 
            .I1(n2424), .I2(VCC_net), .I3(n43738), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15691_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_5539), 
            .I3(n27232), .O(n29767));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15691_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15692_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[4]), .I2(n6_adj_5537), 
            .I3(n27256), .O(n29768));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15692_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n51672), 
            .O(n51678));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_LUT4 i15693_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_5539), 
            .I3(n27227), .O(n29769));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15693_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15694_3_lut (.I0(current[11]), .I1(data_adj_5722[11]), .I2(n28640), 
            .I3(GND_net), .O(n29770));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n3009), .I1(n3011), .I2(n3012), .I3(n51918), 
            .O(n51924));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_12 (.CI(n43738), 
            .I0(n2424), .I1(VCC_net), .CO(n43739));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_11_lut (.I0(GND_net), 
            .I1(n2425), .I2(VCC_net), .I3(n43737), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(n1429), .I1(n36664), .I2(n1430), .I3(n1431), 
            .O(n49699));
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'ha080;
    SB_LUT4 i15695_3_lut (.I0(current[10]), .I1(data_adj_5722[10]), .I2(n28640), 
            .I3(GND_net), .O(n29771));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15695_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_11 (.CI(n43737), 
            .I0(n2425), .I1(VCC_net), .CO(n43738));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_766_2_lut (.I0(GND_net), 
            .I1(n522), .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_766_2 (.CI(VCC_net), 
            .I0(n522), .I1(GND_net), .CO(n43534));
    SB_LUT4 i1_4_lut_adj_1792 (.I0(n3008), .I1(n3010), .I2(n3014), .I3(n51932), 
            .O(n51938));
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_10_lut (.I0(GND_net), 
            .I1(n2426), .I2(VCC_net), .I3(n43736), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39967_4_lut (.I0(n3007), .I1(n51938), .I2(n51924), .I3(n3006), 
            .O(n3039));
    defparam i39967_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15696_3_lut (.I0(current[9]), .I1(data_adj_5722[9]), .I2(n28640), 
            .I3(GND_net), .O(n29772));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15697_3_lut (.I0(current[8]), .I1(data_adj_5722[8]), .I2(n28640), 
            .I3(GND_net), .O(n29773));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15697_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_10 (.CI(n43736), 
            .I0(n2426), .I1(VCC_net), .CO(n43737));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_9_lut (.I0(GND_net), 
            .I1(n2427), .I2(VCC_net), .I3(n43735), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15698_3_lut (.I0(current[7]), .I1(data_adj_5722[7]), .I2(n28640), 
            .I3(GND_net), .O(n29774));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15699_3_lut (.I0(current[6]), .I1(data_adj_5722[6]), .I2(n28640), 
            .I3(GND_net), .O(n29775));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15700_3_lut (.I0(current[5]), .I1(data_adj_5722[5]), .I2(n28640), 
            .I3(GND_net), .O(n29776));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15701_3_lut (.I0(current[4]), .I1(data_adj_5722[4]), .I2(n28640), 
            .I3(GND_net), .O(n29777));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15702_3_lut (.I0(current[3]), .I1(data_adj_5722[3]), .I2(n28640), 
            .I3(GND_net), .O(n29778));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15702_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_9 (.CI(n43735), 
            .I0(n2427), .I1(VCC_net), .CO(n43736));
    SB_LUT4 i15703_3_lut (.I0(current[2]), .I1(data_adj_5722[2]), .I2(n28640), 
            .I3(GND_net), .O(n29779));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15704_3_lut (.I0(current[1]), .I1(data_adj_5722[1]), .I2(n28640), 
            .I3(GND_net), .O(n29780));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_8_lut (.I0(GND_net), 
            .I1(n2428), .I2(VCC_net), .I3(n43734), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_8 (.CI(n43734), 
            .I0(n2428), .I1(VCC_net), .CO(n43735));
    SB_LUT4 i15705_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[5]), .I2(n6_adj_5537), 
            .I3(n27294), .O(n29781));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15705_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15706_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(\PID_CONTROLLER.integral_23__N_3996 [23]), 
            .I2(control_update), .I3(GND_net), .O(n29782));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40361_4_lut (.I0(n49699), .I1(n1422), .I2(n1423), .I3(n51678), 
            .O(n1455));
    defparam i40361_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_7_lut (.I0(GND_net), 
            .I1(n2429), .I2(GND_net), .I3(n43733), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15707_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(\PID_CONTROLLER.integral_23__N_3996 [22]), 
            .I2(control_update), .I3(GND_net), .O(n29783));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_10_lut (.I0(GND_net), 
            .I1(n1026), .I2(VCC_net), .I3(n43533), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position_scaled_23__N_327[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5640));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5517));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_7 (.CI(n43733), 
            .I0(n2429), .I1(GND_net), .CO(n43734));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position_scaled_23__N_327[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5639));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_6_lut (.I0(GND_net), 
            .I1(n2430), .I2(GND_net), .I3(n43732), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_6 (.CI(n43732), 
            .I0(n2430), .I1(GND_net), .CO(n43733));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_9_lut (.I0(GND_net), 
            .I1(n1027), .I2(VCC_net), .I3(n43532), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1040_3_lut (.I0(n1525), 
            .I1(n1592), .I2(n1554_adj_5610), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_5_lut (.I0(GND_net), 
            .I1(n2431), .I2(VCC_net), .I3(n43731), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_5 (.CI(n43731), 
            .I0(n2431), .I1(VCC_net), .CO(n43732));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_4_lut (.I0(GND_net), 
            .I1(n2432), .I2(GND_net), .I3(n43730), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position_scaled_23__N_327[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5638));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_4 (.CI(n43730), 
            .I0(n2432), .I1(GND_net), .CO(n43731));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_9 (.CI(n43532), 
            .I0(n1027), .I1(VCC_net), .CO(n43533));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22658_4_lut (.I0(n526), .I1(n1531), .I2(n1532_adj_5608), 
            .I3(n1533_adj_5609), .O(n36728));
    defparam i22658_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1107_3_lut (.I0(n1624), 
            .I1(n1691), .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1793 (.I0(n1525), .I1(n1526), .I2(n1527), .I3(n1528), 
            .O(n51402));
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1174_3_lut (.I0(n1723), 
            .I1(n1790), .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1794 (.I0(n1529), .I1(n1530), .I2(GND_net), .I3(GND_net), 
            .O(n51684));
    defparam i1_2_lut_adj_1794.LUT_INIT = 16'h8888;
    SB_LUT4 i15806_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n24373), .I3(GND_net), .O(n29882));   // verilog/coms.v(128[12] 303[6])
    defparam i15806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1909_3_lut (.I0(n2810), 
            .I1(n2877), .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_8_lut (.I0(GND_net), 
            .I1(n1028), .I2(VCC_net), .I3(n43531), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position_scaled_23__N_327[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5637));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1241_3_lut (.I0(n1822), 
            .I1(n1889), .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1908_3_lut (.I0(n2809), 
            .I1(n2876), .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1912_3_lut (.I0(n2813), 
            .I1(n2880), .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1911_3_lut (.I0(n2812), 
            .I1(n2879), .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5518));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position_scaled_23__N_327[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5636));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15807_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n24373), .I3(GND_net), .O(n29883));   // verilog/coms.v(128[12] 303[6])
    defparam i15807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position_scaled_23__N_327[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5635));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15808_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n24373), .I3(GND_net), .O(n29884));   // verilog/coms.v(128[12] 303[6])
    defparam i15808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1910_3_lut (.I0(n2811), 
            .I1(n2878), .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_3_lut (.I0(GND_net), 
            .I1(n2433), .I2(VCC_net), .I3(n43729), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_8 (.CI(n43531), 
            .I0(n1028), .I1(VCC_net), .CO(n43532));
    SB_LUT4 i15708_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral_23__N_3996 [21]), 
            .I2(control_update), .I3(GND_net), .O(n29784));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39995_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55788));
    defparam i39995_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_3 (.CI(n43729), 
            .I0(n2433), .I1(VCC_net), .CO(n43730));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1637_2_lut (.I0(GND_net), 
            .I1(n535), .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1637_2 (.CI(VCC_net), 
            .I0(n535), .I1(GND_net), .CO(n43729));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_23_lut (.I0(n55960), 
            .I1(n2313), .I2(VCC_net), .I3(n43728), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n1524), .I1(n51684), .I2(n51402), .I3(n36728), 
            .O(n51406));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_22_lut (.I0(GND_net), 
            .I1(n2314), .I2(VCC_net), .I3(n43727), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position_scaled_23__N_327[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5634));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_22 (.CI(n43727), 
            .I0(n2314), .I1(VCC_net), .CO(n43728));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_21_lut (.I0(GND_net), 
            .I1(n2315), .I2(VCC_net), .I3(n43726), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1915_3_lut (.I0(n2816), 
            .I1(n2883), .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_7_lut (.I0(GND_net), 
            .I1(n1029), .I2(GND_net), .I3(n43530), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15809_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n24373), .I3(GND_net), .O(n29885));   // verilog/coms.v(128[12] 303[6])
    defparam i15809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5463));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15810_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n24373), .I3(GND_net), .O(n29886));   // verilog/coms.v(128[12] 303[6])
    defparam i15810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15811_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n24373), .I3(GND_net), .O(n29887));   // verilog/coms.v(128[12] 303[6])
    defparam i15811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position_scaled_23__N_327[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5633));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40327_1_lut (.I0(n1554_adj_5610), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n56120));
    defparam i40327_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_21 (.CI(n43726), 
            .I0(n2315), .I1(VCC_net), .CO(n43727));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position_scaled_23__N_327[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5632));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_20_lut (.I0(GND_net), 
            .I1(n2316), .I2(VCC_net), .I3(n43725), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1914_3_lut (.I0(n2815), 
            .I1(n2882), .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15812_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n24373), .I3(GND_net), .O(n29888));   // verilog/coms.v(128[12] 303[6])
    defparam i15812_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_20 (.CI(n43725), 
            .I0(n2316), .I1(VCC_net), .CO(n43726));
    SB_LUT4 i15813_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n24373), .I3(GND_net), .O(n29889));   // verilog/coms.v(128[12] 303[6])
    defparam i15813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1913_3_lut (.I0(n2814), 
            .I1(n2881), .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15814_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n24373), .I3(GND_net), .O(n29890));   // verilog/coms.v(128[12] 303[6])
    defparam i15814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1919_3_lut (.I0(n2820), 
            .I1(n2887), .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15709_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .I2(control_update), .I3(GND_net), .O(n29785));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15815_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n24373), .I3(GND_net), .O(n29891));   // verilog/coms.v(128[12] 303[6])
    defparam i15815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15816_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n24373), .I3(GND_net), .O(n29892));   // verilog/coms.v(128[12] 303[6])
    defparam i15816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15817_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n24373), .I3(GND_net), .O(n29893));   // verilog/coms.v(128[12] 303[6])
    defparam i15817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15710_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(control_update), .I3(GND_net), .O(n29786));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1308_rep_19_3_lut (.I0(n1921), 
            .I1(n1988), .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1308_rep_19_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1375_3_lut (.I0(n2020), 
            .I1(n2087), .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15818_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n24373), .I3(GND_net), .O(n29894));   // verilog/coms.v(128[12] 303[6])
    defparam i15818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1918_3_lut (.I0(n2819), 
            .I1(n2886), .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1933_3_lut (.I0(n539), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1932_3_lut (.I0(n2833), 
            .I1(n2900), .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15819_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n24373), .I3(GND_net), .O(n29895));   // verilog/coms.v(128[12] 303[6])
    defparam i15819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position_scaled_23__N_327[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5631));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15820_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n24373), .I3(GND_net), .O(n29896));   // verilog/coms.v(128[12] 303[6])
    defparam i15820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15821_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n24373), .I3(GND_net), .O(n29897));   // verilog/coms.v(128[12] 303[6])
    defparam i15821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i40344_4_lut (.I0(n1522), .I1(n1521), .I2(n1523), .I3(n51406), 
            .O(n1554_adj_5610));
    defparam i40344_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15711_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(control_update), .I3(GND_net), .O(n29787));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15712_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(control_update), .I3(GND_net), .O(n29788));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1442_3_lut (.I0(n2119), 
            .I1(n2186), .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i5_3_lut (.I0(encoder0_position_scaled_23__N_327[4]), 
            .I1(n29), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n540));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1928_3_lut (.I0(n2829), 
            .I1(n2896), .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15822_3_lut (.I0(\data_out_frame[17] [7]), .I1(pwm_setpoint[7]), 
            .I2(n24373), .I3(GND_net), .O(n29898));   // verilog/coms.v(128[12] 303[6])
    defparam i15822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15713_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(control_update), .I3(GND_net), .O(n29789));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_19_lut (.I0(GND_net), 
            .I1(n2317), .I2(VCC_net), .I3(n43724), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_19 (.CI(n43724), 
            .I0(n2317), .I1(VCC_net), .CO(n43725));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_18_lut (.I0(GND_net), 
            .I1(n2318), .I2(VCC_net), .I3(n43723), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15823_3_lut (.I0(\data_out_frame[17] [6]), .I1(pwm_setpoint[6]), 
            .I2(n24373), .I3(GND_net), .O(n29899));   // verilog/coms.v(128[12] 303[6])
    defparam i15823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position_scaled_23__N_327[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5630));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15824_3_lut (.I0(\data_out_frame[17] [5]), .I1(pwm_setpoint[5]), 
            .I2(n24373), .I3(GND_net), .O(n29900));   // verilog/coms.v(128[12] 303[6])
    defparam i15824_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_7 (.CI(n43530), 
            .I0(n1029), .I1(GND_net), .CO(n43531));
    SB_LUT4 i15825_3_lut (.I0(\data_out_frame[17] [4]), .I1(pwm_setpoint[4]), 
            .I2(n24373), .I3(GND_net), .O(n29901));   // verilog/coms.v(128[12] 303[6])
    defparam i15825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15826_3_lut (.I0(\data_out_frame[17] [3]), .I1(pwm_setpoint[3]), 
            .I2(n24373), .I3(GND_net), .O(n29902));   // verilog/coms.v(128[12] 303[6])
    defparam i15826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position_scaled_23__N_327[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5629));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15714_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(control_update), .I3(GND_net), .O(n29790));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15715_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(control_update), .I3(GND_net), .O(n29791));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15716_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(control_update), .I3(GND_net), .O(n29792));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1920_3_lut (.I0(n2821), 
            .I1(n2888), .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1509_3_lut (.I0(n2218), 
            .I1(n2285), .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position_scaled_23__N_327[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5628));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position_scaled_23__N_327[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5627));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1926_3_lut (.I0(n2827), 
            .I1(n2894), .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15827_3_lut (.I0(\data_out_frame[17] [2]), .I1(pwm_setpoint[2]), 
            .I2(n24373), .I3(GND_net), .O(n29903));   // verilog/coms.v(128[12] 303[6])
    defparam i15827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15828_3_lut (.I0(\data_out_frame[17] [1]), .I1(pwm_setpoint[1]), 
            .I2(n24373), .I3(GND_net), .O(n29904));   // verilog/coms.v(128[12] 303[6])
    defparam i15828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_6_lut (.I0(GND_net), 
            .I1(n1030), .I2(GND_net), .I3(n43529), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1925_3_lut (.I0(n2826), 
            .I1(n2893), .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_18 (.CI(n43723), 
            .I0(n2318), .I1(VCC_net), .CO(n43724));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_17_lut (.I0(GND_net), 
            .I1(n2319), .I2(VCC_net), .I3(n43722), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_17 (.CI(n43722), 
            .I0(n2319), .I1(VCC_net), .CO(n43723));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1927_3_lut (.I0(n2828), 
            .I1(n2895), .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1923_3_lut (.I0(n2824), 
            .I1(n2891), .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15717_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(control_update), .I3(GND_net), .O(n29793));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5519));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1921_3_lut (.I0(n2822), 
            .I1(n2889), .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1917_3_lut (.I0(n2818), 
            .I1(n2885), .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15718_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(control_update), .I3(GND_net), .O(n29794));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1916_3_lut (.I0(n2817), 
            .I1(n2884), .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_6 (.CI(n43529), 
            .I0(n1030), .I1(GND_net), .CO(n43530));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_5_lut (.I0(GND_net), 
            .I1(n1031), .I2(VCC_net), .I3(n43528), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_5 (.CI(n43528), 
            .I0(n1031), .I1(VCC_net), .CO(n43529));
    SB_LUT4 i15719_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(control_update), .I3(GND_net), .O(n29795));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position_scaled_23__N_327[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5626));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1931_3_lut (.I0(n2832), 
            .I1(n2899), .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_16_lut (.I0(GND_net), 
            .I1(n2320), .I2(VCC_net), .I3(n43721), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_16 (.CI(n43721), 
            .I0(n2320), .I1(VCC_net), .CO(n43722));
    SB_LUT4 i15829_3_lut (.I0(\data_out_frame[17] [0]), .I1(pwm_setpoint[0]), 
            .I2(n24373), .I3(GND_net), .O(n29905));   // verilog/coms.v(128[12] 303[6])
    defparam i15829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1930_3_lut (.I0(n2831), 
            .I1(n2898), .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5520));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1929_3_lut (.I0(n2830), 
            .I1(n2897), .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position_scaled_23__N_327[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5625));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_175_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n43166), .O(n1552)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_15_lut (.I0(GND_net), 
            .I1(n2321), .I2(VCC_net), .I3(n43720), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_15 (.CI(n43720), 
            .I0(n2321), .I1(VCC_net), .CO(n43721));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1922_3_lut (.I0(n2823), 
            .I1(n2890), .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_14_lut (.I0(GND_net), 
            .I1(n2322), .I2(VCC_net), .I3(n43719), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_14 (.CI(n43719), 
            .I0(n2322), .I1(VCC_net), .CO(n43720));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_4_lut (.I0(GND_net), 
            .I1(n1032), .I2(GND_net), .I3(n43527), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15830_3_lut (.I0(\data_out_frame[16] [7]), .I1(pwm_setpoint[15]), 
            .I2(n24373), .I3(GND_net), .O(n29906));   // verilog/coms.v(128[12] 303[6])
    defparam i15830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15831_3_lut (.I0(\data_out_frame[16] [6]), .I1(pwm_setpoint[14]), 
            .I2(n24373), .I3(GND_net), .O(n29907));   // verilog/coms.v(128[12] 303[6])
    defparam i15831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_13_lut (.I0(GND_net), 
            .I1(n2323), .I2(VCC_net), .I3(n43718), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_13 (.CI(n43718), 
            .I0(n2323), .I1(VCC_net), .CO(n43719));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_4 (.CI(n43527), 
            .I0(n1032), .I1(GND_net), .CO(n43528));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_3_lut (.I0(GND_net), 
            .I1(n1033), .I2(VCC_net), .I3(n43526), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_12_lut (.I0(GND_net), 
            .I1(n2324), .I2(VCC_net), .I3(n43717), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1924_3_lut (.I0(n2825), 
            .I1(n2892), .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_3 (.CI(n43526), 
            .I0(n1033), .I1(VCC_net), .CO(n43527));
    SB_LUT4 i15832_3_lut (.I0(\data_out_frame[16] [5]), .I1(pwm_setpoint[13]), 
            .I2(n24373), .I3(GND_net), .O(n29908));   // verilog/coms.v(128[12] 303[6])
    defparam i15832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15833_3_lut (.I0(\data_out_frame[16] [4]), .I1(pwm_setpoint[12]), 
            .I2(n24373), .I3(GND_net), .O(n29909));   // verilog/coms.v(128[12] 303[6])
    defparam i15833_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_12 (.CI(n43717), 
            .I0(n2324), .I1(VCC_net), .CO(n43718));
    SB_LUT4 i15834_3_lut (.I0(\data_out_frame[16] [3]), .I1(pwm_setpoint[11]), 
            .I2(n24373), .I3(GND_net), .O(n29910));   // verilog/coms.v(128[12] 303[6])
    defparam i15834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_699_2_lut (.I0(GND_net), 
            .I1(n521), .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15720_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(control_update), .I3(GND_net), .O(n29796));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_11_lut (.I0(GND_net), 
            .I1(n2325), .I2(VCC_net), .I3(n43716), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(n2921), .I1(n2923), .I2(n2927), .I3(n2925), 
            .O(n51592));
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_11 (.CI(n43716), 
            .I0(n2325), .I1(VCC_net), .CO(n43717));
    SB_LUT4 i1_3_lut_adj_1797 (.I0(n2926), .I1(n2920), .I2(n2928), .I3(GND_net), 
            .O(n51590));
    defparam i1_3_lut_adj_1797.LUT_INIT = 16'hfefe;
    SB_LUT4 i15835_3_lut (.I0(\data_out_frame[16] [2]), .I1(pwm_setpoint[10]), 
            .I2(n24373), .I3(GND_net), .O(n29911));   // verilog/coms.v(128[12] 303[6])
    defparam i15835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_10_lut (.I0(GND_net), 
            .I1(n2326), .I2(VCC_net), .I3(n43715), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_13 (.CI(n43166), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n43167));
    SB_LUT4 i15721_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(control_update), .I3(GND_net), .O(n29797));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15721_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_10 (.CI(n43715), 
            .I0(n2326), .I1(VCC_net), .CO(n43716));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_9_lut (.I0(GND_net), 
            .I1(n2327), .I2(VCC_net), .I3(n43714), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15722_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(control_update), .I3(GND_net), .O(n29798));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5462));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position_scaled_23__N_327[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5624));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1798 (.I0(n51592), .I1(n2924), .I2(n2922), .I3(GND_net), 
            .O(n51594));
    defparam i1_3_lut_adj_1798.LUT_INIT = 16'hfefe;
    SB_LUT4 i15836_3_lut (.I0(\data_out_frame[16] [1]), .I1(pwm_setpoint[9]), 
            .I2(n24373), .I3(GND_net), .O(n29912));   // verilog/coms.v(128[12] 303[6])
    defparam i15836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15837_3_lut (.I0(\data_out_frame[16] [0]), .I1(pwm_setpoint[8]), 
            .I2(n24373), .I3(GND_net), .O(n29913));   // verilog/coms.v(128[12] 303[6])
    defparam i15837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position_scaled_23__N_327[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5623));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22564_3_lut (.I0(n540), .I1(n2932), .I2(n2933), .I3(GND_net), 
            .O(n36634));
    defparam i22564_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15838_3_lut (.I0(\data_out_frame[15] [7]), .I1(pwm_setpoint[23]), 
            .I2(n24373), .I3(GND_net), .O(n29914));   // verilog/coms.v(128[12] 303[6])
    defparam i15838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1576_3_lut (.I0(n2317), 
            .I1(n2384), .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15839_3_lut (.I0(\data_out_frame[15] [6]), .I1(pwm_setpoint[22]), 
            .I2(n24373), .I3(GND_net), .O(n29915));   // verilog/coms.v(128[12] 303[6])
    defparam i15839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n2918), .I1(n51594), .I2(n2919), .I3(n51590), 
            .O(n51600));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5521));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15840_3_lut (.I0(\data_out_frame[15] [5]), .I1(pwm_setpoint[21]), 
            .I2(n24373), .I3(GND_net), .O(n29916));   // verilog/coms.v(128[12] 303[6])
    defparam i15840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15723_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(control_update), .I3(GND_net), .O(n29799));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22590_3_lut (.I0(n527), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n36660));
    defparam i22590_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(n2929), .I1(n36634), .I2(n2930), .I3(n2931), 
            .O(n49781));
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'ha080;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n27284), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_5457));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15841_3_lut (.I0(\data_out_frame[15] [4]), .I1(pwm_setpoint[20]), 
            .I2(n24373), .I3(GND_net), .O(n29917));   // verilog/coms.v(128[12] 303[6])
    defparam i15841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15842_3_lut (.I0(\data_out_frame[15] [3]), .I1(pwm_setpoint[19]), 
            .I2(n24373), .I3(GND_net), .O(n29918));   // verilog/coms.v(128[12] 303[6])
    defparam i15842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1801 (.I0(n1629), .I1(n36660), .I2(n1630), .I3(n1631), 
            .O(n49707));
    defparam i1_4_lut_adj_1801.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1802 (.I0(n2916), .I1(n2917), .I2(n49781), .I3(n51600), 
            .O(n51606));
    defparam i1_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n51606), 
            .O(n51612));
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'hfffe;
    SB_LUT4 i15843_3_lut (.I0(\data_out_frame[15] [2]), .I1(pwm_setpoint[18]), 
            .I2(n24373), .I3(GND_net), .O(n29919));   // verilog/coms.v(128[12] 303[6])
    defparam i15843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_18_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15844_3_lut (.I0(\data_out_frame[15] [1]), .I1(pwm_setpoint[17]), 
            .I2(n24373), .I3(GND_net), .O(n29920));   // verilog/coms.v(128[12] 303[6])
    defparam i15844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position_scaled_23__N_327[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5622));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5461));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1804 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n51612), 
            .O(n51618));
    defparam i1_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_18_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5460));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15845_3_lut (.I0(\data_out_frame[15] [0]), .I1(pwm_setpoint[16]), 
            .I2(n24373), .I3(GND_net), .O(n29921));   // verilog/coms.v(128[12] 303[6])
    defparam i15845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39999_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n51618), 
            .O(n2940));
    defparam i39999_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15846_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n24373), .I3(GND_net), .O(n29922));   // verilog/coms.v(128[12] 303[6])
    defparam i15846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15847_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n24373), .I3(GND_net), .O(n29923));   // verilog/coms.v(128[12] 303[6])
    defparam i15847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15848_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n24373), .I3(GND_net), .O(n29924));   // verilog/coms.v(128[12] 303[6])
    defparam i15848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1842_3_lut (.I0(n2711), 
            .I1(n2778), .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15724_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(control_update), .I3(GND_net), .O(n29800));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15725_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(control_update), .I3(GND_net), .O(n29801));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1841_3_lut (.I0(n2710), 
            .I1(n2777), .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15849_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n24373), .I3(GND_net), .O(n29925));   // verilog/coms.v(128[12] 303[6])
    defparam i15849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15850_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n24373), .I3(GND_net), .O(n29926));   // verilog/coms.v(128[12] 303[6])
    defparam i15850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15726_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(control_update), .I3(GND_net), .O(n29802));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15851_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n24373), .I3(GND_net), .O(n29927));   // verilog/coms.v(128[12] 303[6])
    defparam i15851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1847_3_lut (.I0(n2716), 
            .I1(n2783), .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15852_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n24373), .I3(GND_net), .O(n29928));   // verilog/coms.v(128[12] 303[6])
    defparam i15852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15853_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n24373), .I3(GND_net), .O(n29929));   // verilog/coms.v(128[12] 303[6])
    defparam i15853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1846_3_lut (.I0(n2715), 
            .I1(n2782), .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15854_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n24373), .I3(GND_net), .O(n29930));   // verilog/coms.v(128[12] 303[6])
    defparam i15854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15855_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n24373), .I3(GND_net), .O(n29931));   // verilog/coms.v(128[12] 303[6])
    defparam i15855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15856_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n24373), .I3(GND_net), .O(n29932));   // verilog/coms.v(128[12] 303[6])
    defparam i15856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1850_3_lut (.I0(n2719), 
            .I1(n2786), .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15857_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n24373), .I3(GND_net), .O(n29933));   // verilog/coms.v(128[12] 303[6])
    defparam i15857_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dti_counter_2279__i7 (.Q(dti_counter[7]), .C(clk16MHz), .D(n48));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i6 (.Q(dti_counter[6]), .C(clk16MHz), .D(n49));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i5 (.Q(dti_counter[5]), .C(clk16MHz), .D(n50));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i4 (.Q(dti_counter[4]), .C(clk16MHz), .D(n51));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i3 (.Q(dti_counter[3]), .C(clk16MHz), .D(n52));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i2 (.Q(dti_counter[2]), .C(clk16MHz), .D(n53));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF dti_counter_2279__i1 (.Q(dti_counter[1]), .C(clk16MHz), .D(n54));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 i33750_3_lut (.I0(n7_adj_5504), .I1(n8589), .I2(n49468), .I3(GND_net), 
            .O(n49477));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33751_rep_33_3_lut (.I0(encoder0_position_scaled_23__N_327[26]), 
            .I1(n900), .I2(n861), .I3(GND_net), .O(n52838));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33751_rep_33_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n10832_bdd_4_lut (.I0(n10832), .I1(n418), .I2(current[15]), 
            .I3(duty[23]), .O(n56554));
    defparam n10832_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1021_1_lut (.I0(n296), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n4748));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1021_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n56554_bdd_3_lut (.I0(n56554), .I1(duty[23]), .I2(n249), .I3(GND_net), 
            .O(pwm_setpoint_23__N_11[23]));
    defparam n56554_bdd_3_lut.LUT_INIT = 16'h9898;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_9 (.CI(n43714), 
            .I0(n2327), .I1(VCC_net), .CO(n43715));
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n1624), .I1(n1626), .I2(n1627), .I3(n1628), 
            .O(n51696));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_8_lut (.I0(GND_net), 
            .I1(n2328), .I2(VCC_net), .I3(n43713), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_8 (.CI(n43713), 
            .I0(n2328), .I1(VCC_net), .CO(n43714));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position_scaled_23__N_327[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5621));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_7_lut (.I0(GND_net), 
            .I1(n2329), .I2(GND_net), .I3(n43712), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n49707), .I1(n1621), .I2(n1623), .I3(n1625), 
            .O(n50497));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_7 (.CI(n43712), 
            .I0(n2329), .I1(GND_net), .CO(n43713));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1849_3_lut (.I0(n2718), 
            .I1(n2785), .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_699_2 (.CI(VCC_net), 
            .I0(n521), .I1(GND_net), .CO(n43526));
    SB_LUT4 add_175_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n43165), .O(n1553)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_6_lut (.I0(GND_net), 
            .I1(n2330), .I2(GND_net), .I3(n43711), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15858_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n24373), .I3(GND_net), .O(n29934));   // verilog/coms.v(128[12] 303[6])
    defparam i15858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15859_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n24373), .I3(GND_net), .O(n29935));   // verilog/coms.v(128[12] 303[6])
    defparam i15859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i706_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_6 (.CI(n43711), 
            .I0(n2330), .I1(GND_net), .CO(n43712));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_5_lut (.I0(GND_net), 
            .I1(n2331), .I2(VCC_net), .I3(n43710), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_5 (.CI(n43710), 
            .I0(n2331), .I1(VCC_net), .CO(n43711));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_9_lut (.I0(n960), 
            .I1(n927), .I2(VCC_net), .I3(n43525), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_175_12 (.CI(n43165), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n43166));
    SB_LUT4 i15860_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n24373), .I3(GND_net), .O(n29936));   // verilog/coms.v(128[12] 303[6])
    defparam i15860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1848_3_lut (.I0(n2717), 
            .I1(n2784), .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_4_lut (.I0(GND_net), 
            .I1(n2332), .I2(GND_net), .I3(n43709), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_4 (.CI(n43709), 
            .I0(n2332), .I1(GND_net), .CO(n43710));
    SB_LUT4 i40326_4_lut (.I0(n1620), .I1(n50497), .I2(n1622), .I3(n51696), 
            .O(n1653));
    defparam i40326_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_3_lut (.I0(GND_net), 
            .I1(n2333), .I2(VCC_net), .I3(n43708), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_8_lut (.I0(GND_net), 
            .I1(n928), .I2(VCC_net), .I3(n43524), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15727_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(control_update), .I3(GND_net), .O(n29803));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i773_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_8 (.CI(n43524), 
            .I0(n928), .I1(VCC_net), .CO(n43525));
    SB_LUT4 i15861_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n24373), .I3(GND_net), .O(n29937));   // verilog/coms.v(128[12] 303[6])
    defparam i15861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15728_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(control_update), .I3(GND_net), .O(n29804));   // verilog/motorControl.v(43[14] 63[8])
    defparam i15728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_175_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n43164), .O(n1554)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_7_lut (.I0(GND_net), 
            .I1(n929), .I2(GND_net), .I3(n43523), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15729_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[6]), .I2(n6_adj_5537), 
            .I3(n27281), .O(n29805));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15729_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15862_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n24373), .I3(GND_net), .O(n29938));   // verilog/coms.v(128[12] 303[6])
    defparam i15862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_281_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[0]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i1_3_lut (.I0(encoder0_position_scaled[0]), .I1(motor_state_23__N_123[0]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i1_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_3 (.CI(n43708), 
            .I0(n2333), .I1(VCC_net), .CO(n43709));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_7 (.CI(n43523), 
            .I0(n929), .I1(GND_net), .CO(n43524));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1570_2_lut (.I0(GND_net), 
            .I1(n534), .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_6_lut (.I0(GND_net), 
            .I1(n930), .I2(GND_net), .I3(n43522), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_281_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[1]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_261_11 (.CI(n43112), .I0(duty[12]), .I1(n56288), .CO(n43113));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1570_2 (.CI(VCC_net), 
            .I0(n534), .I1(GND_net), .CO(n43708));
    SB_LUT4 add_261_10_lut (.I0(current[8]), .I1(duty[11]), .I2(n56288), 
            .I3(n43111), .O(n262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_10_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_6 (.CI(n43522), 
            .I0(n930), .I1(GND_net), .CO(n43523));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_22_lut (.I0(n55986), 
            .I1(n2214), .I2(VCC_net), .I3(n43707), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_21_lut (.I0(GND_net), 
            .I1(n2215), .I2(VCC_net), .I3(n43706), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_5_lut (.I0(GND_net), 
            .I1(n931), .I2(VCC_net), .I3(n43521), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_5 (.CI(n43521), 
            .I0(n931), .I1(VCC_net), .CO(n43522));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_4_lut (.I0(GND_net), 
            .I1(n932), .I2(GND_net), .I3(n43520), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_12 (.CI(n43090), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n43091));
    SB_CARRY add_175_11 (.CI(n43164), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n43165));
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_261_10 (.CI(n43111), .I0(duty[11]), .I1(n56288), .CO(n43112));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_21 (.CI(n43706), 
            .I0(n2215), .I1(VCC_net), .CO(n43707));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_20_lut (.I0(GND_net), 
            .I1(n2216), .I2(VCC_net), .I3(n43705), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_20 (.CI(n43705), 
            .I0(n2216), .I1(VCC_net), .CO(n43706));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_19_lut (.I0(GND_net), 
            .I1(n2217), .I2(VCC_net), .I3(n43704), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_19 (.CI(n43704), 
            .I0(n2217), .I1(VCC_net), .CO(n43705));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_4 (.CI(n43520), 
            .I0(n932), .I1(GND_net), .CO(n43521));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_3_lut (.I0(GND_net), 
            .I1(n933), .I2(VCC_net), .I3(n43519), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_3 (.CI(n43519), 
            .I0(n933), .I1(VCC_net), .CO(n43520));
    SB_LUT4 add_261_9_lut (.I0(current[7]), .I1(duty[10]), .I2(n56288), 
            .I3(n43110), .O(n263)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_9_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_632_2_lut (.I0(GND_net), 
            .I1(n520), .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i840_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_632_2 (.CI(VCC_net), 
            .I0(n520), .I1(GND_net), .CO(n43519));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1043_3_lut (.I0(n1528), 
            .I1(n1595), .I2(n1554_adj_5610), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_276_i2_3_lut (.I0(encoder0_position_scaled[1]), .I1(motor_state_23__N_123[1]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1807 (.I0(n1728), .I1(n1727), .I2(GND_net), .I3(GND_net), 
            .O(n51360));
    defparam i1_2_lut_adj_1807.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1845_3_lut (.I0(n2714), 
            .I1(n2781), .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_18_lut (.I0(GND_net), 
            .I1(n2218), .I2(VCC_net), .I3(n43703), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15863_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n24373), .I3(GND_net), .O(n29939));   // verilog/coms.v(128[12] 303[6])
    defparam i15863_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_18 (.CI(n43703), 
            .I0(n2218), .I1(VCC_net), .CO(n43704));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_17_lut (.I0(GND_net), 
            .I1(n2219), .I2(VCC_net), .I3(n43702), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_8_lut (.I0(n861), 
            .I1(n828), .I2(VCC_net), .I3(n43518), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_17 (.CI(n43702), 
            .I0(n2219), .I1(VCC_net), .CO(n43703));
    SB_LUT4 n10832_bdd_4_lut_40715 (.I0(n10832), .I1(n419), .I2(current[15]), 
            .I3(duty[23]), .O(n56548));
    defparam n10832_bdd_4_lut_40715.LUT_INIT = 16'he4aa;
    SB_LUT4 n56548_bdd_4_lut (.I0(n56548), .I1(duty[22]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[22]));
    defparam n56548_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40710 (.I0(n10832), .I1(n420), .I2(current[15]), 
            .I3(duty[23]), .O(n56542));
    defparam n10832_bdd_4_lut_40710.LUT_INIT = 16'he4aa;
    SB_LUT4 n56542_bdd_4_lut (.I0(n56542), .I1(duty[21]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[21]));
    defparam n56542_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40705 (.I0(n10832), .I1(n421), .I2(current[15]), 
            .I3(duty[23]), .O(n56536));
    defparam n10832_bdd_4_lut_40705.LUT_INIT = 16'he4aa;
    SB_LUT4 n56536_bdd_4_lut (.I0(n56536), .I1(duty[20]), .I2(n250), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[20]));
    defparam n56536_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1041_3_lut (.I0(n1526), 
            .I1(n1593), .I2(n1554_adj_5610), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1108_3_lut (.I0(n1625), 
            .I1(n1692), .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40700 (.I0(n10832), .I1(n422), .I2(current[15]), 
            .I3(duty[23]), .O(n56524));
    defparam n10832_bdd_4_lut_40700.LUT_INIT = 16'he4aa;
    SB_LUT4 n56524_bdd_4_lut (.I0(n56524), .I1(duty[19]), .I2(n251), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[19]));
    defparam n56524_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1175_3_lut (.I0(n1724), 
            .I1(n1791), .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40690 (.I0(n10832), .I1(n423), .I2(current[15]), 
            .I3(duty[23]), .O(n56518));
    defparam n10832_bdd_4_lut_40690.LUT_INIT = 16'he4aa;
    SB_LUT4 n56518_bdd_4_lut (.I0(n56518), .I1(duty[18]), .I2(n252), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[18]));
    defparam n56518_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1242_3_lut (.I0(n1823), 
            .I1(n1890), .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1309_3_lut (.I0(n1922), 
            .I1(n1989), .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40685 (.I0(n10832), .I1(n424), .I2(current[15]), 
            .I3(duty[23]), .O(n56506));
    defparam n10832_bdd_4_lut_40685.LUT_INIT = 16'he4aa;
    SB_LUT4 n56506_bdd_4_lut (.I0(n56506), .I1(duty[17]), .I2(n253), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[17]));
    defparam n56506_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1376_3_lut (.I0(n2021), 
            .I1(n2088), .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_16_lut (.I0(GND_net), 
            .I1(n2220), .I2(VCC_net), .I3(n43701), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22588_3_lut (.I0(n528), .I1(n1732), .I2(n1733), .I3(GND_net), 
            .O(n36658));
    defparam i22588_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15864_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n24373), .I3(GND_net), .O(n29940));   // verilog/coms.v(128[12] 303[6])
    defparam i15864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1443_3_lut (.I0(n2120), 
            .I1(n2187), .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_16 (.CI(n43701), 
            .I0(n2220), .I1(VCC_net), .CO(n43702));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_15_lut (.I0(GND_net), 
            .I1(n2221), .I2(VCC_net), .I3(n43700), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_7_lut (.I0(GND_net), 
            .I1(n829), .I2(GND_net), .I3(n43517), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1844_3_lut (.I0(n2713), 
            .I1(n2780), .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n1724), .I1(n1725), .I2(n51360), .I3(n1726), 
            .O(n51366));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_7 (.CI(n43517), 
            .I0(n829), .I1(GND_net), .CO(n43518));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1843_3_lut (.I0(n2712), 
            .I1(n2779), .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15865_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n24373), .I3(GND_net), .O(n29941));   // verilog/coms.v(128[12] 303[6])
    defparam i15865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_281_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[2]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15866_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n24373), .I3(GND_net), .O(n29942));   // verilog/coms.v(128[12] 303[6])
    defparam i15866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15867_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n24373), .I3(GND_net), .O(n29943));   // verilog/coms.v(128[12] 303[6])
    defparam i15867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1857_3_lut (.I0(n2726), 
            .I1(n2793), .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1809 (.I0(n1729), .I1(n36658), .I2(n1730), .I3(n1731), 
            .O(n49704));
    defparam i1_4_lut_adj_1809.LUT_INIT = 16'ha080;
    SB_LUT4 i15868_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n24373), .I3(GND_net), .O(n29944));   // verilog/coms.v(128[12] 303[6])
    defparam i15868_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_15 (.CI(n43700), 
            .I0(n2221), .I1(VCC_net), .CO(n43701));
    SB_LUT4 i15869_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n24373), .I3(GND_net), .O(n29945));   // verilog/coms.v(128[12] 303[6])
    defparam i15869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_276_i3_3_lut (.I0(encoder0_position_scaled[2]), .I1(motor_state_23__N_123[2]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_6_lut (.I0(GND_net), 
            .I1(n830), .I2(GND_net), .I3(n43516), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1810 (.I0(n1722), .I1(n1723), .I2(n49704), .I3(n51366), 
            .O(n51372));
    defparam i1_4_lut_adj_1810.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1860_3_lut (.I0(n2729), 
            .I1(n2796), .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1854_3_lut (.I0(n2723), 
            .I1(n2790), .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15870_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position_scaled[7]), 
            .I2(n24373), .I3(GND_net), .O(n29946));   // verilog/coms.v(128[12] 303[6])
    defparam i15870_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_6 (.CI(n43516), 
            .I0(n830), .I1(GND_net), .CO(n43517));
    SB_LUT4 add_263_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n43089), .O(encoder1_position_scaled_23__N_75[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_9 (.CI(n43110), .I0(duty[10]), .I1(n56288), .CO(n43111));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_14_lut (.I0(GND_net), 
            .I1(n2222), .I2(VCC_net), .I3(n43699), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15871_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position_scaled[6]), 
            .I2(n24373), .I3(GND_net), .O(n29947));   // verilog/coms.v(128[12] 303[6])
    defparam i15871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position_scaled_23__N_327[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5620));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_14 (.CI(n43699), 
            .I0(n2222), .I1(VCC_net), .CO(n43700));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_13_lut (.I0(GND_net), 
            .I1(n2223), .I2(VCC_net), .I3(n43698), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15350_3_lut (.I0(deadband[14]), .I1(\data_in_frame[15] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29426));   // verilog/coms.v(128[12] 303[6])
    defparam i15350_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i22_3_lut (.I0(encoder0_position_scaled_23__N_327[21]), 
            .I1(n12_adj_5499), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n523));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i845_rep_28_3_lut (.I0(n523), 
            .I1(n1301), .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i845_rep_28_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(pwm_setpoint_23__N_263));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_261_8_lut (.I0(current[6]), .I1(duty[9]), .I2(n56288), 
            .I3(n43109), .O(n264)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_8_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i40307_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n51372), 
            .O(n1752));
    defparam i40307_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY add_261_8 (.CI(n43109), .I0(duty[9]), .I1(n56288), .CO(n43110));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_13 (.CI(n43698), 
            .I0(n2223), .I1(VCC_net), .CO(n43699));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_5_lut (.I0(GND_net), 
            .I1(n831), .I2(VCC_net), .I3(n43515), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15872_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position_scaled[5]), 
            .I2(n24373), .I3(GND_net), .O(n29948));   // verilog/coms.v(128[12] 303[6])
    defparam i15872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_261_7_lut (.I0(current[5]), .I1(duty[8]), .I2(n56288), 
            .I3(n43108), .O(n265)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_7_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1110_3_lut (.I0(n1627), 
            .I1(n1694), .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1811 (.I0(n1825), .I1(n1824), .I2(n1827), .I3(GND_net), 
            .O(n51720));
    defparam i1_3_lut_adj_1811.LUT_INIT = 16'hfefe;
    SB_LUT4 i22586_3_lut (.I0(n529), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n36656));
    defparam i22586_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_12_lut (.I0(GND_net), 
            .I1(n2224), .I2(VCC_net), .I3(n43697), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1812 (.I0(n1823), .I1(n51720), .I2(n1826), .I3(n1828), 
            .O(n51724));
    defparam i1_4_lut_adj_1812.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1510_3_lut (.I0(n2219), 
            .I1(n2286), .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1813 (.I0(n1829), .I1(n36656), .I2(n1830), .I3(n1831), 
            .O(n49744));
    defparam i1_4_lut_adj_1813.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1814 (.I0(n1821), .I1(n49744), .I2(n1822), .I3(n51724), 
            .O(n51730));
    defparam i1_4_lut_adj_1814.LUT_INIT = 16'hfffe;
    SB_LUT4 i40286_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n51730), 
            .O(n1851));
    defparam i40286_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1577_3_lut (.I0(n2318), 
            .I1(n2385), .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15873_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position_scaled[4]), 
            .I2(n24373), .I3(GND_net), .O(n29949));   // verilog/coms.v(128[12] 303[6])
    defparam i15873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1853_3_lut (.I0(n2722), 
            .I1(n2789), .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15874_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position_scaled[3]), 
            .I2(n24373), .I3(GND_net), .O(n29950));   // verilog/coms.v(128[12] 303[6])
    defparam i15874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1852_3_lut (.I0(n2721), 
            .I1(n2788), .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15875_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position_scaled[2]), 
            .I2(n24373), .I3(GND_net), .O(n29951));   // verilog/coms.v(128[12] 303[6])
    defparam i15875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15876_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position_scaled[1]), 
            .I2(n24373), .I3(GND_net), .O(n29952));   // verilog/coms.v(128[12] 303[6])
    defparam i15876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1815 (.I0(n5_adj_5616), .I1(n122), .I2(n4599), 
            .I3(n63_adj_5615), .O(n6_adj_5662));   // verilog/coms.v(128[12] 303[6])
    defparam i1_4_lut_adj_1815.LUT_INIT = 16'heaaa;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1177_rep_21_3_lut (.I0(n1726), 
            .I1(n1793), .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1177_rep_21_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_12 (.CI(n43697), 
            .I0(n2224), .I1(VCC_net), .CO(n43698));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1644_3_lut (.I0(n2417), 
            .I1(n2484), .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_175_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n43163), .O(n1555)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_11_lut (.I0(GND_net), 
            .I1(n2225), .I2(VCC_net), .I3(n43696), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_5 (.CI(n43515), 
            .I0(n831), .I1(VCC_net), .CO(n43516));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_11 (.CI(n43696), 
            .I0(n2225), .I1(VCC_net), .CO(n43697));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_10_lut (.I0(GND_net), 
            .I1(n2226), .I2(VCC_net), .I3(n43695), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_7 (.CI(n43108), .I0(duty[8]), .I1(n56288), .CO(n43109));
    SB_LUT4 i22584_3_lut (.I0(n530), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n36654));
    defparam i22584_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i33746_3_lut (.I0(n5_adj_5506), .I1(n8587), .I2(n49468), .I3(GND_net), 
            .O(n49473));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1816 (.I0(n57092), .I1(n6_adj_5662), .I2(\FRAME_MATCHER.i_31__N_2845 ), 
            .I3(n4452), .O(n8));   // verilog/coms.v(128[12] 303[6])
    defparam i3_4_lut_adj_1816.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(n1925), .I1(n1928), .I2(n1926), .I3(n1927), 
            .O(n51454));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(n122), .I1(n8), .I2(n63), .I3(n5_adj_5458), 
            .O(n56702));   // verilog/coms.v(128[12] 303[6])
    defparam i4_4_lut.LUT_INIT = 16'hefcf;
    SB_LUT4 i1_4_lut_adj_1818 (.I0(n1929), .I1(n36654), .I2(n1930), .I3(n1931), 
            .O(n49729));
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1855_3_lut (.I0(n2724), 
            .I1(n2791), .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15877_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position_scaled[0]), 
            .I2(n24373), .I3(GND_net), .O(n29953));   // verilog/coms.v(128[12] 303[6])
    defparam i15877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_4_lut (.I0(GND_net), 
            .I1(n832), .I2(GND_net), .I3(n43514), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_4 (.CI(n43514), 
            .I0(n832), .I1(GND_net), .CO(n43515));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_3_lut (.I0(GND_net), 
            .I1(n833), .I2(VCC_net), .I3(n43513), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_3 (.CI(n43513), 
            .I0(n833), .I1(VCC_net), .CO(n43514));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_10 (.CI(n43695), 
            .I0(n2226), .I1(VCC_net), .CO(n43696));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_565_2_lut (.I0(GND_net), 
            .I1(n519), .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_9_lut (.I0(GND_net), 
            .I1(n2227), .I2(VCC_net), .I3(n43694), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_6_lut (.I0(current[4]), .I1(duty[7]), .I2(n56288), 
            .I3(n43107), .O(n266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5522));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1819 (.I0(n1922), .I1(n1923), .I2(n1924), .I3(n51454), 
            .O(n51460));
    defparam i1_4_lut_adj_1819.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1858_3_lut (.I0(n2727), 
            .I1(n2794), .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15731_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29807));   // verilog/coms.v(128[12] 303[6])
    defparam i15731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15878_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position_scaled[15]), 
            .I2(n24373), .I3(GND_net), .O(n29954));   // verilog/coms.v(128[12] 303[6])
    defparam i15878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15879_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position_scaled[14]), 
            .I2(n24373), .I3(GND_net), .O(n29955));   // verilog/coms.v(128[12] 303[6])
    defparam i15879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1820 (.I0(n1920), .I1(n1921), .I2(n51460), .I3(n49729), 
            .O(n51466));
    defparam i1_4_lut_adj_1820.LUT_INIT = 16'hfffe;
    SB_LUT4 i15732_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29808));   // verilog/coms.v(128[12] 303[6])
    defparam i15732_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1859_3_lut (.I0(n2728), 
            .I1(n2795), .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15880_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position_scaled[13]), 
            .I2(n24373), .I3(GND_net), .O(n29956));   // verilog/coms.v(128[12] 303[6])
    defparam i15880_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_565_2 (.CI(VCC_net), 
            .I0(n519), .I1(GND_net), .CO(n43513));
    SB_CARRY add_175_10 (.CI(n43163), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n43164));
    SB_CARRY add_263_4 (.CI(n43082), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n43083));
    SB_LUT4 i15881_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position_scaled[12]), 
            .I2(n24373), .I3(GND_net), .O(n29957));   // verilog/coms.v(128[12] 303[6])
    defparam i15881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n43512), 
            .O(n8584)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n43162), .O(n1556)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_9 (.CI(n43162), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n43163));
    SB_LUT4 add_2750_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n43511), 
            .O(n8585)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n43161), .O(n1557)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_9 (.CI(n43694), 
            .I0(n2227), .I1(VCC_net), .CO(n43695));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1863_3_lut (.I0(n2732), 
            .I1(n2799), .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_8 (.CI(n43161), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n43162));
    SB_LUT4 i40265_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n51466), 
            .O(n1950));
    defparam i40265_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1244_3_lut (.I0(n1825), 
            .I1(n1892), .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1821 (.I0(n2024), .I1(n2026), .I2(GND_net), .I3(GND_net), 
            .O(n51740));
    defparam i1_2_lut_adj_1821.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position_scaled_23__N_327[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5619));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2750_6 (.CI(n43511), .I0(n622), .I1(GND_net), .CO(n43512));
    SB_LUT4 i22648_4_lut (.I0(n531), .I1(n2031), .I2(n2032), .I3(n2033), 
            .O(n36718));
    defparam i22648_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 add_175_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n43160), .O(n1558)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2750_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n43510), 
            .O(n8586)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_6 (.CI(n43107), .I0(duty[7]), .I1(n56288), .CO(n43108));
    SB_CARRY add_175_7 (.CI(n43160), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n43161));
    SB_CARRY add_2750_5 (.CI(n43510), .I0(n623), .I1(VCC_net), .CO(n43511));
    SB_LUT4 mux_281_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[3]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1822 (.I0(n2021), .I1(n2027), .I2(n51740), .I3(n2025), 
            .O(n51746));
    defparam i1_4_lut_adj_1822.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_276_i4_3_lut (.I0(encoder0_position_scaled[3]), .I1(motor_state_23__N_123[3]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_2750_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n43509), 
            .O(n8587)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_4 (.CI(n43509), .I0(n516), .I1(GND_net), .CO(n43510));
    SB_CARRY add_263_11 (.CI(n43089), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n43090));
    SB_LUT4 add_263_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n43088), .O(encoder1_position_scaled_23__N_75[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1823 (.I0(n2029), .I1(n51746), .I2(n36718), .I3(n2030), 
            .O(n51748));
    defparam i1_4_lut_adj_1823.LUT_INIT = 16'heccc;
    SB_LUT4 add_175_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n43159), .O(n1559)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_6 (.CI(n43159), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n43160));
    SB_LUT4 add_175_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n43158), .O(n1560)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_5 (.CI(n43158), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n43159));
    SB_LUT4 add_175_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n43157), .O(n1561)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1824 (.I0(n2022), .I1(n2023), .I2(n2028), .I3(GND_net), 
            .O(n51818));
    defparam i1_3_lut_adj_1824.LUT_INIT = 16'hfefe;
    SB_LUT4 i33747_3_lut (.I0(encoder0_position_scaled_23__N_327[28]), .I1(n49473), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_261_5_lut (.I0(current[3]), .I1(duty[6]), .I2(n56288), 
            .I3(n43106), .O(n267)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_2750_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n43508), 
            .O(n8588)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_5 (.CI(n43106), .I0(duty[6]), .I1(n56288), .CO(n43107));
    SB_LUT4 i1_4_lut_adj_1825 (.I0(n51818), .I1(n2019), .I2(n51748), .I3(n2020), 
            .O(n51752));
    defparam i1_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 add_263_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n43081), .O(encoder1_position_scaled_23__N_75[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1862_3_lut (.I0(n2731), 
            .I1(n2798), .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_263_10 (.CI(n43088), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n43089));
    SB_LUT4 add_261_4_lut (.I0(current[2]), .I1(duty[5]), .I2(n56288), 
            .I3(n43105), .O(n268)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mux_281_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[4]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_8_lut (.I0(GND_net), 
            .I1(n2228), .I2(VCC_net), .I3(n43693), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_276_i5_3_lut (.I0(encoder0_position_scaled[4]), .I1(motor_state_23__N_123[4]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i5_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_8 (.CI(n43693), 
            .I0(n2228), .I1(VCC_net), .CO(n43694));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_99[23]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 i15733_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29809));   // verilog/coms.v(128[12] 303[6])
    defparam i15733_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_4 (.CI(n43157), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n43158));
    SB_CARRY add_261_4 (.CI(n43105), .I0(duty[5]), .I1(n56288), .CO(n43106));
    SB_LUT4 LessThan_17_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5576));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5573));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15734_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29810));   // verilog/coms.v(128[12] 303[6])
    defparam i15734_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1861_3_lut (.I0(n2730), 
            .I1(n2797), .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15735_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29811));   // verilog/coms.v(128[12] 303[6])
    defparam i15735_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5603));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38916_4_lut (.I0(n11_adj_5578), .I1(n9_adj_5599), .I2(n7_adj_5601), 
            .I3(n5_adj_5603), .O(n54709));
    defparam i38916_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5600), .I1(current_limit[9]), 
            .I2(n19_adj_5573), .I3(GND_net), .O(n16_adj_5575));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5604));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i39539_3_lut (.I0(n4_adj_5604), .I1(current_limit[5]), .I2(n11_adj_5578), 
            .I3(GND_net), .O(n55332));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39540_3_lut (.I0(n55332), .I1(current_limit[6]), .I2(n13_adj_5577), 
            .I3(GND_net), .O(n55333));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38911_4_lut (.I0(n17_adj_5574), .I1(n15_adj_5576), .I2(n13_adj_5577), 
            .I3(n54709), .O(n54704));
    defparam i38911_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39679_4_lut (.I0(n16_adj_5575), .I1(n6_adj_5602), .I2(n19_adj_5573), 
            .I3(n54702), .O(n55472));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39679_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i38987_3_lut (.I0(n55333), .I1(current_limit[7]), .I2(n15_adj_5576), 
            .I3(GND_net), .O(n54780));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i38987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39763_4_lut (.I0(n54780), .I1(n55472), .I2(n19_adj_5573), 
            .I3(n54704), .O(n55556));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39763_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39764_3_lut (.I0(n55556), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n55557));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39764_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_7_lut (.I0(GND_net), 
            .I1(n2229), .I2(GND_net), .I3(n43692), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_3 (.CI(n43508), .I0(n625), .I1(VCC_net), .CO(n43509));
    SB_LUT4 add_2750_2_lut (.I0(GND_net), .I1(n518), .I2(GND_net), .I3(VCC_net), 
            .O(n8589)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_281_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[5]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i6_3_lut (.I0(encoder0_position_scaled[5]), .I1(motor_state_23__N_123[5]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i6_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_2750_2 (.CI(VCC_net), .I0(n518), .I1(GND_net), .CO(n43508));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39716_3_lut (.I0(n55557), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5572));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i39716_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i40243_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n51752), 
            .O(n2049));
    defparam i40243_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1856_3_lut (.I0(n2725), 
            .I1(n2792), .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15882_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[7]), .I2(n6_adj_5537), 
            .I3(n27287), .O(n29958));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15882_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_7 (.CI(n43692), 
            .I0(n2229), .I1(GND_net), .CO(n43693));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_6_lut (.I0(GND_net), 
            .I1(n2230), .I2(GND_net), .I3(n43691), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_6 (.CI(n43691), 
            .I0(n2230), .I1(GND_net), .CO(n43692));
    SB_LUT4 add_175_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n43156), .O(n1562)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_5_lut (.I0(GND_net), 
            .I1(n2231), .I2(VCC_net), .I3(n43690), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15736_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29812));   // verilog/coms.v(128[12] 303[6])
    defparam i15736_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_175_3 (.CI(n43156), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n43157));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5535), .I3(n43500), .O(displacement_23__N_99[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5534), .I3(n43499), .O(displacement_23__N_99[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n10832_bdd_4_lut_40675 (.I0(n10832), .I1(n425), .I2(current[15]), 
            .I3(duty[23]), .O(n56500));
    defparam n10832_bdd_4_lut_40675.LUT_INIT = 16'he4aa;
    SB_LUT4 n56500_bdd_4_lut (.I0(n56500), .I1(duty[16]), .I2(n254), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[16]));
    defparam n56500_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15883_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[8]), .I2(n5_adj_5538), 
            .I3(n27222), .O(n29959));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15883_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15671_3_lut (.I0(n28795), .I1(\ID_READOUT_FSM.state [0]), .I2(n7974), 
            .I3(GND_net), .O(n29747));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15671_3_lut.LUT_INIT = 16'h4646;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1851_3_lut (.I0(n2720), 
            .I1(n2787), .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_281_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[6]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i7_3_lut (.I0(encoder0_position_scaled[6]), .I1(motor_state_23__N_123[6]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15737_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29813));   // verilog/coms.v(128[12] 303[6])
    defparam i15737_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1865_3_lut (.I0(n538), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5523));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1826 (.I0(n36101), .I1(n49611), .I2(state_adj_5716[0]), 
            .I3(read), .O(n48264));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1826.LUT_INIT = 16'h8280;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_5 (.CI(n43690), 
            .I0(n2231), .I1(VCC_net), .CO(n43691));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_4_lut (.I0(GND_net), 
            .I1(n2232), .I2(GND_net), .I3(n43689), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_99[22]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15738_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29814));   // verilog/coms.v(128[12] 303[6])
    defparam i15738_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1864_3_lut (.I0(n2733), 
            .I1(n2800), .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_4 (.CI(n43689), 
            .I0(n2232), .I1(GND_net), .CO(n43690));
    SB_LUT4 add_175_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1563)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n43499), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5534), .CO(n43500));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_3_lut (.I0(GND_net), 
            .I1(n2233_adj_5612), .I2(VCC_net), .I3(n43688), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_3_lut (.I0(current[1]), .I1(duty[4]), .I2(n56288), 
            .I3(n43104), .O(n269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_3 (.CI(n43688), 
            .I0(n2233_adj_5612), .I1(VCC_net), .CO(n43689));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1503_2_lut (.I0(GND_net), 
            .I1(n533), .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5533), .I3(n43498), .O(displacement_23__N_99[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n43156));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1503_2 (.CI(VCC_net), 
            .I0(n533), .I1(GND_net), .CO(n43688));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_21_lut (.I0(n56010), 
            .I1(n2115), .I2(VCC_net), .I3(n43687), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n43498), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5533), .CO(n43499));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5532), .I3(n43497), .O(displacement_23__N_99[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_20_lut (.I0(GND_net), 
            .I1(n2116), .I2(VCC_net), .I3(n43686), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_20 (.CI(n43686), 
            .I0(n2116), .I1(VCC_net), .CO(n43687));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_19_lut (.I0(GND_net), 
            .I1(n2117), .I2(VCC_net), .I3(n43685), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_19 (.CI(n43685), 
            .I0(n2117), .I1(VCC_net), .CO(n43686));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_18_lut (.I0(GND_net), 
            .I1(n2118), .I2(VCC_net), .I3(n43684), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_18 (.CI(n43684), 
            .I0(n2118), .I1(VCC_net), .CO(n43685));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n43497), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5532), .CO(n43498));
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_99[21]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_99[20]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_99[19]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_99[18]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_99[17]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_99[16]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_99[15]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_99[14]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_99[13]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_99[12]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_99[11]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_99[10]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_99[9]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_99[8]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_99[7]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_99[6]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_99[5]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_99[4]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_99[3]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_99[2]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_99[1]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[23]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[22]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[21]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[20]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[19]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[18]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[17]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[16]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[15]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[14]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[13]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[12]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[11]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_75[10]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[9]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[8]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[7]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[6]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[5]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[4]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[3]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[2]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_75[1]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[23]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 mux_281_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[7]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i8_3_lut (.I0(encoder0_position_scaled[7]), .I1(motor_state_23__N_123[7]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i6_3_lut (.I0(encoder0_position_scaled_23__N_327[5]), 
            .I1(n28), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n539));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15659_3_lut (.I0(n29186), .I1(r_Bit_Index[0]), .I2(n28762), 
            .I3(GND_net), .O(n29735));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15659_3_lut.LUT_INIT = 16'h1414;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[22]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 mux_281_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[8]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[21]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[20]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[19]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[18]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[17]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[16]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[15]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[14]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[13]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[12]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[11]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_51[10]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[9]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[8]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[7]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[6]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[5]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[4]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[3]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[2]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_51[1]));   // verilog/TinyFPGA_B.v(321[10] 334[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_17_lut (.I0(GND_net), 
            .I1(n2119), .I2(VCC_net), .I3(n43683), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5531), .I3(n43496), .O(displacement_23__N_99[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_276_i9_3_lut (.I0(encoder0_position_scaled[8]), .I1(motor_state_23__N_123[8]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i22566_3_lut (.I0(n539), .I1(n2832), .I2(n2833), .I3(GND_net), 
            .O(n36636));
    defparam i22566_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(n2827), .I1(n2826), .I2(n2823), .I3(n2820), 
            .O(n51832));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1828 (.I0(n2821), .I1(n2822), .I2(n2828), .I3(n2825), 
            .O(n51834));
    defparam i1_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 i15656_3_lut (.I0(n29184), .I1(r_Bit_Index_adj_5736[0]), .I2(n28758), 
            .I3(GND_net), .O(n29732));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15656_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i1_4_lut_adj_1829 (.I0(n51834), .I1(n51832), .I2(n2819), .I3(n2824), 
            .O(n51838));
    defparam i1_4_lut_adj_1829.LUT_INIT = 16'hfffe;
    SB_LUT4 i15889_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[9]), .I2(n5_adj_5570), 
            .I3(n27222), .O(n29965));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15889_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1311_3_lut (.I0(n1924), 
            .I1(n1991), .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1830 (.I0(n2829), .I1(n36636), .I2(n2830), .I3(n2831), 
            .O(n49816));
    defparam i1_4_lut_adj_1830.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5524));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1831 (.I0(n2816), .I1(n2817), .I2(n51838), .I3(n2818), 
            .O(n51844));
    defparam i1_4_lut_adj_1831.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1832 (.I0(n2814), .I1(n2815), .I2(n51844), .I3(n49816), 
            .O(n51850));
    defparam i1_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_281_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[9]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i10_3_lut (.I0(encoder0_position_scaled[9]), .I1(motor_state_23__N_123[9]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1833 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n51850), 
            .O(n51856));
    defparam i1_4_lut_adj_1833.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_17 (.CI(n43683), 
            .I0(n2119), .I1(VCC_net), .CO(n43684));
    SB_LUT4 i40030_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n51856), 
            .O(n2841));
    defparam i40030_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1834 (.I0(current_limit[13]), .I1(n24_adj_5572), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n50462));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1834.LUT_INIT = 16'hfffe;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n43496), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5531), .CO(n43497));
    SB_LUT4 mux_281_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[10]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1775_3_lut (.I0(n2612), 
            .I1(n2679), .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_276_i11_3_lut (.I0(encoder0_position_scaled[10]), .I1(motor_state_23__N_123[10]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5530), .I3(n43495), .O(displacement_23__N_99[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n43495), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5530), .CO(n43496));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1774_3_lut (.I0(n2611), 
            .I1(n2678), .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1777_3_lut (.I0(n2614), 
            .I1(n2681), .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1776_3_lut (.I0(n2613), 
            .I1(n2680), .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40057_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55850));
    defparam i40057_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_281_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[11]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1835 (.I0(n2724), .I1(n2727), .I2(n2723), .I3(n2728), 
            .O(n51420));
    defparam i1_4_lut_adj_1835.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5525));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1836 (.I0(n2721), .I1(n2725), .I2(n2726), .I3(n2722), 
            .O(n51422));
    defparam i1_4_lut_adj_1836.LUT_INIT = 16'hfffe;
    SB_LUT4 i22634_4_lut (.I0(n538), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n36704));
    defparam i22634_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 mux_276_i12_3_lut (.I0(encoder0_position_scaled[11]), .I1(motor_state_23__N_123[11]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_281_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[12]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1837 (.I0(n2719), .I1(n2720), .I2(n51422), .I3(n51420), 
            .O(n51428));
    defparam i1_4_lut_adj_1837.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5526));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5527));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_276_i13_3_lut (.I0(encoder0_position_scaled[12]), .I1(motor_state_23__N_123[12]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_3_lut_adj_1838 (.I0(n52823), .I1(n2124), .I2(n2127), .I3(GND_net), 
            .O(n51560));
    defparam i1_3_lut_adj_1838.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1839 (.I0(n2729), .I1(n2730), .I2(GND_net), .I3(GND_net), 
            .O(n51940));
    defparam i1_2_lut_adj_1839.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5529), .I3(n43494), .O(displacement_23__N_99[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n43494), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5529), .CO(n43495));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5528), .I3(n43493), .O(displacement_23__N_99[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n43493), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5528), .CO(n43494));
    SB_LUT4 mux_281_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[13]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5527), .I3(n43492), .O(displacement_23__N_99[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_276_i14_3_lut (.I0(encoder0_position_scaled[13]), .I1(motor_state_23__N_123[13]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1840 (.I0(n2718), .I1(n51940), .I2(n51428), .I3(n36704), 
            .O(n51432));
    defparam i1_4_lut_adj_1840.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1841 (.I0(n2715), .I1(n2716), .I2(n2717), .I3(n51432), 
            .O(n51438));
    defparam i1_4_lut_adj_1841.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n43492), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5527), .CO(n43493));
    SB_LUT4 i1_4_lut_adj_1842 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n51438), 
            .O(n51444));
    defparam i1_4_lut_adj_1842.LUT_INIT = 16'hfffe;
    SB_LUT4 i40060_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n51444), 
            .O(n2742));
    defparam i40060_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5526), .I3(n43491), .O(displacement_23__N_99[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5528));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5529));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40086_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55879));
    defparam i40086_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15890_4_lut (.I0(CS_MISO_c), .I1(data_adj_5722[10]), .I2(n5), 
            .I3(n27222), .O(n29966));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15890_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_16_lut (.I0(GND_net), 
            .I1(n2120), .I2(VCC_net), .I3(n43682), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5530));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n43491), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5526), .CO(n43492));
    SB_LUT4 mux_281_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[14]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i15_3_lut (.I0(encoder0_position_scaled[14]), .I1(motor_state_23__N_123[14]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5525), .I3(n43490), .O(displacement_23__N_99[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n43490), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5525), .CO(n43491));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5524), .I3(n43489), .O(displacement_23__N_99[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n43489), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5524), .CO(n43490));
    SB_LUT4 i1_4_lut_adj_1843 (.I0(current_limit[13]), .I1(n24_adj_5572), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n50464));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1843.LUT_INIT = 16'h8000;
    SB_LUT4 mux_281_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[15]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i16_3_lut (.I0(encoder0_position_scaled[15]), .I1(motor_state_23__N_123[15]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1844 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n50464), .I3(n50462), .O(n296));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1844.LUT_INIT = 16'hb3a2;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5523), .I3(n43488), .O(displacement_23__N_99[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
           .D(n29747));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n43488), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5523), .CO(n43489));
    SB_LUT4 mux_281_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[16]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5522), .I3(n43487), .O(displacement_23__N_99[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_3 (.CI(n43104), .I0(duty[4]), .I1(n56288), .CO(n43105));
    SB_LUT4 mux_276_i17_3_lut (.I0(encoder0_position_scaled[16]), .I1(motor_state_23__N_123[16]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder1_position_scaled_23__I_4_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_359));   // verilog/TinyFPGA_B.v(323[33:52])
    defparam encoder1_position_scaled_23__I_4_4_lut.LUT_INIT = 16'hccc8;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n43487), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5522), .CO(n43488));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5521), .I3(n43486), .O(displacement_23__N_99[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n43486), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5521), .CO(n43487));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5520), .I3(n43485), .O(displacement_23__N_99[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n43485), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5520), .CO(n43486));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_16 (.CI(n43682), 
            .I0(n2120), .I1(VCC_net), .CO(n43683));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_15_lut (.I0(GND_net), 
            .I1(n2121), .I2(VCC_net), .I3(n43681), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5519), .I3(n43484), .O(displacement_23__N_99[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_15 (.CI(n43681), 
            .I0(n2121), .I1(VCC_net), .CO(n43682));
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n7593), 
            .D(n1563), .R(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[23]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[22]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF dti_counter_2279__i0 (.Q(dti_counter[0]), .C(clk16MHz), .D(n55));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n43484), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5519), .CO(n43485));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5518), .I3(n43483), .O(displacement_23__N_99[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n43483), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5518), .CO(n43484));
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[21]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[20]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5517), .I3(n43482), .O(displacement_23__N_99[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n43482), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5517), .CO(n43483));
    SB_LUT4 i40142_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55935));
    defparam i40142_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_14_lut (.I0(GND_net), 
            .I1(n2122), .I2(VCC_net), .I3(n43680), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_14 (.CI(n43680), 
            .I0(n2122), .I1(VCC_net), .CO(n43681));
    SB_LUT4 i40193_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n55986));
    defparam i40193_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[19]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[18]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[17]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[16]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[15]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[14]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[13]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[12]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[11]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[10]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[9]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[8]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[7]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[6]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[5]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[4]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 i22580_3_lut (.I0(n532), .I1(n2132), .I2(n2133), .I3(GND_net), 
            .O(n36650));
    defparam i22580_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[3]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1845 (.I0(n2123), .I1(n51560), .I2(n2128), .I3(n2126), 
            .O(n51564));
    defparam i1_4_lut_adj_1845.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[2]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1846 (.I0(n2129), .I1(n36650), .I2(n2130), .I3(n2131), 
            .O(n49746));
    defparam i1_4_lut_adj_1846.LUT_INIT = 16'ha080;
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[1]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1847 (.I0(n2121), .I1(n49746), .I2(n2122), .I3(n51564), 
            .O(n51570));
    defparam i1_4_lut_adj_1847.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1848 (.I0(n2118), .I1(n2119), .I2(n2120), .I3(n51570), 
            .O(n51576));
    defparam i1_4_lut_adj_1848.LUT_INIT = 16'hfffe;
    SB_LUT4 i40220_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n51576), 
            .O(n2148));
    defparam i40220_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1378_3_lut (.I0(n2023), 
            .I1(n2090), .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22578_3_lut (.I0(n533), .I1(n2232), .I2(n2233_adj_5612), 
            .I3(GND_net), .O(n36648));
    defparam i22578_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1849 (.I0(n2223), .I1(n2227), .I2(n2224), .I3(n2225), 
            .O(n51766));
    defparam i1_4_lut_adj_1849.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1850 (.I0(n2226), .I1(n51766), .I2(n2222), .I3(n2228), 
            .O(n51768));
    defparam i1_4_lut_adj_1850.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1851 (.I0(n2229), .I1(n36648), .I2(n2230), .I3(n2231), 
            .O(n49772));
    defparam i1_4_lut_adj_1851.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1852 (.I0(n2219), .I1(n2220), .I2(n2221), .I3(n51768), 
            .O(n51774));
    defparam i1_4_lut_adj_1852.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1853 (.I0(n2217), .I1(n2218), .I2(n51774), .I3(n49772), 
            .O(n51780));
    defparam i1_4_lut_adj_1853.LUT_INIT = 16'hfffe;
    SB_LUT4 i40196_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n51780), 
            .O(n2247));
    defparam i40196_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1445_3_lut (.I0(n2122), 
            .I1(n2189), .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1854 (.I0(n2321), .I1(n2322), .I2(n2324), .I3(GND_net), 
            .O(n51380));
    defparam i1_3_lut_adj_1854.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1855 (.I0(n2326), .I1(n2325), .I2(GND_net), .I3(GND_net), 
            .O(n51646));
    defparam i1_2_lut_adj_1855.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1039_3_lut (.I0(n1524), 
            .I1(n1591), .I2(n1554_adj_5610), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22642_4_lut (.I0(n534), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n36712));
    defparam i22642_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1856 (.I0(n2328), .I1(n51646), .I2(n2323), .I3(n2327), 
            .O(n51652));
    defparam i1_4_lut_adj_1856.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1857 (.I0(n2329), .I1(n51652), .I2(n36712), .I3(n2330), 
            .O(n51654));
    defparam i1_4_lut_adj_1857.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1106_3_lut (.I0(n1623), 
            .I1(n1690), .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1858 (.I0(n2316), .I1(n2318), .I2(n2320), .I3(n51380), 
            .O(n51386));
    defparam i1_4_lut_adj_1858.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1859 (.I0(n2317), .I1(n2315), .I2(n2319), .I3(n51654), 
            .O(n51089));
    defparam i1_4_lut_adj_1859.LUT_INIT = 16'hfffe;
    SB_LUT4 i40171_4_lut (.I0(n2314), .I1(n2313), .I2(n51089), .I3(n51386), 
            .O(n2346));
    defparam i40171_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1173_3_lut (.I0(n1722), 
            .I1(n1789), .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1512_3_lut (.I0(n2221), 
            .I1(n2288), .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40670 (.I0(n10832), .I1(n426), .I2(current[15]), 
            .I3(duty[23]), .O(n56458));
    defparam n10832_bdd_4_lut_40670.LUT_INIT = 16'he4aa;
    SB_LUT4 n56458_bdd_4_lut (.I0(n56458), .I1(duty[15]), .I2(n255), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[15]));
    defparam n56458_bdd_4_lut.LUT_INIT = 16'haad8;
    GND i1 (.Y(GND_net));
    SB_LUT4 mux_281_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[17]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i18_3_lut (.I0(encoder0_position_scaled[17]), .I1(motor_state_23__N_123[17]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1240_3_lut (.I0(n1821), 
            .I1(n1888), .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHC_214 (.Q(GHC), .C(clk16MHz), .E(n28583), .D(GHC_N_514), 
            .R(n29049));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i1_4_lut_adj_1860 (.I0(n2423), .I1(n2424), .I2(n2425), .I3(n2428), 
            .O(n51802));
    defparam i1_4_lut_adj_1860.LUT_INIT = 16'hfffe;
    SB_LUT4 i21950_2_lut (.I0(duty[15]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4914));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21950_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1307_3_lut (.I0(n1920), 
            .I1(n1987), .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5531));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n10832_bdd_4_lut_40636 (.I0(n10832), .I1(n427), .I2(current[15]), 
            .I3(duty[23]), .O(n56452));
    defparam n10832_bdd_4_lut_40636.LUT_INIT = 16'he4aa;
    SB_LUT4 n56452_bdd_4_lut (.I0(n56452), .I1(duty[14]), .I2(n256), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[14]));
    defparam n56452_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1374_3_lut (.I0(n2019), 
            .I1(n2086), .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40631 (.I0(n10832), .I1(n428), .I2(current[15]), 
            .I3(duty[23]), .O(n56446));
    defparam n10832_bdd_4_lut_40631.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_281_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[18]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n56446_bdd_4_lut (.I0(n56446), .I1(duty[13]), .I2(n257), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[13]));
    defparam n56446_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1441_3_lut (.I0(n2118), 
            .I1(n2185), .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40626 (.I0(n10832), .I1(n429), .I2(current[15]), 
            .I3(duty[23]), .O(n56440));
    defparam n10832_bdd_4_lut_40626.LUT_INIT = 16'he4aa;
    SB_LUT4 n56440_bdd_4_lut (.I0(n56440), .I1(duty[12]), .I2(n258), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[12]));
    defparam n56440_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_13_lut (.I0(GND_net), 
            .I1(n2123), .I2(VCC_net), .I3(n43679), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1508_3_lut (.I0(n2217), 
            .I1(n2284), .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_13 (.CI(n43679), 
            .I0(n2123), .I1(VCC_net), .CO(n43680));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5516), .I3(n43481), .O(displacement_23__N_99[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1575_3_lut (.I0(n2316), 
            .I1(n2383), .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1642_3_lut (.I0(n2415), 
            .I1(n2482), .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_12_lut (.I0(GND_net), 
            .I1(n2124), .I2(VCC_net), .I3(n43678), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1643_3_lut (.I0(n2416), 
            .I1(n2483), .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n43481), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5516), .CO(n43482));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1711_3_lut (.I0(n2516), 
            .I1(n2583), .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_276_i19_3_lut (.I0(encoder0_position_scaled[18]), .I1(motor_state_23__N_123[18]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 n10832_bdd_4_lut_40621 (.I0(n10832), .I1(n430), .I2(current[11]), 
            .I3(duty[23]), .O(n56410));
    defparam n10832_bdd_4_lut_40621.LUT_INIT = 16'he4aa;
    SB_LUT4 n56410_bdd_4_lut (.I0(n56410), .I1(duty[11]), .I2(n259), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[11]));
    defparam n56410_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1710_3_lut (.I0(n2515), 
            .I1(n2582), .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40596 (.I0(n10832), .I1(n431), .I2(current[10]), 
            .I3(duty[23]), .O(n56404));
    defparam n10832_bdd_4_lut_40596.LUT_INIT = 16'he4aa;
    SB_LUT4 n56404_bdd_4_lut (.I0(n56404), .I1(duty[10]), .I2(n260), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[10]));
    defparam n56404_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1709_3_lut (.I0(n2514), 
            .I1(n2581), .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22678_4_lut (.I0(n519), .I1(n831), .I2(n832), .I3(n833), 
            .O(n36748));
    defparam i22678_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 n10832_bdd_4_lut_40591 (.I0(n10832), .I1(n432), .I2(current[9]), 
            .I3(duty[23]), .O(n56392));
    defparam n10832_bdd_4_lut_40591.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_281_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[19]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i20_3_lut (.I0(encoder0_position_scaled[19]), .I1(motor_state_23__N_123[19]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i40217_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56010));
    defparam i40217_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40240_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56033));
    defparam i40240_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_281_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[20]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i21_3_lut (.I0(encoder0_position_scaled[20]), .I1(motor_state_23__N_123[20]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i21_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_12 (.CI(n43678), 
            .I0(n2124), .I1(VCC_net), .CO(n43679));
    SB_LUT4 i15245_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n24373), .I3(GND_net), .O(n29321));   // verilog/coms.v(128[12] 303[6])
    defparam i15245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_281_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15), .I3(n15_adj_5485), .O(motor_state_23__N_123[21]));   // verilog/TinyFPGA_B.v(284[5] 286[10])
    defparam mux_281_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_276_i22_3_lut (.I0(encoder0_position_scaled[21]), .I1(motor_state_23__N_123[21]), 
            .I2(n15_adj_5457), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(283[5] 286[10])
    defparam mux_276_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1861 (.I0(n2420), .I1(n51802), .I2(n2426), .I3(n2427), 
            .O(n51806));
    defparam i1_4_lut_adj_1861.LUT_INIT = 16'hfffe;
    SB_LUT4 i40262_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56055));
    defparam i40262_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5532));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_11_lut (.I0(GND_net), 
            .I1(n52823), .I2(VCC_net), .I3(n43677), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5515), .I3(n43480), .O(displacement_23__N_99[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n43480), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5515), .CO(n43481));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i26_3_lut (.I0(encoder0_position_scaled_23__N_327[25]), 
            .I1(n8_adj_5503), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i573_rep_32_3_lut (.I0(n519), 
            .I1(n901), .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i573_rep_32_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR GHB_212 (.Q(GHB), .C(clk16MHz), .E(n28583), .D(GHB_N_500), 
            .R(n29049));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_11 (.CI(n43677), 
            .I0(n52823), .I1(VCC_net), .CO(n43678));
    SB_LUT4 i15182_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n49594), .I3(GND_net), .O(n29258));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_10_lut (.I0(GND_net), 
            .I1(n2126), .I2(VCC_net), .I3(n43676), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5533));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_10 (.CI(n43676), 
            .I0(n2126), .I1(VCC_net), .CO(n43677));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5514), .I3(n43479), .O(displacement_23__N_99[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n43479), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5514), .CO(n43480));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_9_lut (.I0(GND_net), 
            .I1(n2127), .I2(VCC_net), .I3(n43675), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_9 (.CI(n43675), 
            .I0(n2127), .I1(VCC_net), .CO(n43676));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5513), .I3(n43478), .O(displacement_23__N_99[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n43478), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5513), .CO(n43479));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_8_lut (.I0(GND_net), 
            .I1(n2128), .I2(VCC_net), .I3(n43674), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_2_lut (.I0(GND_net), .I1(duty[3]), .I2(n211), .I3(GND_net), 
            .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_261_2 (.CI(GND_net), .I0(duty[3]), .I1(n211), .CO(n43104));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5512), .I3(VCC_net), .O(displacement_23__N_99[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1862 (.I0(n2418), .I1(n2416), .I2(n2419), .I3(n2422), 
            .O(n50765));
    defparam i1_4_lut_adj_1862.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5534));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5535));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_8 (.CI(n43674), 
            .I0(n2128), .I1(VCC_net), .CO(n43675));
    SB_LUT4 n56392_bdd_4_lut (.I0(n56392), .I1(duty[9]), .I2(n261), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[9]));
    defparam n56392_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i22742_4_lut (.I0(n829), .I1(n828), .I2(n36748), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i22742_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i33744_3_lut (.I0(n4_adj_5507), .I1(n8586), .I2(n49468), .I3(GND_net), 
            .O(n49471));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33745_3_lut (.I0(encoder0_position_scaled_23__N_327[29]), .I1(n49471), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5512), .CO(n43478));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_7_lut (.I0(GND_net), 
            .I1(n2129), .I2(GND_net), .I3(n43673), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n10832_bdd_4_lut_40581 (.I0(n10832), .I1(n433), .I2(current[8]), 
            .I3(duty[23]), .O(n56362));
    defparam n10832_bdd_4_lut_40581.LUT_INIT = 16'he4aa;
    SB_LUT4 n56362_bdd_4_lut (.I0(n56362), .I1(duty[8]), .I2(n262), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[8]));
    defparam n56362_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40558 (.I0(n10832), .I1(n434), .I2(current[7]), 
            .I3(duty[23]), .O(n56356));
    defparam n10832_bdd_4_lut_40558.LUT_INIT = 16'he4aa;
    SB_LUT4 n56356_bdd_4_lut (.I0(n56356), .I1(duty[7]), .I2(n263), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[7]));
    defparam n56356_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i770_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_7 (.CI(n43673), 
            .I0(n2129), .I1(GND_net), .CO(n43674));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_6_lut (.I0(GND_net), 
            .I1(n2130), .I2(GND_net), .I3(n43672), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n10832_bdd_4_lut_40553 (.I0(n10832), .I1(n435), .I2(current[6]), 
            .I3(duty[23]), .O(n56350));
    defparam n10832_bdd_4_lut_40553.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_6 (.CI(n43672), 
            .I0(n2130), .I1(GND_net), .CO(n43673));
    SB_LUT4 n56350_bdd_4_lut (.I0(n56350), .I1(duty[6]), .I2(n264), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[6]));
    defparam n56350_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR GHA_210 (.Q(GHA), .C(clk16MHz), .E(n28583), .D(GHA_N_478), 
            .R(n29049));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i28_3_lut (.I0(encoder0_position_scaled_23__N_327[27]), 
            .I1(n6_adj_5505), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n625));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_5_lut (.I0(GND_net), 
            .I1(n2131), .I2(VCC_net), .I3(n43671), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_5 (.CI(n43671), 
            .I0(n2131), .I1(VCC_net), .CO(n43672));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i29_3_lut (.I0(encoder0_position_scaled_23__N_327[28]), 
            .I1(n5_adj_5506), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_263_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n43103), .O(encoder1_position_scaled_23__N_75[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_4_lut (.I0(GND_net), 
            .I1(n2132), .I2(GND_net), .I3(n43670), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i30_3_lut (.I0(encoder0_position_scaled_23__N_327[29]), 
            .I1(n4_adj_5507), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n623));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_4 (.CI(n43670), 
            .I0(n2132), .I1(GND_net), .CO(n43671));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_3_lut (.I0(GND_net), 
            .I1(n2133), .I2(VCC_net), .I3(n43669), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_3 (.CI(n43669), 
            .I0(n2133), .I1(VCC_net), .CO(n43670));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1436_2_lut (.I0(GND_net), 
            .I1(n532), .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1436_2 (.CI(VCC_net), 
            .I0(n532), .I1(GND_net), .CO(n43669));
    SB_LUT4 add_263_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n43102), .O(encoder1_position_scaled_23__N_75[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_20_lut (.I0(n56033), 
            .I1(n2016), .I2(VCC_net), .I3(n43668), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_19_lut (.I0(GND_net), 
            .I1(n2017), .I2(VCC_net), .I3(n43667), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_19 (.CI(n43667), 
            .I0(n2017), .I1(VCC_net), .CO(n43668));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i31_3_lut (.I0(encoder0_position_scaled_23__N_327[30]), 
            .I1(n3_adj_5508), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n622));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_18_lut (.I0(GND_net), 
            .I1(n2018), .I2(VCC_net), .I3(n43666), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33751_3_lut (.I0(encoder0_position_scaled_23__N_327[26]), .I1(n49477), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33751_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_18 (.CI(n43666), 
            .I0(n2018), .I1(VCC_net), .CO(n43667));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_17_lut (.I0(GND_net), 
            .I1(n2019), .I2(VCC_net), .I3(n43665), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_17 (.CI(n43665), 
            .I0(n2019), .I1(VCC_net), .CO(n43666));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_16_lut (.I0(GND_net), 
            .I1(n2020), .I2(VCC_net), .I3(n43664), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_16 (.CI(n43664), 
            .I0(n2020), .I1(VCC_net), .CO(n43665));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_15_lut (.I0(GND_net), 
            .I1(n2021), .I2(VCC_net), .I3(n43663), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_15 (.CI(n43663), 
            .I0(n2021), .I1(VCC_net), .CO(n43664));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_14_lut (.I0(GND_net), 
            .I1(n2022), .I2(VCC_net), .I3(n43662), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_14 (.CI(n43662), 
            .I0(n2022), .I1(VCC_net), .CO(n43663));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_13_lut (.I0(GND_net), 
            .I1(n2023), .I2(VCC_net), .I3(n43661), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_13 (.CI(n43661), 
            .I0(n2023), .I1(VCC_net), .CO(n43662));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_12_lut (.I0(GND_net), 
            .I1(n2024), .I2(VCC_net), .I3(n43660), .O(n2091_adj_5611)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_12 (.CI(n43660), 
            .I0(n2024), .I1(VCC_net), .CO(n43661));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_11_lut (.I0(GND_net), 
            .I1(n2025), .I2(VCC_net), .I3(n43659), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n43468), .O(n330)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n43467), .O(n334)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1863 (.I0(control_mode[0]), .I1(n27284), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_5485));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i1_2_lut_3_lut_adj_1863.LUT_INIT = 16'hefef;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n6_adj_5668), .D(commutation_state_7__N_264[0]), .S(commutation_state_7__N_272));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY add_263_24 (.CI(n43102), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n43103));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_11 (.CI(n43659), 
            .I0(n2025), .I1(VCC_net), .CO(n43660));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i904_rep_27_3_lut (.I0(n1325), 
            .I1(n1392), .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i904_rep_27_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_10_lut (.I0(GND_net), 
            .I1(n2026), .I2(VCC_net), .I3(n43658), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_14 (.CI(n43467), .I0(GND_net), .I1(n2), 
            .CO(n43468));
    SB_LUT4 unary_minus_19_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5466), 
            .I3(n43466), .O(n335)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_10 (.CI(n43658), 
            .I0(n2026), .I1(VCC_net), .CO(n43659));
    SB_CARRY unary_minus_19_add_3_13 (.CI(n43466), .I0(GND_net), .I1(n14_adj_5466), 
            .CO(n43467));
    SB_LUT4 unary_minus_19_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5467), 
            .I3(n43465), .O(n336)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_12 (.CI(n43465), .I0(GND_net), .I1(n15_adj_5467), 
            .CO(n43466));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_9_lut (.I0(GND_net), 
            .I1(n2027), .I2(VCC_net), .I3(n43657), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5468), 
            .I3(n43464), .O(n337)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_9 (.CI(n43657), 
            .I0(n2027), .I1(VCC_net), .CO(n43658));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_8_lut (.I0(GND_net), 
            .I1(n2028), .I2(VCC_net), .I3(n43656), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_8 (.CI(n43656), 
            .I0(n2028), .I1(VCC_net), .CO(n43657));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_7_lut (.I0(GND_net), 
            .I1(n2029), .I2(GND_net), .I3(n43655), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33743_3_lut (.I0(encoder0_position_scaled_23__N_327[30]), .I1(n49469), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15343_3_lut (.I0(deadband[20]), .I1(\data_in_frame[14] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29419));   // verilog/coms.v(128[12] 303[6])
    defparam i15343_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5667));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(delay_counter[28]), .I1(n12_adj_5667), .I2(delay_counter[25]), 
            .I3(delay_counter[30]), .O(n27140));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1864 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n27137));
    defparam i2_3_lut_adj_1864.LUT_INIT = 16'hfefe;
    SB_CARRY unary_minus_19_add_3_11 (.CI(n43464), .I0(GND_net), .I1(n16_adj_5468), 
            .CO(n43465));
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5484));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 unary_minus_19_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5469), 
            .I3(n43463), .O(n338)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1865 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5483));
    defparam i6_4_lut_adj_1865.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5483), .I1(delay_counter[2]), .I2(n14_adj_5484), 
            .I3(delay_counter[6]), .O(n27143));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4658_4_lut (.I0(n27143), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5613));
    defparam i4658_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1866 (.I0(n24_adj_5613), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n51177));
    defparam i2_4_lut_adj_1866.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1867 (.I0(n51177), .I1(delay_counter[18]), .I2(n27137), 
            .I3(GND_net), .O(n50777));
    defparam i2_3_lut_adj_1867.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1868 (.I0(delay_counter[23]), .I1(n50777), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5663));
    defparam i2_4_lut_adj_1868.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut_adj_1869 (.I0(n7_adj_5663), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n27140), .O(n62));
    defparam i4_4_lut_adj_1869.LUT_INIT = 16'hfffe;
    SB_LUT4 i5785_3_lut (.I0(n62), .I1(\ID_READOUT_FSM.state [0]), .I2(delay_counter[31]), 
            .I3(GND_net), .O(n20976));
    defparam i5785_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i1_2_lut_adj_1870 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5664));
    defparam i1_2_lut_adj_1870.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1871 (.I0(delay_counter[9]), .I1(n4_adj_5664), 
            .I2(delay_counter[10]), .I3(n27143), .O(n51094));
    defparam i2_4_lut_adj_1871.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1872 (.I0(n51094), .I1(n27137), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n50786));
    defparam i2_4_lut_adj_1872.LUT_INIT = 16'hffec;
    SB_CARRY unary_minus_19_add_3_10 (.CI(n43463), .I0(GND_net), .I1(n17_adj_5469), 
            .CO(n43464));
    SB_LUT4 unary_minus_19_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5470), 
            .I3(n43462), .O(n339)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5665));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_7 (.CI(n43655), 
            .I0(n2029), .I1(GND_net), .CO(n43656));
    SB_LUT4 i2_4_lut_adj_1873 (.I0(delay_counter[22]), .I1(n50786), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5666));
    defparam i2_4_lut_adj_1873.LUT_INIT = 16'ha8a0;
    SB_LUT4 i21877_4_lut (.I0(n7_adj_5666), .I1(delay_counter[31]), .I2(n27140), 
            .I3(n8_adj_5665), .O(n1650));   // verilog/TinyFPGA_B.v(389[14:38])
    defparam i21877_4_lut.LUT_INIT = 16'h3230;
    SB_CARRY unary_minus_19_add_3_9 (.CI(n43462), .I0(GND_net), .I1(n18_adj_5470), 
            .CO(n43463));
    SB_LUT4 i2_2_lut (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5659));   // verilog/TinyFPGA_B.v(387[12:17])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 unary_minus_19_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5471), 
            .I3(n43461), .O(n340)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1874 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_5658));   // verilog/TinyFPGA_B.v(387[12:17])
    defparam i6_4_lut_adj_1874.LUT_INIT = 16'hfffe;
    SB_LUT4 add_263_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n43101), .O(encoder1_position_scaled_23__N_75[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_8 (.CI(n43461), .I0(GND_net), .I1(n19_adj_5471), 
            .CO(n43462));
    SB_LUT4 unary_minus_19_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5472), 
            .I3(n43460), .O(n341)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut (.I0(ID[3]), .I1(n14_adj_5658), .I2(n10_adj_5659), 
            .I3(ID[6]), .O(n27117));   // verilog/TinyFPGA_B.v(387[12:17])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_263_23 (.CI(n43101), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n43102));
    SB_CARRY unary_minus_19_add_3_7 (.CI(n43460), .I0(GND_net), .I1(n20_adj_5472), 
            .CO(n43461));
    SB_LUT4 i15099_4_lut (.I0(n7593), .I1(n1650), .I2(n20976), .I3(n27118), 
            .O(n29146));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    defparam i15099_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i5050_2_lut (.I0(n2_adj_5509), .I1(encoder0_position_scaled_23__N_327[31]), 
            .I2(GND_net), .I3(GND_net), .O(n621));
    defparam i5050_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i500_4_lut (.I0(n621), .I1(n8584), 
            .I2(n51706), .I3(n5_adj_5482), .O(n828));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i500_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_6_lut (.I0(GND_net), 
            .I1(n2030), .I2(GND_net), .I3(n43654), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_6 (.CI(n43654), 
            .I0(n2030), .I1(GND_net), .CO(n43655));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_5_lut (.I0(GND_net), 
            .I1(n2031), .I2(VCC_net), .I3(n43653), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5473), 
            .I3(n43459), .O(n342)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_6 (.CI(n43459), .I0(GND_net), .I1(n21_adj_5473), 
            .CO(n43460));
    SB_LUT4 i21658_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(91[16:31])
    defparam i21658_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21657_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(89[16:31])
    defparam i21657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21656_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(87[16:31])
    defparam i21656_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_5 (.CI(n43653), 
            .I0(n2031), .I1(VCC_net), .CO(n43654));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_4_lut (.I0(GND_net), 
            .I1(n2032), .I2(GND_net), .I3(n43652), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_4 (.CI(n43652), 
            .I0(n2032), .I1(GND_net), .CO(n43653));
    SB_LUT4 unary_minus_19_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5474), 
            .I3(n43458), .O(n343)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_3_lut (.I0(GND_net), 
            .I1(n2033), .I2(VCC_net), .I3(n43651), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_3 (.CI(n43651), 
            .I0(n2033), .I1(VCC_net), .CO(n43652));
    SB_CARRY unary_minus_19_add_3_5 (.CI(n43458), .I0(GND_net), .I1(n22_adj_5474), 
            .CO(n43459));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1369_2_lut (.I0(GND_net), 
            .I1(n531), .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1369_2 (.CI(VCC_net), 
            .I0(n531), .I1(GND_net), .CO(n43651));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_19_lut (.I0(n56055), 
            .I1(n1917), .I2(VCC_net), .I3(n43650), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_18_lut (.I0(GND_net), 
            .I1(n1918), .I2(VCC_net), .I3(n43649), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_18 (.CI(n43649), 
            .I0(n1918), .I1(VCC_net), .CO(n43650));
    SB_LUT4 unary_minus_19_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5475), 
            .I3(n43457), .O(n344)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_4 (.CI(n43457), .I0(GND_net), .I1(n23_adj_5475), 
            .CO(n43458));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_17_lut (.I0(GND_net), 
            .I1(n1919), .I2(VCC_net), .I3(n43648), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_17 (.CI(n43648), 
            .I0(n1919), .I1(VCC_net), .CO(n43649));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_16_lut (.I0(GND_net), 
            .I1(n1920), .I2(VCC_net), .I3(n43647), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_16 (.CI(n43647), 
            .I0(n1920), .I1(VCC_net), .CO(n43648));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_15_lut (.I0(GND_net), 
            .I1(n1921), .I2(VCC_net), .I3(n43646), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_15 (.CI(n43646), 
            .I0(n1921), .I1(VCC_net), .CO(n43647));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_14_lut (.I0(GND_net), 
            .I1(n1922), .I2(VCC_net), .I3(n43645), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2279_add_4_9_lut (.I0(n54247), .I1(n35823), .I2(dti_counter[7]), 
            .I3(n43993), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 dti_counter_2279_add_4_8_lut (.I0(n54248), .I1(n35823), .I2(dti_counter[6]), 
            .I3(n43992), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 unary_minus_19_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5476), 
            .I3(n43456), .O(n345)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2279_add_4_8 (.CI(n43992), .I0(n35823), .I1(dti_counter[6]), 
            .CO(n43993));
    SB_CARRY unary_minus_19_add_3_3 (.CI(n43456), .I0(GND_net), .I1(n24_adj_5476), 
            .CO(n43457));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_14 (.CI(n43645), 
            .I0(n1922), .I1(VCC_net), .CO(n43646));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_13_lut (.I0(GND_net), 
            .I1(n1923), .I2(VCC_net), .I3(n43644), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n25_adj_5477), 
            .I3(VCC_net), .O(n54237)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 dti_counter_2279_add_4_7_lut (.I0(n54249), .I1(n35823), .I2(dti_counter[5]), 
            .I3(n43991), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2279_add_4_7 (.CI(n43991), .I0(n35823), .I1(dti_counter[5]), 
            .CO(n43992));
    SB_CARRY unary_minus_19_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5477), 
            .CO(n43456));
    SB_LUT4 dti_counter_2279_add_4_6_lut (.I0(n54250), .I1(n35823), .I2(dti_counter[4]), 
            .I3(n43990), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 add_5097_32_lut (.I0(GND_net), .I1(encoder0_position[31]), .I2(VCC_net), 
            .I3(n43455), .O(encoder0_position_scaled_23__N_327[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2279_add_4_6 (.CI(n43990), .I0(n35823), .I1(dti_counter[4]), 
            .CO(n43991));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_13 (.CI(n43644), 
            .I0(n1923), .I1(VCC_net), .CO(n43645));
    SB_LUT4 dti_counter_2279_add_4_5_lut (.I0(n54251), .I1(n35823), .I2(dti_counter[3]), 
            .I3(n43989), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2279_add_4_5 (.CI(n43989), .I0(n35823), .I1(dti_counter[3]), 
            .CO(n43990));
    SB_LUT4 add_263_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n43100), .O(encoder1_position_scaled_23__N_75[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2279_add_4_4_lut (.I0(n54252), .I1(n35823), .I2(dti_counter[2]), 
            .I3(n43988), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 add_5097_31_lut (.I0(GND_net), .I1(encoder0_position[30]), .I2(VCC_net), 
            .I3(n43454), .O(encoder0_position_scaled_23__N_327[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_31 (.CI(n43454), .I0(encoder0_position[30]), .I1(VCC_net), 
            .CO(n43455));
    SB_LUT4 add_5097_30_lut (.I0(GND_net), .I1(encoder0_position[29]), .I2(VCC_net), 
            .I3(n43453), .O(encoder0_position_scaled_23__N_327[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_12_lut (.I0(GND_net), 
            .I1(n1924), .I2(VCC_net), .I3(n43643), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2279_add_4_4 (.CI(n43988), .I0(n35823), .I1(dti_counter[2]), 
            .CO(n43989));
    SB_LUT4 dti_counter_2279_add_4_3_lut (.I0(n54253), .I1(n35823), .I2(dti_counter[1]), 
            .I3(n43987), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_12 (.CI(n43643), 
            .I0(n1924), .I1(VCC_net), .CO(n43644));
    SB_CARRY dti_counter_2279_add_4_3 (.CI(n43987), .I0(n35823), .I1(dti_counter[1]), 
            .CO(n43988));
    SB_LUT4 dti_counter_2279_add_4_2_lut (.I0(n54290), .I1(n2573), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2279_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY dti_counter_2279_add_4_2 (.CI(VCC_net), .I0(n2573), .I1(dti_counter[0]), 
            .CO(n43987));
    SB_LUT4 add_2800_25_lut (.I0(n56209), .I1(n2_adj_5618), .I2(n1059), 
            .I3(n43986), .O(encoder0_position_scaled_23__N_51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2800_24_lut (.I0(n56195), .I1(n2_adj_5618), .I2(n1158), 
            .I3(n43985), .O(encoder0_position_scaled_23__N_51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_24 (.CI(n43985), .I0(n2_adj_5618), .I1(n1158), .CO(n43986));
    SB_LUT4 add_2800_23_lut (.I0(n56181), .I1(n2_adj_5618), .I2(n1257), 
            .I3(n43984), .O(encoder0_position_scaled_23__N_51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_11_lut (.I0(GND_net), 
            .I1(n1925), .I2(VCC_net), .I3(n43642), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_23 (.CI(n43984), .I0(n2_adj_5618), .I1(n1257), .CO(n43985));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_11 (.CI(n43642), 
            .I0(n1925), .I1(VCC_net), .CO(n43643));
    SB_LUT4 add_2800_22_lut (.I0(n56167), .I1(n2_adj_5618), .I2(n1356), 
            .I3(n43983), .O(encoder0_position_scaled_23__N_51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_22 (.CI(n43983), .I0(n2_adj_5618), .I1(n1356), .CO(n43984));
    SB_LUT4 add_2800_21_lut (.I0(n56150), .I1(n2_adj_5618), .I2(n1455), 
            .I3(n43982), .O(encoder0_position_scaled_23__N_51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i971_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2800_21 (.CI(n43982), .I0(n2_adj_5618), .I1(n1455), .CO(n43983));
    SB_CARRY add_5097_30 (.CI(n43453), .I0(encoder0_position[29]), .I1(VCC_net), 
            .CO(n43454));
    SB_LUT4 add_2800_20_lut (.I0(n56120), .I1(n2_adj_5618), .I2(n1554_adj_5610), 
            .I3(n43981), .O(encoder0_position_scaled_23__N_51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_20 (.CI(n43981), .I0(n2_adj_5618), .I1(n1554_adj_5610), 
            .CO(n43982));
    SB_LUT4 add_2800_19_lut (.I0(n56116), .I1(n2_adj_5618), .I2(n1653), 
            .I3(n43980), .O(encoder0_position_scaled_23__N_51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_19 (.CI(n43980), .I0(n2_adj_5618), .I1(n1653), .CO(n43981));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_10_lut (.I0(GND_net), 
            .I1(n1926), .I2(VCC_net), .I3(n43641), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_10 (.CI(n43641), 
            .I0(n1926), .I1(VCC_net), .CO(n43642));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2800_18_lut (.I0(n56096), .I1(n2_adj_5618), .I2(n1752), 
            .I3(n43979), .O(encoder0_position_scaled_23__N_51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_18 (.CI(n43979), .I0(n2_adj_5618), .I1(n1752), .CO(n43980));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_9_lut (.I0(GND_net), 
            .I1(n1927), .I2(VCC_net), .I3(n43640), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2800_17_lut (.I0(n56075), .I1(n2_adj_5618), .I2(n1851), 
            .I3(n43978), .O(encoder0_position_scaled_23__N_51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_17 (.CI(n43978), .I0(n2_adj_5618), .I1(n1851), .CO(n43979));
    SB_LUT4 add_2800_16_lut (.I0(n56055), .I1(n2_adj_5618), .I2(n1950), 
            .I3(n43977), .O(encoder0_position_scaled_23__N_51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_16 (.CI(n43977), .I0(n2_adj_5618), .I1(n1950), .CO(n43978));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_9 (.CI(n43640), 
            .I0(n1927), .I1(VCC_net), .CO(n43641));
    SB_LUT4 add_5097_29_lut (.I0(GND_net), .I1(encoder0_position[28]), .I2(VCC_net), 
            .I3(n43452), .O(encoder0_position_scaled_23__N_327[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2800_15_lut (.I0(n56033), .I1(n2_adj_5618), .I2(n2049), 
            .I3(n43976), .O(encoder0_position_scaled_23__N_51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_8_lut (.I0(GND_net), 
            .I1(n1928), .I2(VCC_net), .I3(n43639), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_15 (.CI(n43976), .I0(n2_adj_5618), .I1(n2049), .CO(n43977));
    SB_LUT4 add_2800_14_lut (.I0(n56010), .I1(n2_adj_5618), .I2(n2148), 
            .I3(n43975), .O(encoder0_position_scaled_23__N_51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i841_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_8 (.CI(n43639), 
            .I0(n1928), .I1(VCC_net), .CO(n43640));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_7_lut (.I0(GND_net), 
            .I1(n1929), .I2(GND_net), .I3(n43638), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_7 (.CI(n43638), 
            .I0(n1929), .I1(GND_net), .CO(n43639));
    SB_CARRY add_2800_14 (.CI(n43975), .I0(n2_adj_5618), .I1(n2148), .CO(n43976));
    SB_LUT4 add_2800_13_lut (.I0(n55986), .I1(n2_adj_5618), .I2(n2247), 
            .I3(n43974), .O(encoder0_position_scaled_23__N_51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_13 (.CI(n43974), .I0(n2_adj_5618), .I1(n2247), .CO(n43975));
    SB_LUT4 add_2800_12_lut (.I0(n55960), .I1(n2_adj_5618), .I2(n2346), 
            .I3(n43973), .O(encoder0_position_scaled_23__N_51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_12 (.CI(n43973), .I0(n2_adj_5618), .I1(n2346), .CO(n43974));
    SB_LUT4 add_2800_11_lut (.I0(n55935), .I1(n2_adj_5618), .I2(n2445), 
            .I3(n43972), .O(encoder0_position_scaled_23__N_51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_11 (.CI(n43972), .I0(n2_adj_5618), .I1(n2445), .CO(n43973));
    SB_LUT4 add_2800_10_lut (.I0(n55883), .I1(n2_adj_5618), .I2(n2544), 
            .I3(n43971), .O(encoder0_position_scaled_23__N_51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_10 (.CI(n43971), .I0(n2_adj_5618), .I1(n2544), .CO(n43972));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_6_lut (.I0(GND_net), 
            .I1(n1930), .I2(GND_net), .I3(n43637), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_29 (.CI(n43452), .I0(encoder0_position[28]), .I1(VCC_net), 
            .CO(n43453));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_6 (.CI(n43637), 
            .I0(n1930), .I1(GND_net), .CO(n43638));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_5_lut (.I0(GND_net), 
            .I1(n1931), .I2(VCC_net), .I3(n43636), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2800_9_lut (.I0(n55879), .I1(n2_adj_5618), .I2(n2643), 
            .I3(n43970), .O(encoder0_position_scaled_23__N_51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_9 (.CI(n43970), .I0(n2_adj_5618), .I1(n2643), .CO(n43971));
    SB_LUT4 add_2800_8_lut (.I0(n55850), .I1(n2_adj_5618), .I2(n2742), 
            .I3(n43969), .O(encoder0_position_scaled_23__N_51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_8 (.CI(n43969), .I0(n2_adj_5618), .I1(n2742), .CO(n43970));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_5 (.CI(n43636), 
            .I0(n1931), .I1(VCC_net), .CO(n43637));
    SB_LUT4 add_2800_7_lut (.I0(n55819), .I1(n2_adj_5618), .I2(n2841), 
            .I3(n43968), .O(encoder0_position_scaled_23__N_51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_7 (.CI(n43968), .I0(n2_adj_5618), .I1(n2841), .CO(n43969));
    SB_LUT4 add_2800_6_lut (.I0(n55788), .I1(n2_adj_5618), .I2(n2940), 
            .I3(n43967), .O(encoder0_position_scaled_23__N_51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_6 (.CI(n43967), .I0(n2_adj_5618), .I1(n2940), .CO(n43968));
    SB_LUT4 add_2800_5_lut (.I0(n55756), .I1(n2_adj_5618), .I2(n3039), 
            .I3(n43966), .O(encoder0_position_scaled_23__N_51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_4_lut (.I0(GND_net), 
            .I1(n1932), .I2(GND_net), .I3(n43635), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_4 (.CI(n43635), 
            .I0(n1932), .I1(GND_net), .CO(n43636));
    SB_CARRY add_2800_5 (.CI(n43966), .I0(n2_adj_5618), .I1(n3039), .CO(n43967));
    SB_LUT4 add_2800_4_lut (.I0(n55724), .I1(n2_adj_5618), .I2(n3138), 
            .I3(n43965), .O(encoder0_position_scaled_23__N_51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_4 (.CI(n43965), .I0(n2_adj_5618), .I1(n3138), .CO(n43966));
    SB_LUT4 add_5097_28_lut (.I0(GND_net), .I1(encoder0_position[27]), .I2(VCC_net), 
            .I3(n43451), .O(encoder0_position_scaled_23__N_327[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_28 (.CI(n43451), .I0(encoder0_position[27]), .I1(VCC_net), 
            .CO(n43452));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_3_lut (.I0(GND_net), 
            .I1(n1933), .I2(VCC_net), .I3(n43634), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_3 (.CI(n43634), 
            .I0(n1933), .I1(VCC_net), .CO(n43635));
    SB_LUT4 add_2800_3_lut (.I0(n56270), .I1(n2_adj_5618), .I2(n3237), 
            .I3(n43964), .O(encoder0_position_scaled_23__N_51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1302_2_lut (.I0(GND_net), 
            .I1(n530), .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5097_27_lut (.I0(GND_net), .I1(encoder0_position[26]), .I2(VCC_net), 
            .I3(n43450), .O(encoder0_position_scaled_23__N_327[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_27 (.CI(n43450), .I0(encoder0_position[26]), .I1(VCC_net), 
            .CO(n43451));
    SB_LUT4 add_5097_26_lut (.I0(GND_net), .I1(encoder0_position[25]), .I2(VCC_net), 
            .I3(n43449), .O(encoder0_position_scaled_23__N_327[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_26 (.CI(n43449), .I0(encoder0_position[25]), .I1(VCC_net), 
            .CO(n43450));
    SB_LUT4 add_5097_25_lut (.I0(GND_net), .I1(encoder0_position[24]), .I2(VCC_net), 
            .I3(n43448), .O(encoder0_position_scaled_23__N_327[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_3 (.CI(n43964), .I0(n2_adj_5618), .I1(n3237), .CO(n43965));
    SB_LUT4 add_2800_2_lut (.I0(n56237), .I1(n2_adj_5618), .I2(n36808), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2800_2 (.CI(VCC_net), .I0(n2_adj_5618), .I1(n36808), 
            .CO(n43964));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_33_lut (.I0(GND_net), 
            .I1(n3204), .I2(VCC_net), .I3(n43963), .O(n3271)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_25 (.CI(n43448), .I0(encoder0_position[24]), .I1(VCC_net), 
            .CO(n43449));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1302_2 (.CI(VCC_net), 
            .I0(n530), .I1(GND_net), .CO(n43634));
    SB_LUT4 add_5097_24_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(VCC_net), 
            .I3(n43447), .O(encoder0_position_scaled_23__N_327[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_32_lut (.I0(GND_net), 
            .I1(n3205), .I2(VCC_net), .I3(n43962), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_24 (.CI(n43447), .I0(encoder0_position[23]), .I1(VCC_net), 
            .CO(n43448));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_32 (.CI(n43962), 
            .I0(n3205), .I1(VCC_net), .CO(n43963));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_31_lut (.I0(GND_net), 
            .I1(n3206), .I2(VCC_net), .I3(n43961), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_18_lut (.I0(n56075), 
            .I1(n1818), .I2(VCC_net), .I3(n43633), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_17_lut (.I0(GND_net), 
            .I1(n1819), .I2(VCC_net), .I3(n43632), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5097_23_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(VCC_net), 
            .I3(n43446), .O(encoder0_position_scaled_23__N_327[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_23 (.CI(n43446), .I0(encoder0_position[22]), .I1(VCC_net), 
            .CO(n43447));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_31 (.CI(n43961), 
            .I0(n3206), .I1(VCC_net), .CO(n43962));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_17 (.CI(n43632), 
            .I0(n1819), .I1(VCC_net), .CO(n43633));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_16_lut (.I0(GND_net), 
            .I1(n1820), .I2(VCC_net), .I3(n43631), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_16 (.CI(n43631), 
            .I0(n1820), .I1(VCC_net), .CO(n43632));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_30_lut (.I0(GND_net), 
            .I1(n3207), .I2(VCC_net), .I3(n43960), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5097_22_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(VCC_net), 
            .I3(n43445), .O(encoder0_position_scaled_23__N_327[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_15_lut (.I0(GND_net), 
            .I1(n1821), .I2(VCC_net), .I3(n43630), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_30 (.CI(n43960), 
            .I0(n3207), .I1(VCC_net), .CO(n43961));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_29_lut (.I0(GND_net), 
            .I1(n3208), .I2(VCC_net), .I3(n43959), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_22 (.CI(n43445), .I0(encoder0_position[21]), .I1(VCC_net), 
            .CO(n43446));
    SB_LUT4 add_5097_21_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(VCC_net), 
            .I3(n43444), .O(encoder0_position_scaled_23__N_327[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_15 (.CI(n43630), 
            .I0(n1821), .I1(VCC_net), .CO(n43631));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_29 (.CI(n43959), 
            .I0(n3208), .I1(VCC_net), .CO(n43960));
    SB_CARRY add_5097_21 (.CI(n43444), .I0(encoder0_position[20]), .I1(VCC_net), 
            .CO(n43445));
    SB_LUT4 add_5097_20_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(VCC_net), 
            .I3(n43443), .O(encoder0_position_scaled_23__N_327[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_20 (.CI(n43443), .I0(encoder0_position[19]), .I1(VCC_net), 
            .CO(n43444));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_28_lut (.I0(GND_net), 
            .I1(n3209), .I2(VCC_net), .I3(n43958), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_28 (.CI(n43958), 
            .I0(n3209), .I1(VCC_net), .CO(n43959));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_27_lut (.I0(GND_net), 
            .I1(n3210), .I2(VCC_net), .I3(n43957), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_14_lut (.I0(GND_net), 
            .I1(n1822), .I2(VCC_net), .I3(n43629), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_14 (.CI(n43629), 
            .I0(n1822), .I1(VCC_net), .CO(n43630));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_13_lut (.I0(GND_net), 
            .I1(n1823), .I2(VCC_net), .I3(n43628), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5097_19_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(VCC_net), 
            .I3(n43442), .O(encoder0_position_scaled_23__N_327[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_27 (.CI(n43957), 
            .I0(n3210), .I1(VCC_net), .CO(n43958));
    SB_CARRY add_5097_19 (.CI(n43442), .I0(encoder0_position[18]), .I1(VCC_net), 
            .CO(n43443));
    SB_LUT4 add_5097_18_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(VCC_net), 
            .I3(n43441), .O(encoder0_position_scaled_23__N_327[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_26_lut (.I0(GND_net), 
            .I1(n3211), .I2(VCC_net), .I3(n43956), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_26 (.CI(n43956), 
            .I0(n3211), .I1(VCC_net), .CO(n43957));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_13 (.CI(n43628), 
            .I0(n1823), .I1(VCC_net), .CO(n43629));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_25_lut (.I0(GND_net), 
            .I1(n3212), .I2(VCC_net), .I3(n43955), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_18 (.CI(n43441), .I0(encoder0_position[17]), .I1(VCC_net), 
            .CO(n43442));
    SB_LUT4 add_5097_17_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(VCC_net), 
            .I3(n43440), .O(encoder0_position_scaled_23__N_327[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_12_lut (.I0(GND_net), 
            .I1(n1824), .I2(VCC_net), .I3(n43627), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_17 (.CI(n43440), .I0(encoder0_position[16]), .I1(VCC_net), 
            .CO(n43441));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_12 (.CI(n43627), 
            .I0(n1824), .I1(VCC_net), .CO(n43628));
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(clk16MHz), .D(n29257));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_LUT4 add_5097_16_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(VCC_net), 
            .I3(n43439), .O(encoder0_position_scaled_23__N_327[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_16 (.CI(n43439), .I0(encoder0_position[15]), .I1(VCC_net), 
            .CO(n43440));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_25 (.CI(n43955), 
            .I0(n3212), .I1(VCC_net), .CO(n43956));
    SB_LUT4 add_5097_15_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(VCC_net), 
            .I3(n43438), .O(encoder0_position_scaled_23__N_327[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_24_lut (.I0(GND_net), 
            .I1(n3213), .I2(VCC_net), .I3(n43954), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_15 (.CI(n43438), .I0(encoder0_position[14]), .I1(VCC_net), 
            .CO(n43439));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_24 (.CI(n43954), 
            .I0(n3213), .I1(VCC_net), .CO(n43955));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_23_lut (.I0(GND_net), 
            .I1(n3214), .I2(VCC_net), .I3(n43953), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5097_14_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(VCC_net), 
            .I3(n43437), .O(encoder0_position_scaled_23__N_327[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_14 (.CI(n43437), .I0(encoder0_position[13]), .I1(VCC_net), 
            .CO(n43438));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_23 (.CI(n43953), 
            .I0(n3214), .I1(VCC_net), .CO(n43954));
    SB_LUT4 add_5097_13_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(VCC_net), 
            .I3(n43436), .O(encoder0_position_scaled_23__N_327[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_22_lut (.I0(GND_net), 
            .I1(n3215), .I2(VCC_net), .I3(n43952), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_22 (.CI(n43952), 
            .I0(n3215), .I1(VCC_net), .CO(n43953));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_21_lut (.I0(GND_net), 
            .I1(n3216), .I2(VCC_net), .I3(n43951), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_21 (.CI(n43951), 
            .I0(n3216), .I1(VCC_net), .CO(n43952));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_11_lut (.I0(GND_net), 
            .I1(n1825), .I2(VCC_net), .I3(n43626), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_11 (.CI(n43626), 
            .I0(n1825), .I1(VCC_net), .CO(n43627));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_10_lut (.I0(GND_net), 
            .I1(n1826), .I2(VCC_net), .I3(n43625), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_10 (.CI(n43625), 
            .I0(n1826), .I1(VCC_net), .CO(n43626));
    SB_CARRY add_5097_13 (.CI(n43436), .I0(encoder0_position[12]), .I1(VCC_net), 
            .CO(n43437));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_20_lut (.I0(GND_net), 
            .I1(n3217), .I2(VCC_net), .I3(n43950), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_9_lut (.I0(GND_net), 
            .I1(n1827), .I2(VCC_net), .I3(n43624), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_20 (.CI(n43950), 
            .I0(n3217), .I1(VCC_net), .CO(n43951));
    SB_LUT4 add_5097_12_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(VCC_net), 
            .I3(n43435), .O(encoder0_position_scaled_23__N_327[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_19_lut (.I0(GND_net), 
            .I1(n3218), .I2(VCC_net), .I3(n43949), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_19 (.CI(n43949), 
            .I0(n3218), .I1(VCC_net), .CO(n43950));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_9 (.CI(n43624), 
            .I0(n1827), .I1(VCC_net), .CO(n43625));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_18_lut (.I0(GND_net), 
            .I1(n3219), .I2(VCC_net), .I3(n43948), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_8_lut (.I0(GND_net), 
            .I1(n1828), .I2(VCC_net), .I3(n43623), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_8 (.CI(n43623), 
            .I0(n1828), .I1(VCC_net), .CO(n43624));
    SB_CARRY add_5097_12 (.CI(n43435), .I0(encoder0_position[11]), .I1(VCC_net), 
            .CO(n43436));
    SB_LUT4 add_5097_11_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(VCC_net), 
            .I3(n43434), .O(encoder0_position_scaled_23__N_327[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_11 (.CI(n43434), .I0(encoder0_position[10]), .I1(VCC_net), 
            .CO(n43435));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_18 (.CI(n43948), 
            .I0(n3219), .I1(VCC_net), .CO(n43949));
    SB_LUT4 add_5097_10_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(VCC_net), 
            .I3(n43433), .O(encoder0_position_scaled_23__N_327[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_17_lut (.I0(GND_net), 
            .I1(n3220), .I2(VCC_net), .I3(n43947), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_17 (.CI(n43947), 
            .I0(n3220), .I1(VCC_net), .CO(n43948));
    SB_CARRY add_5097_10 (.CI(n43433), .I0(encoder0_position[9]), .I1(VCC_net), 
            .CO(n43434));
    SB_LUT4 add_5097_9_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(VCC_net), 
            .I3(n43432), .O(encoder0_position_scaled_23__N_327[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_9 (.CI(n43432), .I0(encoder0_position[8]), .I1(VCC_net), 
            .CO(n43433));
    SB_LUT4 add_5097_8_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(VCC_net), 
            .I3(n43431), .O(encoder0_position_scaled_23__N_327[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_8 (.CI(n43431), .I0(encoder0_position[7]), .I1(VCC_net), 
            .CO(n43432));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_16_lut (.I0(GND_net), 
            .I1(n3221), .I2(VCC_net), .I3(n43946), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_7_lut (.I0(GND_net), 
            .I1(n1829), .I2(GND_net), .I3(n43622), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_16 (.CI(n43946), 
            .I0(n3221), .I1(VCC_net), .CO(n43947));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_15_lut (.I0(GND_net), 
            .I1(n3222), .I2(VCC_net), .I3(n43945), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5097_7_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(VCC_net), 
            .I3(n43430), .O(encoder0_position_scaled_23__N_327[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_15 (.CI(n43945), 
            .I0(n3222), .I1(VCC_net), .CO(n43946));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_14_lut (.I0(GND_net), 
            .I1(n3223), .I2(VCC_net), .I3(n43944), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_7 (.CI(n43430), .I0(encoder0_position[6]), .I1(VCC_net), 
            .CO(n43431));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_7 (.CI(n43622), 
            .I0(n1829), .I1(GND_net), .CO(n43623));
    SB_LUT4 add_5097_6_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(VCC_net), 
            .I3(n43429), .O(encoder0_position_scaled_23__N_327[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_14 (.CI(n43944), 
            .I0(n3223), .I1(VCC_net), .CO(n43945));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_6_lut (.I0(GND_net), 
            .I1(n1830), .I2(GND_net), .I3(n43621), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_6 (.CI(n43429), .I0(encoder0_position[5]), .I1(VCC_net), 
            .CO(n43430));
    SB_LUT4 add_5097_5_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(VCC_net), 
            .I3(n43428), .O(encoder0_position_scaled_23__N_327[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_6 (.CI(n43621), 
            .I0(n1830), .I1(GND_net), .CO(n43622));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_13_lut (.I0(GND_net), 
            .I1(n3224), .I2(VCC_net), .I3(n43943), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_5_lut (.I0(GND_net), 
            .I1(n1831), .I2(VCC_net), .I3(n43620), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_5 (.CI(n43620), 
            .I0(n1831), .I1(VCC_net), .CO(n43621));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_13 (.CI(n43943), 
            .I0(n3224), .I1(VCC_net), .CO(n43944));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_12_lut (.I0(GND_net), 
            .I1(n3225), .I2(VCC_net), .I3(n43942), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_4_lut (.I0(GND_net), 
            .I1(n1832), .I2(GND_net), .I3(n43619), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_5 (.CI(n43428), .I0(encoder0_position[4]), .I1(VCC_net), 
            .CO(n43429));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_4 (.CI(n43619), 
            .I0(n1832), .I1(GND_net), .CO(n43620));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_12 (.CI(n43942), 
            .I0(n3225), .I1(VCC_net), .CO(n43943));
    SB_LUT4 add_5097_4_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(VCC_net), 
            .I3(n43427), .O(encoder0_position_scaled_23__N_327[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_4 (.CI(n43427), .I0(encoder0_position[3]), .I1(VCC_net), 
            .CO(n43428));
    SB_LUT4 add_5097_3_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(VCC_net), 
            .I3(n43426), .O(encoder0_position_scaled_23__N_327[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5097_3 (.CI(n43426), .I0(encoder0_position[2]), .I1(VCC_net), 
            .CO(n43427));
    SB_LUT4 add_5097_2_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(VCC_net), 
            .I3(n43425), .O(encoder0_position_scaled_23__N_327[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5097_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_11_lut (.I0(GND_net), 
            .I1(n3226), .I2(VCC_net), .I3(n43941), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_3_lut (.I0(GND_net), 
            .I1(n1833), .I2(VCC_net), .I3(n43618), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_11 (.CI(n43941), 
            .I0(n3226), .I1(VCC_net), .CO(n43942));
    SB_CARRY add_5097_2 (.CI(n43425), .I0(encoder0_position[1]), .I1(VCC_net), 
            .CO(n43426));
    SB_CARRY add_5097_1 (.CI(GND_net), .I0(encoder0_position[0]), .I1(encoder0_position[0]), 
            .CO(n43425));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_10_lut (.I0(GND_net), 
            .I1(n3227), .I2(VCC_net), .I3(n43940), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_3 (.CI(n43618), 
            .I0(n1833), .I1(VCC_net), .CO(n43619));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1235_2_lut (.I0(GND_net), 
            .I1(n529), .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1235_2 (.CI(VCC_net), 
            .I0(n529), .I1(GND_net), .CO(n43618));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_10 (.CI(n43940), 
            .I0(n3227), .I1(VCC_net), .CO(n43941));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1038_3_lut (.I0(n1523), 
            .I1(n1590), .I2(n1554_adj_5610), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_9_lut (.I0(GND_net), 
            .I1(n3228), .I2(VCC_net), .I3(n43939), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_9 (.CI(n43939), 
            .I0(n3228), .I1(VCC_net), .CO(n43940));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_8_lut (.I0(GND_net), 
            .I1(n3229), .I2(GND_net), .I3(n43938), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLA_211 (.Q(INLA_c_0), .C(clk16MHz), .E(n28583), .D(GLA_N_495), 
            .R(n29049));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1105_3_lut (.I0(n1622), 
            .I1(n1689), .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_8 (.CI(n43938), 
            .I0(n3229), .I1(GND_net), .CO(n43939));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_7_lut (.I0(n3298), 
            .I1(n3230), .I2(GND_net), .I3(n43937), .O(n54294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_7 (.CI(n43937), 
            .I0(n3230), .I1(GND_net), .CO(n43938));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_17_lut (.I0(n56096), 
            .I1(n1719), .I2(VCC_net), .I3(n43617), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_16_lut (.I0(GND_net), 
            .I1(n1720), .I2(VCC_net), .I3(n43616), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_6_lut (.I0(GND_net), 
            .I1(n3231), .I2(VCC_net), .I3(n43936), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i975_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_6 (.CI(n43936), 
            .I0(n3231), .I1(VCC_net), .CO(n43937));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_5_lut (.I0(GND_net), 
            .I1(n3232), .I2(GND_net), .I3(n43935), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLB_213 (.Q(INLB_c_0), .C(clk16MHz), .E(n28583), .D(GLB_N_509), 
            .R(n29049));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_16 (.CI(n43616), 
            .I0(n1720), .I1(VCC_net), .CO(n43617));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_15_lut (.I0(GND_net), 
            .I1(n1721), .I2(VCC_net), .I3(n43615), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_15 (.CI(n43615), 
            .I0(n1721), .I1(VCC_net), .CO(n43616));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_14_lut (.I0(GND_net), 
            .I1(n1722), .I2(VCC_net), .I3(n43614), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_14 (.CI(n43614), 
            .I0(n1722), .I1(VCC_net), .CO(n43615));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_5 (.CI(n43935), 
            .I0(n3232), .I1(GND_net), .CO(n43936));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_4_lut (.I0(GND_net), 
            .I1(n3233), .I2(VCC_net), .I3(n43934), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_13_lut (.I0(GND_net), 
            .I1(n1723), .I2(VCC_net), .I3(n43613), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_22 (.CI(n43100), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n43101));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_4 (.CI(n43934), 
            .I0(n3233), .I1(VCC_net), .CO(n43935));
    SB_LUT4 add_263_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n43099), .O(encoder1_position_scaled_23__N_75[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2173_3_lut (.I0(GND_net), 
            .I1(n543), .I2(GND_net), .I3(n43933), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_3 (.CI(n43933), 
            .I0(n543), .I1(GND_net), .CO(n43934));
    SB_CARRY add_263_3 (.CI(n43081), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n43082));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2173_2 (.CI(VCC_net), 
            .I0(n544), .I1(VCC_net), .CO(n43933));
    SB_LUT4 add_263_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n43087), .O(encoder1_position_scaled_23__N_75[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_31_lut (.I0(n55724), 
            .I1(n3105), .I2(VCC_net), .I3(n43932), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_30_lut (.I0(GND_net), 
            .I1(n3106), .I2(VCC_net), .I3(n43931), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_30 (.CI(n43931), 
            .I0(n3106), .I1(VCC_net), .CO(n43932));
    SB_CARRY add_263_21 (.CI(n43099), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n43100));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_29_lut (.I0(GND_net), 
            .I1(n3107), .I2(VCC_net), .I3(n43930), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_13 (.CI(n43613), 
            .I0(n1723), .I1(VCC_net), .CO(n43614));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_29 (.CI(n43930), 
            .I0(n3107), .I1(VCC_net), .CO(n43931));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_12_lut (.I0(GND_net), 
            .I1(n1724), .I2(VCC_net), .I3(n43612), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_12 (.CI(n43612), 
            .I0(n1724), .I1(VCC_net), .CO(n43613));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_28_lut (.I0(GND_net), 
            .I1(n3108), .I2(VCC_net), .I3(n43929), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_11_lut (.I0(GND_net), 
            .I1(n1725), .I2(VCC_net), .I3(n43611), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_11 (.CI(n43611), 
            .I0(n1725), .I1(VCC_net), .CO(n43612));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_10_lut (.I0(GND_net), 
            .I1(n1726), .I2(VCC_net), .I3(n43610), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_28 (.CI(n43929), 
            .I0(n3108), .I1(VCC_net), .CO(n43930));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_27_lut (.I0(GND_net), 
            .I1(n3109), .I2(VCC_net), .I3(n43928), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_27 (.CI(n43928), 
            .I0(n3109), .I1(VCC_net), .CO(n43929));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_26_lut (.I0(GND_net), 
            .I1(n3110), .I2(VCC_net), .I3(n43927), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_26 (.CI(n43927), 
            .I0(n3110), .I1(VCC_net), .CO(n43928));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_25_lut (.I0(GND_net), 
            .I1(n3111), .I2(VCC_net), .I3(n43926), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_10 (.CI(n43610), 
            .I0(n1726), .I1(VCC_net), .CO(n43611));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_9_lut (.I0(GND_net), 
            .I1(n1727), .I2(VCC_net), .I3(n43609), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_25 (.CI(n43926), 
            .I0(n3111), .I1(VCC_net), .CO(n43927));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_24_lut (.I0(GND_net), 
            .I1(n3112), .I2(VCC_net), .I3(n43925), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_9 (.CI(n43609), 
            .I0(n1727), .I1(VCC_net), .CO(n43610));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_8_lut (.I0(GND_net), 
            .I1(n1728), .I2(VCC_net), .I3(n43608), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_8 (.CI(n43608), 
            .I0(n1728), .I1(VCC_net), .CO(n43609));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_24 (.CI(n43925), 
            .I0(n3112), .I1(VCC_net), .CO(n43926));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1042_3_lut (.I0(n1527), 
            .I1(n1594), .I2(n1554_adj_5610), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_23_lut (.I0(GND_net), 
            .I1(n3113), .I2(VCC_net), .I3(n43924), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_7_lut (.I0(GND_net), 
            .I1(n1729), .I2(GND_net), .I3(n43607), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_23 (.CI(n43924), 
            .I0(n3113), .I1(VCC_net), .CO(n43925));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_22_lut (.I0(GND_net), 
            .I1(n3114), .I2(VCC_net), .I3(n43923), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_22 (.CI(n43923), 
            .I0(n3114), .I1(VCC_net), .CO(n43924));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_21_lut (.I0(GND_net), 
            .I1(n3115), .I2(VCC_net), .I3(n43922), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_7 (.CI(n43607), 
            .I0(n1729), .I1(GND_net), .CO(n43608));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_21 (.CI(n43922), 
            .I0(n3115), .I1(VCC_net), .CO(n43923));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_20_lut (.I0(GND_net), 
            .I1(n3116), .I2(VCC_net), .I3(n43921), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_20 (.CI(n43921), 
            .I0(n3116), .I1(VCC_net), .CO(n43922));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_19_lut (.I0(GND_net), 
            .I1(n3117), .I2(VCC_net), .I3(n43920), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_6_lut (.I0(GND_net), 
            .I1(n1730), .I2(GND_net), .I3(n43606), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_19 (.CI(n43920), 
            .I0(n3117), .I1(VCC_net), .CO(n43921));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_18_lut (.I0(GND_net), 
            .I1(n3118), .I2(VCC_net), .I3(n43919), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_18 (.CI(n43919), 
            .I0(n3118), .I1(VCC_net), .CO(n43920));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_6 (.CI(n43606), 
            .I0(n1730), .I1(GND_net), .CO(n43607));
    SB_LUT4 add_263_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_359), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_17_lut (.I0(GND_net), 
            .I1(n3119), .I2(VCC_net), .I3(n43918), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_17 (.CI(n43918), 
            .I0(n3119), .I1(VCC_net), .CO(n43919));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_5_lut (.I0(GND_net), 
            .I1(n1731), .I2(VCC_net), .I3(n43605), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_16_lut (.I0(GND_net), 
            .I1(n3120), .I2(VCC_net), .I3(n43917), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_9 (.CI(n43087), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n43088));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_16 (.CI(n43917), 
            .I0(n3120), .I1(VCC_net), .CO(n43918));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_15_lut (.I0(GND_net), 
            .I1(n3121), .I2(VCC_net), .I3(n43916), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_15 (.CI(n43916), 
            .I0(n3121), .I1(VCC_net), .CO(n43917));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_14_lut (.I0(GND_net), 
            .I1(n3122), .I2(VCC_net), .I3(n43915), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_14 (.CI(n43915), 
            .I0(n3122), .I1(VCC_net), .CO(n43916));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_5 (.CI(n43605), 
            .I0(n1731), .I1(VCC_net), .CO(n43606));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_13_lut (.I0(GND_net), 
            .I1(n3123), .I2(VCC_net), .I3(n43914), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_13 (.CI(n43914), 
            .I0(n3123), .I1(VCC_net), .CO(n43915));
    SB_LUT4 add_263_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n43098), .O(encoder1_position_scaled_23__N_75[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_12_lut (.I0(GND_net), 
            .I1(n3124), .I2(VCC_net), .I3(n43913), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_12 (.CI(n43913), 
            .I0(n3124), .I1(VCC_net), .CO(n43914));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_11_lut (.I0(GND_net), 
            .I1(n3125), .I2(VCC_net), .I3(n43912), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_11 (.CI(n43912), 
            .I0(n3125), .I1(VCC_net), .CO(n43913));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_10_lut (.I0(GND_net), 
            .I1(n3126), .I2(VCC_net), .I3(n43911), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_10 (.CI(n43911), 
            .I0(n3126), .I1(VCC_net), .CO(n43912));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_9_lut (.I0(GND_net), 
            .I1(n3127), .I2(VCC_net), .I3(n43910), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_4_lut (.I0(GND_net), 
            .I1(n1732), .I2(GND_net), .I3(n43604), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_4 (.CI(n43604), 
            .I0(n1732), .I1(GND_net), .CO(n43605));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_9 (.CI(n43910), 
            .I0(n3127), .I1(VCC_net), .CO(n43911));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_3_lut (.I0(GND_net), 
            .I1(n1733), .I2(VCC_net), .I3(n43603), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n10832_bdd_4_lut_40548 (.I0(n10832), .I1(n436), .I2(current[5]), 
            .I3(duty[23]), .O(n56344));
    defparam n10832_bdd_4_lut_40548.LUT_INIT = 16'he4aa;
    SB_LUT4 n56344_bdd_4_lut (.I0(n56344), .I1(duty[5]), .I2(n265), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[5]));
    defparam n56344_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_3 (.CI(n43603), 
            .I0(n1733), .I1(VCC_net), .CO(n43604));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1172_3_lut (.I0(n1721), 
            .I1(n1788), .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40543 (.I0(n10832), .I1(n437), .I2(current[4]), 
            .I3(duty[23]), .O(n56338));
    defparam n10832_bdd_4_lut_40543.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_8_lut (.I0(GND_net), 
            .I1(n3128), .I2(VCC_net), .I3(n43909), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_8 (.CI(n43909), 
            .I0(n3128), .I1(VCC_net), .CO(n43910));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1168_2_lut (.I0(GND_net), 
            .I1(n528), .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1168_2 (.CI(VCC_net), 
            .I0(n528), .I1(GND_net), .CO(n43603));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_16_lut (.I0(GND_net), 
            .I1(n1620), .I2(VCC_net), .I3(n43602), .O(n1687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_7_lut (.I0(GND_net), 
            .I1(n3129), .I2(GND_net), .I3(n43908), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_7 (.CI(n43908), 
            .I0(n3129), .I1(GND_net), .CO(n43909));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_6_lut (.I0(GND_net), 
            .I1(n3130), .I2(GND_net), .I3(n43907), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n56338_bdd_4_lut (.I0(n56338), .I1(duty[4]), .I2(n266), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[4]));
    defparam n56338_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_6 (.CI(n43907), 
            .I0(n3130), .I1(GND_net), .CO(n43908));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_5_lut (.I0(GND_net), 
            .I1(n3131), .I2(VCC_net), .I3(n43906), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_5 (.CI(n43906), 
            .I0(n3131), .I1(VCC_net), .CO(n43907));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_4_lut (.I0(GND_net), 
            .I1(n3132), .I2(GND_net), .I3(n43905), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_4 (.CI(n43905), 
            .I0(n3132), .I1(GND_net), .CO(n43906));
    SB_CARRY add_263_20 (.CI(n43098), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n43099));
    SB_LUT4 i21942_2_lut_2_lut (.I0(duty[23]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4906));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21942_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1239_3_lut (.I0(n1820), 
            .I1(n1887), .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n10832_bdd_4_lut_40538 (.I0(n10832), .I1(n438), .I2(current[3]), 
            .I3(duty[23]), .O(n56332));
    defparam n10832_bdd_4_lut_40538.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_3_lut (.I0(GND_net), 
            .I1(n3133), .I2(VCC_net), .I3(n43904), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_3 (.CI(n43904), 
            .I0(n3133), .I1(VCC_net), .CO(n43905));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2106_2_lut (.I0(GND_net), 
            .I1(n542), .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2106_2 (.CI(VCC_net), 
            .I0(n542), .I1(GND_net), .CO(n43904));
    SB_LUT4 n56332_bdd_4_lut (.I0(n56332), .I1(duty[3]), .I2(n267), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[3]));
    defparam n56332_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_30_lut (.I0(GND_net), 
            .I1(n3006), .I2(VCC_net), .I3(n43903), .O(n3073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_29_lut (.I0(GND_net), 
            .I1(n3007), .I2(VCC_net), .I3(n43902), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_29 (.CI(n43902), 
            .I0(n3007), .I1(VCC_net), .CO(n43903));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_15_lut (.I0(GND_net), 
            .I1(n1621), .I2(VCC_net), .I3(n43601), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5618), .I3(n44246), .O(n2_adj_5509)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_28_lut (.I0(GND_net), 
            .I1(n3008), .I2(VCC_net), .I3(n43901), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_15 (.CI(n43601), 
            .I0(n1621), .I1(VCC_net), .CO(n43602));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_28 (.CI(n43901), 
            .I0(n3008), .I1(VCC_net), .CO(n43902));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5619), .I3(n44245), .O(n3_adj_5508)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1306_3_lut (.I0(n1919), 
            .I1(n1986), .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_27_lut (.I0(GND_net), 
            .I1(n3009), .I2(VCC_net), .I3(n43900), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_14_lut (.I0(GND_net), 
            .I1(n1622), .I2(VCC_net), .I3(n43600), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_32 (.CI(n44245), 
            .I0(GND_net), .I1(n3_adj_5619), .CO(n44246));
    SB_LUT4 i21943_2_lut_2_lut (.I0(duty[22]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4907));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21943_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_14 (.CI(n43600), 
            .I0(n1622), .I1(VCC_net), .CO(n43601));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_13_lut (.I0(GND_net), 
            .I1(n1623), .I2(VCC_net), .I3(n43599), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5620), .I3(n44244), .O(n4_adj_5507)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_27 (.CI(n43900), 
            .I0(n3009), .I1(VCC_net), .CO(n43901));
    SB_LUT4 add_261_23_lut (.I0(current[15]), .I1(duty[23]), .I2(n56288), 
            .I3(n43124), .O(n249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_23_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_31 (.CI(n44244), 
            .I0(GND_net), .I1(n4_adj_5620), .CO(n44245));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_26_lut (.I0(GND_net), 
            .I1(n3010), .I2(VCC_net), .I3(n43899), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_13 (.CI(n43599), 
            .I0(n1623), .I1(VCC_net), .CO(n43600));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_26 (.CI(n43899), 
            .I0(n3010), .I1(VCC_net), .CO(n43900));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1373_3_lut (.I0(n2018), 
            .I1(n2085), .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1440_3_lut (.I0(n2117), 
            .I1(n2184), .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_12_lut (.I0(GND_net), 
            .I1(n1624), .I2(VCC_net), .I3(n43598), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_12 (.CI(n43598), 
            .I0(n1624), .I1(VCC_net), .CO(n43599));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_25_lut (.I0(GND_net), 
            .I1(n3011), .I2(VCC_net), .I3(n43898), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_263), 
            .I3(n43210), .O(n356)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5621), .I3(n44243), .O(n5_adj_5506)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_22_lut (.I0(current[15]), .I1(duty[23]), .I2(n56288), 
            .I3(n43123), .O(n250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_22_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_25 (.CI(n43898), 
            .I0(n3011), .I1(VCC_net), .CO(n43899));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_11_lut (.I0(GND_net), 
            .I1(n1625), .I2(VCC_net), .I3(n43597), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_25_lut (.I0(n4748), .I1(GND_net), .I2(pwm_setpoint_23__N_263), 
            .I3(n43209), .O(n4884)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_24_lut (.I0(GND_net), 
            .I1(n3012), .I2(VCC_net), .I3(n43897), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_25 (.CI(n43209), .I0(GND_net), .I1(pwm_setpoint_23__N_263), 
            .CO(n43210));
    SB_LUT4 unary_minus_21_add_3_24_lut (.I0(n4748), .I1(GND_net), .I2(n3), 
            .I3(n43208), .O(n4885)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_261_22 (.CI(n43123), .I0(duty[23]), .I1(n56288), .CO(n43124));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_30 (.CI(n44243), 
            .I0(GND_net), .I1(n5_adj_5621), .CO(n44244));
    SB_CARRY unary_minus_21_add_3_24 (.CI(n43208), .I0(GND_net), .I1(n3), 
            .CO(n43209));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1109_3_lut (.I0(n1626), 
            .I1(n1693), .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1507_3_lut (.I0(n2216), 
            .I1(n2283), .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_24 (.CI(n43897), 
            .I0(n3012), .I1(VCC_net), .CO(n43898));
    SB_LUT4 unary_minus_21_add_3_23_lut (.I0(n4748), .I1(GND_net), .I2(n4_adj_5460), 
            .I3(n43207), .O(n4886)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_23_lut (.I0(GND_net), 
            .I1(n3013), .I2(VCC_net), .I3(n43896), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_23 (.CI(n43896), 
            .I0(n3013), .I1(VCC_net), .CO(n43897));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_11 (.CI(n43597), 
            .I0(n1625), .I1(VCC_net), .CO(n43598));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_10_lut (.I0(GND_net), 
            .I1(n1626), .I2(VCC_net), .I3(n43596), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_23 (.CI(n43207), .I0(GND_net), .I1(n4_adj_5460), 
            .CO(n43208));
    SB_LUT4 add_261_21_lut (.I0(current[15]), .I1(duty[22]), .I2(n56288), 
            .I3(n43122), .O(n251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_21_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 unary_minus_21_add_3_22_lut (.I0(n4748), .I1(GND_net), .I2(n5_adj_5461), 
            .I3(n43206), .O(n4887)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_22 (.CI(n43206), .I0(GND_net), .I1(n5_adj_5461), 
            .CO(n43207));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_22_lut (.I0(GND_net), 
            .I1(n3014), .I2(VCC_net), .I3(n43895), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_22 (.CI(n43895), 
            .I0(n3014), .I1(VCC_net), .CO(n43896));
    SB_CARRY add_261_21 (.CI(n43122), .I0(duty[22]), .I1(n56288), .CO(n43123));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5622), .I3(n44242), .O(n6_adj_5505)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_21_lut (.I0(GND_net), 
            .I1(n3015), .I2(VCC_net), .I3(n43894), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_29 (.CI(n44242), 
            .I0(GND_net), .I1(n6_adj_5622), .CO(n44243));
    SB_LUT4 unary_minus_21_add_3_21_lut (.I0(n4748), .I1(GND_net), .I2(n6), 
            .I3(n43205), .O(n4888)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_21 (.CI(n43205), .I0(GND_net), .I1(n6), 
            .CO(n43206));
    SB_LUT4 n10832_bdd_4_lut_40533 (.I0(n10832), .I1(n439), .I2(current[2]), 
            .I3(duty[23]), .O(n56314));
    defparam n10832_bdd_4_lut_40533.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_21 (.CI(n43894), 
            .I0(n3015), .I1(VCC_net), .CO(n43895));
    SB_LUT4 add_263_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n43097), .O(encoder1_position_scaled_23__N_75[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1574_3_lut (.I0(n2315), 
            .I1(n2382), .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n56314_bdd_4_lut (.I0(n56314), .I1(duty[2]), .I2(n268), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[2]));
    defparam n56314_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1176_3_lut (.I0(n1725), 
            .I1(n1792), .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_261_20_lut (.I0(current[15]), .I1(duty[21]), .I2(n56288), 
            .I3(n43121), .O(n252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_20_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 unary_minus_21_add_3_20_lut (.I0(n4748), .I1(GND_net), .I2(n7), 
            .I3(n43204), .O(n4889)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_261_20 (.CI(n43121), .I0(duty[21]), .I1(n56288), .CO(n43122));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_20_lut (.I0(GND_net), 
            .I1(n3016), .I2(VCC_net), .I3(n43893), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_261_19_lut (.I0(current[15]), .I1(duty[20]), .I2(n56288), 
            .I3(n43120), .O(n253)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_19_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5623), .I3(n44241), .O(n7_adj_5504)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_10 (.CI(n43596), 
            .I0(n1626), .I1(VCC_net), .CO(n43597));
    SB_CARRY add_261_19 (.CI(n43120), .I0(duty[20]), .I1(n56288), .CO(n43121));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_9_lut (.I0(GND_net), 
            .I1(n1627), .I2(VCC_net), .I3(n43595), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_9 (.CI(n43595), 
            .I0(n1627), .I1(VCC_net), .CO(n43596));
    SB_LUT4 add_261_18_lut (.I0(current[15]), .I1(duty[19]), .I2(n56288), 
            .I3(n43119), .O(n254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_18_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_8_lut (.I0(GND_net), 
            .I1(n1628), .I2(VCC_net), .I3(n43594), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_8 (.CI(n43594), 
            .I0(n1628), .I1(VCC_net), .CO(n43595));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_28 (.CI(n44241), 
            .I0(GND_net), .I1(n7_adj_5623), .CO(n44242));
    SB_CARRY unary_minus_21_add_3_20 (.CI(n43204), .I0(GND_net), .I1(n7), 
            .CO(n43205));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5624), .I3(n44240), .O(n8_adj_5503)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_19_lut (.I0(n4748), .I1(GND_net), .I2(n8_adj_5462), 
            .I3(n43203), .O(n4890)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_263_19 (.CI(n43097), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n43098));
    SB_CARRY add_261_18 (.CI(n43119), .I0(duty[19]), .I1(n56288), .CO(n43120));
    SB_LUT4 add_261_17_lut (.I0(current[15]), .I1(duty[18]), .I2(n56288), 
            .I3(n43118), .O(n255)) /* synthesis syn_instantiated=1 */ ;
    defparam add_261_17_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_20 (.CI(n43893), 
            .I0(n3016), .I1(VCC_net), .CO(n43894));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_19_lut (.I0(GND_net), 
            .I1(n3017), .I2(VCC_net), .I3(n43892), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_19 (.CI(n43203), .I0(GND_net), .I1(n8_adj_5462), 
            .CO(n43204));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i27_3_lut (.I0(encoder0_position_scaled_23__N_327[26]), 
            .I1(n7_adj_5504), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_19 (.CI(n43892), 
            .I0(n3017), .I1(VCC_net), .CO(n43893));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_18_lut (.I0(GND_net), 
            .I1(n3018), .I2(VCC_net), .I3(n43891), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_7_lut (.I0(GND_net), 
            .I1(n1629), .I2(GND_net), .I3(n43593), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_18_lut (.I0(n4748), .I1(GND_net), .I2(n9), 
            .I3(n43202), .O(n4891)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_7 (.CI(n43593), 
            .I0(n1629), .I1(GND_net), .CO(n43594));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_6_lut (.I0(GND_net), 
            .I1(n1630), .I2(GND_net), .I3(n43592), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_6 (.CI(n43592), 
            .I0(n1630), .I1(GND_net), .CO(n43593));
    SB_CARRY unary_minus_21_add_3_18 (.CI(n43202), .I0(GND_net), .I1(n9), 
            .CO(n43203));
    SB_LUT4 unary_minus_21_add_3_17_lut (.I0(n4748), .I1(GND_net), .I2(n10), 
            .I3(n43201), .O(n4892)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_27 (.CI(n44240), 
            .I0(GND_net), .I1(n8_adj_5624), .CO(n44241));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5625), .I3(n44239), .O(n9_adj_5502)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_26 (.CI(n44239), 
            .I0(GND_net), .I1(n9_adj_5625), .CO(n44240));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_18 (.CI(n43891), 
            .I0(n3018), .I1(VCC_net), .CO(n43892));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_17_lut (.I0(GND_net), 
            .I1(n3019), .I2(VCC_net), .I3(n43890), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_17 (.CI(n43890), 
            .I0(n3019), .I1(VCC_net), .CO(n43891));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5626), .I3(n44238), .O(n10_adj_5501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_17 (.CI(n43201), .I0(GND_net), .I1(n10), 
            .CO(n43202));
    SB_CARRY add_261_17 (.CI(n43118), .I0(duty[18]), .I1(n56288), .CO(n43119));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_16_lut (.I0(GND_net), 
            .I1(n3020), .I2(VCC_net), .I3(n43889), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_16 (.CI(n43889), 
            .I0(n3020), .I1(VCC_net), .CO(n43890));
    SB_LUT4 add_263_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n43086), .O(encoder1_position_scaled_23__N_75[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_15_lut (.I0(GND_net), 
            .I1(n3021), .I2(VCC_net), .I3(n43888), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_15 (.CI(n43888), 
            .I0(n3021), .I1(VCC_net), .CO(n43889));
    SB_LUT4 unary_minus_21_add_3_16_lut (.I0(n4748), .I1(GND_net), .I2(n11), 
            .I3(n43200), .O(n4893)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_263_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n43096), .O(encoder1_position_scaled_23__N_75[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_14_lut (.I0(GND_net), 
            .I1(n3022), .I2(VCC_net), .I3(n43887), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_18 (.CI(n43096), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n43097));
    SB_CARRY add_263_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_359), 
            .CO(n43081));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_14 (.CI(n43887), 
            .I0(n3022), .I1(VCC_net), .CO(n43888));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_25 (.CI(n44238), 
            .I0(GND_net), .I1(n10_adj_5626), .CO(n44239));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5627), .I3(n44237), .O(n11_adj_5500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n10832_bdd_4_lut_40519 (.I0(n10832), .I1(n440), .I2(current[1]), 
            .I3(duty[23]), .O(n56308));
    defparam n10832_bdd_4_lut_40519.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_24 (.CI(n44237), 
            .I0(GND_net), .I1(n11_adj_5627), .CO(n44238));
    SB_CARRY unary_minus_21_add_3_16 (.CI(n43200), .I0(GND_net), .I1(n11), 
            .CO(n43201));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5628), .I3(n44236), .O(n12_adj_5499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_23 (.CI(n44236), 
            .I0(GND_net), .I1(n12_adj_5628), .CO(n44237));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_5_lut (.I0(GND_net), 
            .I1(n1631), .I2(VCC_net), .I3(n43591), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_13_lut (.I0(GND_net), 
            .I1(n3023), .I2(VCC_net), .I3(n43886), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_13 (.CI(n43886), 
            .I0(n3023), .I1(VCC_net), .CO(n43887));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_12_lut (.I0(GND_net), 
            .I1(n3024), .I2(VCC_net), .I3(n43885), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5629), .I3(n44235), .O(n13_adj_5498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_8 (.CI(n43086), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n43087));
    SB_LUT4 n56308_bdd_4_lut (.I0(n56308), .I1(duty[1]), .I2(n269), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[1]));
    defparam n56308_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_5 (.CI(n43591), 
            .I0(n1631), .I1(VCC_net), .CO(n43592));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_22 (.CI(n44235), 
            .I0(GND_net), .I1(n13_adj_5629), .CO(n44236));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_12 (.CI(n43885), 
            .I0(n3024), .I1(VCC_net), .CO(n43886));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_11_lut (.I0(GND_net), 
            .I1(n3025), .I2(VCC_net), .I3(n43884), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_4_lut (.I0(GND_net), 
            .I1(n1632), .I2(GND_net), .I3(n43590), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_11 (.CI(n43884), 
            .I0(n3025), .I1(VCC_net), .CO(n43885));
    SB_LUT4 i21944_2_lut_2_lut (.I0(duty[21]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4908));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21944_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_10_lut (.I0(GND_net), 
            .I1(n3026), .I2(VCC_net), .I3(n43883), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5630), .I3(n44234), .O(n14_adj_5497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_10 (.CI(n43883), 
            .I0(n3026), .I1(VCC_net), .CO(n43884));
    SB_LUT4 i1_4_lut_adj_1875 (.I0(n4_adj_5507), .I1(n5_adj_5506), .I2(n518), 
            .I3(n6_adj_5505), .O(n5_adj_5482));
    defparam i1_4_lut_adj_1875.LUT_INIT = 16'heeea;
    SB_LUT4 unary_minus_21_add_3_15_lut (.I0(n4748), .I1(GND_net), .I2(n12), 
            .I3(n43199), .O(n4894)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_4 (.CI(n43590), 
            .I0(n1632), .I1(GND_net), .CO(n43591));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_21 (.CI(n44234), 
            .I0(GND_net), .I1(n14_adj_5630), .CO(n44235));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_9_lut (.I0(GND_net), 
            .I1(n3027), .I2(VCC_net), .I3(n43882), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_15 (.CI(n43199), .I0(GND_net), .I1(n12), 
            .CO(n43200));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_9 (.CI(n43882), 
            .I0(n3027), .I1(VCC_net), .CO(n43883));
    SB_LUT4 i21945_2_lut_2_lut (.I0(duty[20]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4909));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21945_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_8_lut (.I0(GND_net), 
            .I1(n3028), .I2(VCC_net), .I3(n43881), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_8 (.CI(n43881), 
            .I0(n3028), .I1(VCC_net), .CO(n43882));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5631), .I3(n44233), .O(n15_adj_5496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_3_lut (.I0(GND_net), 
            .I1(n1633), .I2(VCC_net), .I3(n43589), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_3 (.CI(n43589), 
            .I0(n1633), .I1(VCC_net), .CO(n43590));
    SB_LUT4 i21946_2_lut_2_lut (.I0(duty[19]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4910));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21946_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1101_2_lut (.I0(GND_net), 
            .I1(n527), .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_7_lut (.I0(GND_net), 
            .I1(n3029), .I2(GND_net), .I3(n43880), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1101_2 (.CI(VCC_net), 
            .I0(n527), .I1(GND_net), .CO(n43589));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_7 (.CI(n43880), 
            .I0(n3029), .I1(GND_net), .CO(n43881));
    SB_LUT4 unary_minus_21_add_3_14_lut (.I0(n4748), .I1(GND_net), .I2(n13), 
            .I3(n43198), .O(n4895)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i21947_2_lut_2_lut (.I0(duty[18]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4911));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21947_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY unary_minus_21_add_3_14 (.CI(n43198), .I0(GND_net), .I1(n13), 
            .CO(n43199));
    SB_DFFESR GLC_215 (.Q(INLC_c_0), .C(clk16MHz), .E(n28583), .D(GLC_N_523), 
            .R(n29049));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i15344_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_5478), 
            .I3(n27232), .O(n29420));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15344_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_263_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n43085), .O(encoder1_position_scaled_23__N_75[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_20 (.CI(n44233), 
            .I0(GND_net), .I1(n15_adj_5631), .CO(n44234));
    SB_LUT4 i38617_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5605), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[0]), .O(n54290));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38617_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 add_263_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n43095), .O(encoder1_position_scaled_23__N_75[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5632), .I3(n44232), .O(n16_adj_5495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_19 (.CI(n44232), 
            .I0(GND_net), .I1(n16_adj_5632), .CO(n44233));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_6_lut (.I0(GND_net), 
            .I1(n3030), .I2(GND_net), .I3(n43879), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_6 (.CI(n43879), 
            .I0(n3030), .I1(GND_net), .CO(n43880));
    SB_LUT4 unary_minus_21_add_3_13_lut (.I0(n4748), .I1(GND_net), .I2(n14), 
            .I3(n43197), .O(n4896)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_15_lut (.I0(n56120), 
            .I1(n1521), .I2(VCC_net), .I3(n43588), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5633), .I3(n44231), .O(n17_adj_5494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_5_lut (.I0(GND_net), 
            .I1(n3031), .I2(VCC_net), .I3(n43878), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_5 (.CI(n43878), 
            .I0(n3031), .I1(VCC_net), .CO(n43879));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_4_lut (.I0(GND_net), 
            .I1(n3032), .I2(GND_net), .I3(n43877), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_14_lut (.I0(GND_net), 
            .I1(n1522), .I2(VCC_net), .I3(n43587), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_13 (.CI(n43197), .I0(GND_net), .I1(n14), 
            .CO(n43198));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_14 (.CI(n43587), 
            .I0(n1522), .I1(VCC_net), .CO(n43588));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_4 (.CI(n43877), 
            .I0(n3032), .I1(GND_net), .CO(n43878));
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(n4748), .I1(GND_net), .I2(n15_adj_5463), 
            .I3(n43196), .O(n4897)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_12 (.CI(n43196), .I0(GND_net), .I1(n15_adj_5463), 
            .CO(n43197));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_18 (.CI(n44231), 
            .I0(GND_net), .I1(n17_adj_5633), .CO(n44232));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_13_lut (.I0(GND_net), 
            .I1(n1523), .I2(VCC_net), .I3(n43586), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5634), .I3(n44230), .O(n18_adj_5493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(n4748), .I1(GND_net), .I2(n16), 
            .I3(n43195), .O(n4898)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_17 (.CI(n44230), 
            .I0(GND_net), .I1(n18_adj_5634), .CO(n44231));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_3_lut (.I0(GND_net), 
            .I1(n3033), .I2(VCC_net), .I3(n43876), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_3 (.CI(n43876), 
            .I0(n3033), .I1(VCC_net), .CO(n43877));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_2039_2_lut (.I0(GND_net), 
            .I1(n541), .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_13 (.CI(n43586), 
            .I0(n1523), .I1(VCC_net), .CO(n43587));
    SB_CARRY add_263_17 (.CI(n43095), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n43096));
    SB_LUT4 add_263_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n43094), .O(encoder1_position_scaled_23__N_75[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1243_3_lut (.I0(n1824), 
            .I1(n1891), .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_2039_2 (.CI(VCC_net), 
            .I0(n541), .I1(GND_net), .CO(n43876));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_29_lut (.I0(n55788), 
            .I1(n2907), .I2(VCC_net), .I3(n43875), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_28_lut (.I0(GND_net), 
            .I1(n2908), .I2(VCC_net), .I3(n43874), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38593_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5605), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[1]), .O(n54253));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38593_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5635), .I3(n44229), .O(n19_adj_5492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_28 (.CI(n43874), 
            .I0(n2908), .I1(VCC_net), .CO(n43875));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_27_lut (.I0(GND_net), 
            .I1(n2909), .I2(VCC_net), .I3(n43873), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_16 (.CI(n44229), 
            .I0(GND_net), .I1(n19_adj_5635), .CO(n44230));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_27 (.CI(n43873), 
            .I0(n2909), .I1(VCC_net), .CO(n43874));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_26_lut (.I0(GND_net), 
            .I1(n2910), .I2(VCC_net), .I3(n43872), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5636), .I3(n44228), .O(n20_adj_5491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_26 (.CI(n43872), 
            .I0(n2910), .I1(VCC_net), .CO(n43873));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_25_lut (.I0(GND_net), 
            .I1(n2911), .I2(VCC_net), .I3(n43871), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38680_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5605), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[2]), .O(n54252));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38680_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_15 (.CI(n44228), 
            .I0(GND_net), .I1(n20_adj_5636), .CO(n44229));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_25 (.CI(n43871), 
            .I0(n2911), .I1(VCC_net), .CO(n43872));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_24_lut (.I0(GND_net), 
            .I1(n2912), .I2(VCC_net), .I3(n43870), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5637), .I3(n44227), .O(n21_adj_5490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_24 (.CI(n43870), 
            .I0(n2912), .I1(VCC_net), .CO(n43871));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_23_lut (.I0(GND_net), 
            .I1(n2913), .I2(VCC_net), .I3(n43869), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_14 (.CI(n44227), 
            .I0(GND_net), .I1(n21_adj_5637), .CO(n44228));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_23 (.CI(n43869), 
            .I0(n2913), .I1(VCC_net), .CO(n43870));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_12_lut (.I0(GND_net), 
            .I1(n1524), .I2(VCC_net), .I3(n43585), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_12 (.CI(n43585), 
            .I0(n1524), .I1(VCC_net), .CO(n43586));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5638), .I3(n44226), .O(n22_adj_5489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_11_lut (.I0(GND_net), 
            .I1(n1525), .I2(VCC_net), .I3(n43584), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_22_lut (.I0(GND_net), 
            .I1(n2914), .I2(VCC_net), .I3(n43868), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_22 (.CI(n43868), 
            .I0(n2914), .I1(VCC_net), .CO(n43869));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_21_lut (.I0(GND_net), 
            .I1(n2915), .I2(VCC_net), .I3(n43867), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_13 (.CI(n44226), 
            .I0(GND_net), .I1(n22_adj_5638), .CO(n44227));
    SB_CARRY unary_minus_21_add_3_11 (.CI(n43195), .I0(GND_net), .I1(n16), 
            .CO(n43196));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_21 (.CI(n43867), 
            .I0(n2915), .I1(VCC_net), .CO(n43868));
    SB_CARRY add_263_7 (.CI(n43085), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n43086));
    SB_LUT4 i38678_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5605), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[3]), .O(n54251));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38678_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_20_lut (.I0(GND_net), 
            .I1(n2916), .I2(VCC_net), .I3(n43866), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_20 (.CI(n43866), 
            .I0(n2916), .I1(VCC_net), .CO(n43867));
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(n4748), .I1(GND_net), .I2(n17), 
            .I3(n43194), .O(n4899)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_19_lut (.I0(GND_net), 
            .I1(n2917), .I2(VCC_net), .I3(n43865), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38677_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5605), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[4]), .O(n54250));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38677_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5639), .I3(n44225), .O(n23_adj_5488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_19 (.CI(n43865), 
            .I0(n2917), .I1(VCC_net), .CO(n43866));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_18_lut (.I0(GND_net), 
            .I1(n2918), .I2(VCC_net), .I3(n43864), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_12 (.CI(n44225), 
            .I0(GND_net), .I1(n23_adj_5639), .CO(n44226));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5640), .I3(n44224), .O(n24_adj_5487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_16 (.CI(n43094), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n43095));
    SB_CARRY unary_minus_21_add_3_10 (.CI(n43194), .I0(GND_net), .I1(n17), 
            .CO(n43195));
    SB_LUT4 i21948_2_lut_2_lut (.I0(duty[17]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4912));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21948_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_11 (.CI(n44224), 
            .I0(GND_net), .I1(n24_adj_5640), .CO(n44225));
    SB_LUT4 i15360_4_lut_4_lut (.I0(n28689), .I1(state[0]), .I2(state[1]), 
            .I3(state_3__N_639[1]), .O(n29436));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15360_4_lut_4_lut.LUT_INIT = 16'hfa7a;
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
           .D(n48472));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i38676_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5605), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[5]), .O(n54249));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38676_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5641), .I3(n44223), .O(n25_adj_5486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_18 (.CI(n43864), 
            .I0(n2918), .I1(VCC_net), .CO(n43865));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_17_lut (.I0(GND_net), 
            .I1(n2919), .I2(VCC_net), .I3(n43863), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38630_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5605), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[6]), .O(n54248));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38630_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 n10832_bdd_4_lut_40514 (.I0(n10832), .I1(n441), .I2(current[0]), 
            .I3(duty[23]), .O(n56302));
    defparam n10832_bdd_4_lut_40514.LUT_INIT = 16'he4aa;
    SB_LUT4 add_263_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n43084), .O(encoder1_position_scaled_23__N_75[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(n4748), .I1(GND_net), .I2(n18), 
            .I3(n43193), .O(n4900)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_17 (.CI(n43863), 
            .I0(n2919), .I1(VCC_net), .CO(n43864));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_16_lut (.I0(GND_net), 
            .I1(n2920), .I2(VCC_net), .I3(n43862), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38589_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5605), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[7]), .O(n54247));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i38589_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i21949_2_lut_2_lut (.I0(duty[16]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n4913));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21949_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY unary_minus_21_add_3_9 (.CI(n43193), .I0(GND_net), .I1(n18), 
            .CO(n43194));
    SB_LUT4 i1_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5605), 
            .I2(commutation_state_prev[0]), .I3(dti_N_527), .O(n28559));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i2_2_lut_3_lut (.I0(hall1), .I1(hall3), .I2(hall2), .I3(GND_net), 
            .O(commutation_state_7__N_272));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n49501));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i33742_3_lut (.I0(n3_adj_5508), .I1(n8585), .I2(n49468), .I3(GND_net), 
            .O(n49469));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33742_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(clk16MHz), .D(n29714));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(clk16MHz), .D(n29713));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(clk16MHz), .D(n29712));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(clk16MHz), .D(n29711));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(clk16MHz), .D(n29710));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(clk16MHz), .D(n29709));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(clk16MHz), .D(n29708));   // verilog/TinyFPGA_B.v(368[10] 396[6])
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_10 (.CI(n44223), 
            .I0(GND_net), .I1(n25_adj_5641), .CO(n44224));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_16 (.CI(n43862), 
            .I0(n2920), .I1(VCC_net), .CO(n43863));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_15_lut (.I0(GND_net), 
            .I1(n2921), .I2(VCC_net), .I3(n43861), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5642), .I3(n44222), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_15 (.CI(n43861), 
            .I0(n2921), .I1(VCC_net), .CO(n43862));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_14_lut (.I0(GND_net), 
            .I1(n2922), .I2(VCC_net), .I3(n43860), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_9 (.CI(n44222), 
            .I0(GND_net), .I1(n26_adj_5642), .CO(n44223));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_14 (.CI(n43860), 
            .I0(n2922), .I1(VCC_net), .CO(n43861));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_13_lut (.I0(GND_net), 
            .I1(n2923), .I2(VCC_net), .I3(n43859), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5643), .I3(n44221), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_13 (.CI(n43859), 
            .I0(n2923), .I1(VCC_net), .CO(n43860));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_12_lut (.I0(GND_net), 
            .I1(n2924), .I2(VCC_net), .I3(n43858), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_8 (.CI(n44221), 
            .I0(GND_net), .I1(n27_adj_5643), .CO(n44222));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_12 (.CI(n43858), 
            .I0(n2924), .I1(VCC_net), .CO(n43859));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_11_lut (.I0(GND_net), 
            .I1(n2925), .I2(VCC_net), .I3(n43857), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5644), .I3(n44220), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_11 (.CI(n43857), 
            .I0(n2925), .I1(VCC_net), .CO(n43858));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_10_lut (.I0(GND_net), 
            .I1(n2926), .I2(VCC_net), .I3(n43856), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_7 (.CI(n44220), 
            .I0(GND_net), .I1(n28_adj_5644), .CO(n44221));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_10 (.CI(n43856), 
            .I0(n2926), .I1(VCC_net), .CO(n43857));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_9_lut (.I0(GND_net), 
            .I1(n2927), .I2(VCC_net), .I3(n43855), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5645), .I3(n44219), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_9 (.CI(n43855), 
            .I0(n2927), .I1(VCC_net), .CO(n43856));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_8_lut (.I0(GND_net), 
            .I1(n2928), .I2(VCC_net), .I3(n43854), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_6 (.CI(n44219), 
            .I0(GND_net), .I1(n29_adj_5645), .CO(n44220));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_8 (.CI(n43854), 
            .I0(n2928), .I1(VCC_net), .CO(n43855));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_7_lut (.I0(GND_net), 
            .I1(n2929), .I2(GND_net), .I3(n43853), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5646), .I3(n44218), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_7 (.CI(n43853), 
            .I0(n2929), .I1(GND_net), .CO(n43854));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_6_lut (.I0(GND_net), 
            .I1(n2930), .I2(GND_net), .I3(n43852), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_5 (.CI(n44218), 
            .I0(GND_net), .I1(n30_adj_5646), .CO(n44219));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_6 (.CI(n43852), 
            .I0(n2930), .I1(GND_net), .CO(n43853));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_5_lut (.I0(GND_net), 
            .I1(n2931), .I2(VCC_net), .I3(n43851), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5647), .I3(n44217), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_5 (.CI(n43851), 
            .I0(n2931), .I1(VCC_net), .CO(n43852));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_4_lut (.I0(GND_net), 
            .I1(n2932), .I2(GND_net), .I3(n43850), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_4 (.CI(n44217), 
            .I0(GND_net), .I1(n31_adj_5647), .CO(n44218));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_4 (.CI(n43850), 
            .I0(n2932), .I1(GND_net), .CO(n43851));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_3_lut (.I0(GND_net), 
            .I1(n2933), .I2(VCC_net), .I3(n43849), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5648), .I3(n44216), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_3 (.CI(n43849), 
            .I0(n2933), .I1(VCC_net), .CO(n43850));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1972_2_lut (.I0(GND_net), 
            .I1(n540), .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_3 (.CI(n44216), 
            .I0(GND_net), .I1(n32_adj_5648), .CO(n44217));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1972_2 (.CI(VCC_net), 
            .I0(n540), .I1(GND_net), .CO(n43849));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_28_lut (.I0(n55819), 
            .I1(n2808), .I2(VCC_net), .I3(n43848), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5649), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_27_lut (.I0(GND_net), 
            .I1(n2809), .I2(VCC_net), .I3(n43847), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_27 (.CI(n43847), 
            .I0(n2809), .I1(VCC_net), .CO(n43848));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_11 (.CI(n43584), 
            .I0(n1525), .I1(VCC_net), .CO(n43585));
    SB_CARRY encoder0_position_scaled_23__I_0_227_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5649), .CO(n44216));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_10_lut (.I0(GND_net), 
            .I1(n1526), .I2(VCC_net), .I3(n43583), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_26_lut (.I0(GND_net), 
            .I1(n2810), .I2(VCC_net), .I3(n43846), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_26 (.CI(n43846), 
            .I0(n2810), .I1(VCC_net), .CO(n43847));
    SB_LUT4 i38925_2_lut_4_lut (.I0(duty[8]), .I1(n338), .I2(duty[4]), 
            .I3(n342), .O(n54718));
    defparam i38925_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(n4748), .I1(GND_net), .I2(n19), 
            .I3(n43192), .O(n4901)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_25_lut (.I0(GND_net), 
            .I1(n2811), .I2(VCC_net), .I3(n43845), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_25 (.CI(n43845), 
            .I0(n2811), .I1(VCC_net), .CO(n43846));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_10 (.CI(n43583), 
            .I0(n1526), .I1(VCC_net), .CO(n43584));
    SB_CARRY unary_minus_21_add_3_8 (.CI(n43192), .I0(GND_net), .I1(n19), 
            .CO(n43193));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_24_lut (.I0(GND_net), 
            .I1(n2812), .I2(VCC_net), .I3(n43844), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(n4748), .I1(GND_net), .I2(n20_adj_5464), 
            .I3(n43191), .O(n4902)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_24 (.CI(n43844), 
            .I0(n2812), .I1(VCC_net), .CO(n43845));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_23_lut (.I0(GND_net), 
            .I1(n2813), .I2(VCC_net), .I3(n43843), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_9_lut (.I0(GND_net), 
            .I1(n1527), .I2(VCC_net), .I3(n43582), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_9 (.CI(n43582), 
            .I0(n1527), .I1(VCC_net), .CO(n43583));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_8_lut (.I0(GND_net), 
            .I1(n1528), .I2(VCC_net), .I3(n43581), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_23 (.CI(n43843), 
            .I0(n2813), .I1(VCC_net), .CO(n43844));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_8 (.CI(n43581), 
            .I0(n1528), .I1(VCC_net), .CO(n43582));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_22_lut (.I0(GND_net), 
            .I1(n2814), .I2(VCC_net), .I3(n43842), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_22 (.CI(n43842), 
            .I0(n2814), .I1(VCC_net), .CO(n43843));
    SB_LUT4 add_263_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n43093), .O(encoder1_position_scaled_23__N_75[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_15 (.CI(n43093), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n43094));
    SB_CARRY add_263_6 (.CI(n43084), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n43085));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_7_lut (.I0(GND_net), 
            .I1(n1529), .I2(GND_net), .I3(n43580), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_21_lut (.I0(GND_net), 
            .I1(n2815), .I2(VCC_net), .I3(n43841), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_7 (.CI(n43580), 
            .I0(n1529), .I1(GND_net), .CO(n43581));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_6_lut (.I0(GND_net), 
            .I1(n1530), .I2(GND_net), .I3(n43579), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_6 (.CI(n43579), 
            .I0(n1530), .I1(GND_net), .CO(n43580));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_21 (.CI(n43841), 
            .I0(n2815), .I1(VCC_net), .CO(n43842));
    SB_CARRY unary_minus_21_add_3_7 (.CI(n43191), .I0(GND_net), .I1(n20_adj_5464), 
            .CO(n43192));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_5_lut (.I0(GND_net), 
            .I1(n1531), .I2(VCC_net), .I3(n43578), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_20_lut (.I0(GND_net), 
            .I1(n2816), .I2(VCC_net), .I3(n43840), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_263_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n43092), .O(encoder1_position_scaled_23__N_75[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_263_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_20 (.CI(n43840), 
            .I0(n2816), .I1(VCC_net), .CO(n43841));
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(n4748), .I1(GND_net), .I2(n21), 
            .I3(n43190), .O(n4903)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_19_lut (.I0(GND_net), 
            .I1(n2817), .I2(VCC_net), .I3(n43839), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_5 (.CI(n43578), 
            .I0(n1531), .I1(VCC_net), .CO(n43579));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_4_lut (.I0(GND_net), 
            .I1(n1532_adj_5608), .I2(GND_net), .I3(n43577), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_19 (.CI(n43839), 
            .I0(n2817), .I1(VCC_net), .CO(n43840));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_18_lut (.I0(GND_net), 
            .I1(n2818), .I2(VCC_net), .I3(n43838), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_18 (.CI(n43838), 
            .I0(n2818), .I1(VCC_net), .CO(n43839));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_4 (.CI(n43577), 
            .I0(n1532_adj_5608), .I1(GND_net), .CO(n43578));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_3_lut (.I0(GND_net), 
            .I1(n1533_adj_5609), .I2(VCC_net), .I3(n43576), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_17_lut (.I0(GND_net), 
            .I1(n2819), .I2(VCC_net), .I3(n43837), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_17 (.CI(n43837), 
            .I0(n2819), .I1(VCC_net), .CO(n43838));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_3 (.CI(n43576), 
            .I0(n1533_adj_5609), .I1(VCC_net), .CO(n43577));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1034_2_lut (.I0(GND_net), 
            .I1(n526), .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_6 (.CI(n43190), .I0(GND_net), .I1(n21), 
            .CO(n43191));
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(n296), .I1(GND_net), .I2(n22), 
            .I3(n43189), .O(n4904)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY unary_minus_21_add_3_5 (.CI(n43189), .I0(GND_net), .I1(n22), 
            .CO(n43190));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_16_lut (.I0(GND_net), 
            .I1(n2820), .I2(VCC_net), .I3(n43836), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21964_2_lut (.I0(duty[1]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4928));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21964_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5582));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_16 (.CI(n43836), 
            .I0(n2820), .I1(VCC_net), .CO(n43837));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_15_lut (.I0(GND_net), 
            .I1(n2821), .I2(VCC_net), .I3(n43835), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(n379), .I1(GND_net), .I2(n23), 
            .I3(n43188), .O(n4_adj_5480)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1034_2 (.CI(VCC_net), 
            .I0(n526), .I1(GND_net), .CO(n43576));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_15 (.CI(n43835), 
            .I0(n2821), .I1(VCC_net), .CO(n43836));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_14_lut (.I0(n56150), 
            .I1(n1422), .I2(VCC_net), .I3(n43575), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_14_lut (.I0(GND_net), 
            .I1(n2822), .I2(VCC_net), .I3(n43834), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_13_lut (.I0(GND_net), 
            .I1(n1423), .I2(VCC_net), .I3(n43574), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_263_14 (.CI(n43092), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n43093));
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5583));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_14 (.CI(n43834), 
            .I0(n2822), .I1(VCC_net), .CO(n43835));
    SB_CARRY unary_minus_21_add_3_4 (.CI(n43188), .I0(GND_net), .I1(n23), 
            .CO(n43189));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_13_lut (.I0(GND_net), 
            .I1(n2823), .I2(VCC_net), .I3(n43833), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5465), 
            .I3(n43187), .O(n379)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5579));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5587));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5580_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_478));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5580_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_13 (.CI(n43833), 
            .I0(n2823), .I1(VCC_net), .CO(n43834));
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5584));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5585));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_12_lut (.I0(GND_net), 
            .I1(n2824), .I2(VCC_net), .I3(n43832), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_13 (.CI(n43574), 
            .I0(n1423), .I1(VCC_net), .CO(n43575));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_12 (.CI(n43832), 
            .I0(n2824), .I1(VCC_net), .CO(n43833));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_12_lut (.I0(GND_net), 
            .I1(n1424), .I2(VCC_net), .I3(n43573), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_12 (.CI(n43573), 
            .I0(n1424), .I1(VCC_net), .CO(n43574));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_11_lut (.I0(GND_net), 
            .I1(n1425), .I2(VCC_net), .I3(n43572), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_3 (.CI(n43187), .I0(GND_net), .I1(n24_adj_5465), 
            .CO(n43188));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_11_lut (.I0(GND_net), 
            .I1(n2825), .I2(VCC_net), .I3(n43831), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_11 (.CI(n43831), 
            .I0(n2825), .I1(VCC_net), .CO(n43832));
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(n4_adj_5480), .I1(GND_net), 
            .I2(n25), .I3(VCC_net), .O(n54231)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_10_lut (.I0(GND_net), 
            .I1(n2826), .I2(VCC_net), .I3(n43830), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_11 (.CI(n43572), 
            .I0(n1425), .I1(VCC_net), .CO(n43573));
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5580));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_1039_25_lut (.I0(GND_net), .I1(n4883), .I2(n4906), .I3(n43340), 
            .O(n418)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n43187));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_10 (.CI(n43830), 
            .I0(n2826), .I1(VCC_net), .CO(n43831));
    SB_LUT4 add_1039_24_lut (.I0(GND_net), .I1(n4883), .I2(n4907), .I3(n43339), 
            .O(n419)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i5_2_lut (.I0(current[2]), .I1(duty[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5589));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38899_4_lut (.I0(n11_adj_5584), .I1(n9_adj_5585), .I2(n7_adj_5587), 
            .I3(n5_adj_5589), .O(n54692));
    defparam i38899_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_9_lut (.I0(GND_net), 
            .I1(n2827), .I2(VCC_net), .I3(n43829), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_9 (.CI(n43829), 
            .I0(n2827), .I1(VCC_net), .CO(n43830));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_8_lut (.I0(GND_net), 
            .I1(n2828), .I2(VCC_net), .I3(n43828), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_10_lut (.I0(GND_net), 
            .I1(n1426), .I2(VCC_net), .I3(n43571), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_10 (.CI(n43571), 
            .I0(n1426), .I1(VCC_net), .CO(n43572));
    SB_CARRY add_1039_24 (.CI(n43339), .I0(n4883), .I1(n4907), .CO(n43340));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_9_lut (.I0(GND_net), 
            .I1(n1427), .I2(VCC_net), .I3(n43570), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_9 (.CI(n43570), 
            .I0(n1427), .I1(VCC_net), .CO(n43571));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_8_lut (.I0(GND_net), 
            .I1(n1428), .I2(VCC_net), .I3(n43569), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_8 (.CI(n43569), 
            .I0(n1428), .I1(VCC_net), .CO(n43570));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_8 (.CI(n43828), 
            .I0(n2828), .I1(VCC_net), .CO(n43829));
    SB_LUT4 add_175_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n43186), .O(n1532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_7_lut (.I0(GND_net), 
            .I1(n2829), .I2(GND_net), .I3(n43827), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_7 (.CI(n43827), 
            .I0(n2829), .I1(GND_net), .CO(n43828));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_6_lut (.I0(GND_net), 
            .I1(n2830), .I2(GND_net), .I3(n43826), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_6 (.CI(n43826), 
            .I0(n2830), .I1(GND_net), .CO(n43827));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_5_lut (.I0(GND_net), 
            .I1(n2831), .I2(VCC_net), .I3(n43825), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_5 (.CI(n43825), 
            .I0(n2831), .I1(VCC_net), .CO(n43826));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_4_lut (.I0(GND_net), 
            .I1(n2832), .I2(GND_net), .I3(n43824), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_7_lut (.I0(GND_net), 
            .I1(n1429), .I2(GND_net), .I3(n43568), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_4 (.CI(n43824), 
            .I0(n2832), .I1(GND_net), .CO(n43825));
    SB_LUT4 add_1039_23_lut (.I0(GND_net), .I1(n4883), .I2(n4908), .I3(n43338), 
            .O(n420)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_23 (.CI(n43338), .I0(n4883), .I1(n4908), .CO(n43339));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_3_lut (.I0(GND_net), 
            .I1(n2833), .I2(VCC_net), .I3(n43823), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_3 (.CI(n43823), 
            .I0(n2833), .I1(VCC_net), .CO(n43824));
    SB_LUT4 add_1039_22_lut (.I0(GND_net), .I1(n4884), .I2(n4909), .I3(n43337), 
            .O(n421)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_22 (.CI(n43337), .I0(n4884), .I1(n4909), .CO(n43338));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1905_2_lut (.I0(GND_net), 
            .I1(n539), .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_21_lut (.I0(GND_net), .I1(n4885), .I2(n4910), .I3(n43336), 
            .O(n422)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_175_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n43185), .O(n1533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1905_2 (.CI(VCC_net), 
            .I0(n539), .I1(GND_net), .CO(n43823));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_27_lut (.I0(n55850), 
            .I1(n2709), .I2(VCC_net), .I3(n43822), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_26_lut (.I0(GND_net), 
            .I1(n2710), .I2(VCC_net), .I3(n43821), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_21 (.CI(n43336), .I0(n4885), .I1(n4910), .CO(n43337));
    SB_LUT4 add_1039_20_lut (.I0(GND_net), .I1(n4886), .I2(n4911), .I3(n43335), 
            .O(n423)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_175_32 (.CI(n43185), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n43186));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_26 (.CI(n43821), 
            .I0(n2710), .I1(VCC_net), .CO(n43822));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_7 (.CI(n43568), 
            .I0(n1429), .I1(GND_net), .CO(n43569));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_25_lut (.I0(GND_net), 
            .I1(n2711), .I2(VCC_net), .I3(n43820), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_25 (.CI(n43820), 
            .I0(n2711), .I1(VCC_net), .CO(n43821));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_24_lut (.I0(GND_net), 
            .I1(n2712), .I2(VCC_net), .I3(n43819), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_24 (.CI(n43819), 
            .I0(n2712), .I1(VCC_net), .CO(n43820));
    SB_CARRY add_1039_20 (.CI(n43335), .I0(n4886), .I1(n4911), .CO(n43336));
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_11[0]));   // verilog/TinyFPGA_B.v(103[9] 129[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_6_lut (.I0(GND_net), 
            .I1(n1430), .I2(GND_net), .I3(n43567), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1039_19_lut (.I0(GND_net), .I1(n4887), .I2(n4912), .I3(n43334), 
            .O(n424)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_19 (.CI(n43334), .I0(n4887), .I1(n4912), .CO(n43335));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_6 (.CI(n43567), 
            .I0(n1430), .I1(GND_net), .CO(n43568));
    SB_LUT4 add_1039_18_lut (.I0(GND_net), .I1(n4888), .I2(n4913), .I3(n43333), 
            .O(n425)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1039_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5582_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_495));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5582_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_967_5_lut (.I0(GND_net), 
            .I1(n1431), .I2(VCC_net), .I3(n43566), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1039_18 (.CI(n43333), .I0(n4888), .I1(n4913), .CO(n43334));
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_967_5 (.CI(n43566), 
            .I0(n1431), .I1(VCC_net), .CO(n43567));
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_23_lut (.I0(GND_net), 
            .I1(n2713), .I2(VCC_net), .I3(n43818), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_227_add_1838_23 (.CI(n43818), 
            .I0(n2713), .I1(VCC_net), .CO(n43819));
    SB_LUT4 add_175_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n43184), .O(n1534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_175_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_add_1838_22_lut (.I0(GND_net), 
            .I1(n2714), .I2(VCC_net), .I3(n43817), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_227_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5586), .I1(duty[9]), .I2(n19_adj_5579), 
            .I3(GND_net), .O(n16_adj_5581));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    \quadrature_decoder(1)_U0  quad_counter0 (.b_prev(b_prev), .n2269(clk16MHz), 
            .GND_net(GND_net), .a_new({a_new[1], Open_0}), .position_31__N_4108(position_31__N_4108), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .n29393(n29393), .n2233(n2233), .encoder0_position({encoder0_position}), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(302[49] 308[6])
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5598));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i39537_3_lut (.I0(n4_adj_5598), .I1(duty[5]), .I2(n11_adj_5584), 
            .I3(GND_net), .O(n55330));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39538_3_lut (.I0(n55330), .I1(duty[6]), .I2(n13_adj_5583), 
            .I3(GND_net), .O(n55331));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38895_4_lut (.I0(n17_adj_5580), .I1(n15_adj_5582), .I2(n13_adj_5583), 
            .I3(n54692), .O(n54688));
    defparam i38895_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39677_4_lut (.I0(n16_adj_5581), .I1(n6_adj_5588), .I2(n19_adj_5579), 
            .I3(n54686), .O(n55470));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39677_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i38991_3_lut (.I0(n55331), .I1(duty[7]), .I2(n15_adj_5582), 
            .I3(GND_net), .O(n54784));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i38991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39761_4_lut (.I0(n54784), .I1(n55470), .I2(n19_adj_5579), 
            .I3(n54688), .O(n55554));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39761_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39762_3_lut (.I0(n55554), .I1(duty[10]), .I2(current[10]), 
            .I3(GND_net), .O(n55555));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39762_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39718_3_lut (.I0(n55555), .I1(duty[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5541));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i39718_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15744_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29820));   // verilog/coms.v(128[12] 303[6])
    defparam i15744_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1876 (.I0(duty[14]), .I1(n24_adj_5541), .I2(duty[12]), 
            .I3(duty[13]), .O(n50454));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1876.LUT_INIT = 16'hfffe;
    SB_LUT4 i15745_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29821));   // verilog/coms.v(128[12] 303[6])
    defparam i15745_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1877 (.I0(duty[14]), .I1(n24_adj_5541), .I2(duty[12]), 
            .I3(duty[13]), .O(n50459));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1877.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1878 (.I0(duty[15]), .I1(current[15]), .I2(n50459), 
            .I3(n50454), .O(n32_adj_5540));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_1878.LUT_INIT = 16'hb3a2;
    SB_LUT4 i15746_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29822));   // verilog/coms.v(128[12] 303[6])
    defparam i15746_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1879 (.I0(duty[18]), .I1(n32_adj_5540), .I2(duty[16]), 
            .I3(duty[17]), .O(n50546));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1879.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1880 (.I0(duty[18]), .I1(n32_adj_5540), .I2(duty[16]), 
            .I3(duty[17]), .O(n50549));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1880.LUT_INIT = 16'h8000;
    SB_LUT4 i40323_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56116));
    defparam i40323_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1881 (.I0(duty[19]), .I1(current[15]), .I2(n50549), 
            .I3(n50546), .O(n40));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_1881.LUT_INIT = 16'hb3a2;
    SB_LUT4 i33743_rep_51_3_lut (.I0(encoder0_position_scaled_23__N_327[30]), 
            .I1(n896), .I2(n861), .I3(GND_net), .O(n52856));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i33743_rep_51_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1882 (.I0(duty[22]), .I1(n40), .I2(duty[20]), 
            .I3(duty[21]), .O(n50599));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1882.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1883 (.I0(duty[22]), .I1(n40), .I2(duty[20]), 
            .I3(duty[21]), .O(n50597));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1883.LUT_INIT = 16'h8000;
    SB_LUT4 i15747_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29823));   // verilog/coms.v(128[12] 303[6])
    defparam i15747_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22640_4_lut (.I0(n535), .I1(n2431), .I2(n2432), .I3(n2433), 
            .O(n36710));
    defparam i22640_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1884 (.I0(n2429), .I1(n2430), .I2(GND_net), .I3(GND_net), 
            .O(n51996));
    defparam i1_2_lut_adj_1884.LUT_INIT = 16'h8888;
    SB_LUT4 i21963_2_lut (.I0(duty[2]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4927));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21963_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i21962_2_lut (.I0(duty[3]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4926));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21962_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i21961_2_lut (.I0(duty[4]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4925));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21961_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i21960_2_lut (.I0(duty[5]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4924));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21960_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i21959_2_lut (.I0(duty[6]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4923));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21959_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i7_3_lut (.I0(encoder0_position_scaled_23__N_327[6]), 
            .I1(n27), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n538));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i635_rep_31_3_lut (.I0(n928), 
            .I1(n995), .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i635_rep_31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21958_2_lut (.I0(duty[7]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4922));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21958_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i8_3_lut (.I0(encoder0_position_scaled_23__N_327[7]), 
            .I1(n26), .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), 
            .O(n537));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1797_3_lut (.I0(n537), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21957_2_lut (.I0(duty[8]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4921));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21957_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i21956_2_lut (.I0(duty[9]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4920));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21956_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i9_3_lut (.I0(encoder0_position_scaled_23__N_327[8]), 
            .I1(n25_adj_5486), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n536));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1729_3_lut (.I0(n536), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1796_3_lut (.I0(n2633), 
            .I1(n2700), .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21955_2_lut (.I0(duty[10]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4919));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21955_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i10_3_lut (.I0(encoder0_position_scaled_23__N_327[9]), 
            .I1(n24_adj_5487), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n535));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15748_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29824));   // verilog/coms.v(128[12] 303[6])
    defparam i15748_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1661_3_lut (.I0(n535), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1728_3_lut (.I0(n2533), 
            .I1(n2600), .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1795_3_lut (.I0(n2632), 
            .I1(n2699), .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1794_3_lut (.I0(n2631), 
            .I1(n2698), .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21954_2_lut (.I0(duty[11]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4918));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21954_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1793_3_lut (.I0(n2630), 
            .I1(n2697), .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40374_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56167));
    defparam i40374_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1885 (.I0(n2414), .I1(n50765), .I2(n2415), .I3(n51806), 
            .O(n51812));
    defparam i1_4_lut_adj_1885.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1792_3_lut (.I0(n2629), 
            .I1(n2696), .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i14_3_lut (.I0(encoder0_position_scaled_23__N_327[13]), 
            .I1(n20_adj_5491), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n531));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1389_3_lut (.I0(n531), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1456_3_lut (.I0(n2133), 
            .I1(n2200), .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1523_3_lut (.I0(n2232), 
            .I1(n2299), .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1590_3_lut (.I0(n2331), 
            .I1(n2398), .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1657_3_lut (.I0(n2430), 
            .I1(n2497), .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1724_3_lut (.I0(n2529), 
            .I1(n2596), .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1791_3_lut (.I0(n2628), 
            .I1(n2695), .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i15_3_lut (.I0(encoder0_position_scaled_23__N_327[14]), 
            .I1(n19_adj_5492), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n530));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1321_3_lut (.I0(n530), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1388_3_lut (.I0(n2033), 
            .I1(n2100), .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1455_3_lut (.I0(n2132), 
            .I1(n2199), .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1522_3_lut (.I0(n2231), 
            .I1(n2298), .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1589_3_lut (.I0(n2330), 
            .I1(n2397), .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1656_rep_40_3_lut (.I0(n2429), 
            .I1(n2496), .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1656_rep_40_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1886 (.I0(n2417), .I1(n51996), .I2(n2421), .I3(n36710), 
            .O(n51794));
    defparam i1_4_lut_adj_1886.LUT_INIT = 16'hfefa;
    SB_LUT4 i15749_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29825));   // verilog/coms.v(128[12] 303[6])
    defparam i15749_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40145_4_lut (.I0(n2412), .I1(n51794), .I2(n51812), .I3(n2413), 
            .O(n2445));
    defparam i40145_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i40416_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56209));
    defparam i40416_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position_scaled_23__N_327[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5618));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1723_3_lut (.I0(n2528), 
            .I1(n2595), .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1790_3_lut (.I0(n2627), 
            .I1(n2694), .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i16_3_lut (.I0(encoder0_position_scaled_23__N_327[15]), 
            .I1(n18_adj_5493), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n529));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1253_rep_20_3_lut (.I0(n529), 
            .I1(n1901), .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1253_rep_20_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1320_3_lut (.I0(n1933), 
            .I1(n2000), .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1387_3_lut (.I0(n2032), 
            .I1(n2099), .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1454_3_lut (.I0(n2131), 
            .I1(n2198), .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1521_3_lut (.I0(n2230), 
            .I1(n2297), .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1588_3_lut (.I0(n2329), 
            .I1(n2396), .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1655_3_lut (.I0(n2428), 
            .I1(n2495), .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39478_3_lut (.I0(n2626), .I1(n2693), .I2(n2643), .I3(GND_net), 
            .O(n2725));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39478_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21953_2_lut (.I0(duty[12]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4917));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21953_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i17_3_lut (.I0(encoder0_position_scaled_23__N_327[16]), 
            .I1(n17_adj_5494), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n528));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1185_3_lut (.I0(n528), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1252_3_lut (.I0(n1833), 
            .I1(n1900), .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1319_3_lut (.I0(n1932), 
            .I1(n1999), .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1386_3_lut (.I0(n2031), 
            .I1(n2098), .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1453_3_lut (.I0(n2130), 
            .I1(n2197), .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21764_1_lut_2_lut (.I0(n24565), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n2573));
    defparam i21764_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1520_3_lut (.I0(n2229), 
            .I1(n2296), .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1587_3_lut (.I0(n2328), 
            .I1(n2395), .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15750_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29826));   // verilog/coms.v(128[12] 303[6])
    defparam i15750_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i572_3_lut_4_lut (.I0(n861), 
            .I1(encoder0_position_scaled_23__N_327[31]), .I2(n52838), .I3(n49477), 
            .O(n932));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i572_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1579_3_lut (.I0(n2320), 
            .I1(n2387), .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i568_3_lut_4_lut (.I0(n861), 
            .I1(encoder0_position_scaled_23__N_327[31]), .I2(n52856), .I3(n49469), 
            .O(n928));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i568_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1654_rep_37_3_lut (.I0(n2427), 
            .I1(n2494), .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1654_rep_37_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22572_3_lut (.I0(n536), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n36642));
    defparam i22572_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1721_3_lut (.I0(n2526), 
            .I1(n2593), .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1788_3_lut (.I0(n2625), 
            .I1(n2692), .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i18_3_lut (.I0(encoder0_position_scaled_23__N_327[17]), 
            .I1(n16_adj_5495), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n527));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1117_3_lut (.I0(n527), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1184_3_lut (.I0(n1733), 
            .I1(n1800), .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1251_3_lut (.I0(n1832), 
            .I1(n1899), .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1318_3_lut (.I0(n1931), 
            .I1(n1998), .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1385_3_lut (.I0(n2030), 
            .I1(n2097), .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1452_rep_48_3_lut (.I0(n2129), 
            .I1(n2196), .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1452_rep_48_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1519_3_lut (.I0(n2228), 
            .I1(n2295), .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1586_3_lut (.I0(n2327), 
            .I1(n2394), .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15751_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29827));   // verilog/coms.v(128[12] 303[6])
    defparam i15751_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1653_rep_43_3_lut (.I0(n2426), 
            .I1(n2493), .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1653_rep_43_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1720_3_lut (.I0(n2525), 
            .I1(n2592), .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1787_3_lut (.I0(n2624), 
            .I1(n2691), .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i19_3_lut (.I0(encoder0_position_scaled_23__N_327[18]), 
            .I1(n15_adj_5496), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n526));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1049_3_lut (.I0(n526), .I1(n1601), 
            .I2(n1554_adj_5610), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1116_3_lut (.I0(n1633), 
            .I1(n1700), .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1183_3_lut (.I0(n1732), 
            .I1(n1799), .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15183_3_lut (.I0(deadband[0]), .I1(\data_in_frame[16] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29259));   // verilog/coms.v(128[12] 303[6])
    defparam i15183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1250_3_lut (.I0(n1831), 
            .I1(n1898), .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1317_3_lut (.I0(n1930), 
            .I1(n1997), .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_1887 (.I0(n2_adj_5509), .I1(n3_adj_5508), 
            .I2(encoder0_position_scaled_23__N_327[31]), .I3(GND_net), .O(n51706));
    defparam i1_2_lut_3_lut_adj_1887.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1384_3_lut (.I0(n2029), 
            .I1(n2096), .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1451_rep_45_3_lut (.I0(n2128), 
            .I1(n2195), .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1451_rep_45_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1518_3_lut (.I0(n2227), 
            .I1(n2294), .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1585_3_lut (.I0(n2326), 
            .I1(n2393), .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1652_rep_38_3_lut (.I0(n2425), 
            .I1(n2492), .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1652_rep_38_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1719_3_lut (.I0(n2524), 
            .I1(n2591), .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1786_3_lut (.I0(n2623), 
            .I1(n2690), .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i981_rep_26_3_lut (.I0(n525), 
            .I1(n1501), .I2(n1455), .I3(GND_net), .O(n1533_adj_5609));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i981_rep_26_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1048_3_lut (.I0(n1533_adj_5609), 
            .I1(n1600), .I2(n1554_adj_5610), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33741_2_lut_3_lut (.I0(n2_adj_5509), .I1(n3_adj_5508), .I2(n5_adj_5482), 
            .I3(GND_net), .O(n49468));
    defparam i33741_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1115_3_lut (.I0(n1632), 
            .I1(n1699), .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1182_3_lut (.I0(n1731), 
            .I1(n1798), .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1249_3_lut (.I0(n1830), 
            .I1(n1897), .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1316_3_lut (.I0(n1929), 
            .I1(n1996), .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5477));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1383_3_lut (.I0(n2028), 
            .I1(n2095), .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1450_rep_46_3_lut (.I0(n2127), 
            .I1(n2194), .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1450_rep_46_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1517_3_lut (.I0(n2226), 
            .I1(n2293), .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1584_3_lut (.I0(n2325), 
            .I1(n2392), .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5476));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1651_rep_39_3_lut (.I0(n2424), 
            .I1(n2491), .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1651_rep_39_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40496_1_lut_4_lut (.I0(current[15]), .I1(duty[23]), .I2(n50597), 
            .I3(n50599), .O(n56288));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i40496_1_lut_4_lut.LUT_INIT = 16'h4c5d;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1718_3_lut (.I0(n2523), 
            .I1(n2590), .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1785_3_lut (.I0(n2622), 
            .I1(n2689), .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532_adj_5608));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1047_3_lut (.I0(n1532_adj_5608), 
            .I1(n1599), .I2(n1554_adj_5610), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1114_3_lut (.I0(n1631), 
            .I1(n1698), .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1181_3_lut (.I0(n1730), 
            .I1(n1797), .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1248_3_lut (.I0(n1829), 
            .I1(n1896), .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21763_2_lut (.I0(n24565), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n35823));
    defparam i21763_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1888 (.I0(n2525), .I1(n2527), .I2(n2524), .I3(n2523), 
            .O(n51530));
    defparam i1_4_lut_adj_1888.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_4_lut (.I0(current[15]), .I1(duty[23]), .I2(n50597), 
            .I3(n50599), .O(n209));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb3a2;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1315_3_lut (.I0(n1928), 
            .I1(n1995), .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1382_3_lut (.I0(n2027), 
            .I1(n2094), .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i769_rep_29_3_lut (.I0(n1126), 
            .I1(n1193), .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i769_rep_29_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1449_rep_50_3_lut (.I0(n2126), 
            .I1(n2193), .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1449_rep_50_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1516_3_lut (.I0(n2225), 
            .I1(n2292), .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1583_3_lut (.I0(n2324), 
            .I1(n2391), .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1650_3_lut (.I0(n2423), 
            .I1(n2490), .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1717_3_lut (.I0(n2522), 
            .I1(n2589), .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1784_3_lut (.I0(n2621), 
            .I1(n2688), .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1889 (.I0(n2526), .I1(n51530), .I2(n2522), .I3(n2528), 
            .O(n51532));
    defparam i1_4_lut_adj_1889.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i836_3_lut.LUT_INIT = 16'hacac;
    motorControl control (.GND_net(GND_net), .\Kp[8] (Kp[8]), .\Ki[1] (Ki[1]), 
            .\PID_CONTROLLER.integral_23__N_3996 ({\PID_CONTROLLER.integral_23__N_3996 }), 
            .\Ki[0] (Ki[0]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[2] (Ki[2]), 
            .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[3] (Ki[3]), .\Kp[9] (Kp[9]), 
            .\Ki[15] (Ki[15]), .\Kp[10] (Kp[10]), .\Ki[4] (Ki[4]), .\Kp[11] (Kp[11]), 
            .\Ki[5] (Ki[5]), .IntegralLimit({IntegralLimit}), .\Ki[6] (Ki[6]), 
            .\Ki[7] (Ki[7]), .\Kp[12] (Kp[12]), .\Kp[3] (Kp[3]), .\Ki[9] (Ki[9]), 
            .PWMLimit({PWMLimit}), .\Kp[4] (Kp[4]), .\Kp[14] (Kp[14]), 
            .\Kp[5] (Kp[5]), .\Kp[1] (Kp[1]), .\Kp[2] (Kp[2]), .\Kp[0] (Kp[0]), 
            .\Kp[13] (Kp[13]), .\Ki[8] (Ki[8]), .\Ki[10] (Ki[10]), .\Kp[15] (Kp[15]), 
            .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .duty({duty}), .clk16MHz(clk16MHz), 
            .control_update(control_update), .deadband({deadband}), .VCC_net(VCC_net), 
            .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), .n29289(n29289), 
            .setpoint({setpoint}), .motor_state({motor_state}), .n29804(n29804), 
            .n29803(n29803), .n29802(n29802), .n29801(n29801), .n29800(n29800), 
            .n29799(n29799), .n29798(n29798), .n29797(n29797), .n29796(n29796), 
            .n29795(n29795), .n29794(n29794), .n29793(n29793), .n29792(n29792), 
            .n29791(n29791), .n29790(n29790), .n29789(n29789), .n29788(n29788), 
            .n29787(n29787), .n29786(n29786), .n29785(n29785), .n29784(n29784), 
            .n29783(n29783), .n29782(n29782)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(288[16] 300[4])
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1046_3_lut (.I0(n1531), 
            .I1(n1598), .I2(n1554_adj_5610), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1113_3_lut (.I0(n1630), 
            .I1(n1697), .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1180_3_lut (.I0(n1729), 
            .I1(n1796), .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1247_3_lut (.I0(n1828), 
            .I1(n1895), .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1314_3_lut (.I0(n1927), 
            .I1(n1994), .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1381_rep_18_3_lut (.I0(n2026), 
            .I1(n2093), .I2(n2049), .I3(GND_net), .O(n52823));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1381_rep_18_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21668_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27117), .I3(n1650), .O(n35728));   // verilog/TinyFPGA_B.v(386[7:11])
    defparam i21668_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfbb;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1448_rep_47_3_lut (.I0(n52823), 
            .I1(n2192), .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1448_rep_47_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1515_3_lut (.I0(n2224), 
            .I1(n2291), .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1582_3_lut (.I0(n2323), 
            .I1(n2390), .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1649_3_lut (.I0(n2422), 
            .I1(n2489), .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1716_3_lut (.I0(n2521), 
            .I1(n2588), .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1783_3_lut (.I0(n2620), 
            .I1(n2687), .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27117), .I3(GND_net), .O(n7593));   // verilog/TinyFPGA_B.v(386[7:11])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5588));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38893_2_lut_4_lut (.I0(current[8]), .I1(duty[8]), .I2(current[4]), 
            .I3(duty[4]), .O(n54686));
    defparam i38893_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27117), .I3(n1650), .O(n7974));   // verilog/TinyFPGA_B.v(386[7:11])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5586));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_1890 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27117), .I3(GND_net), .O(n27118));   // verilog/TinyFPGA_B.v(386[7:11])
    defparam i1_2_lut_3_lut_adj_1890.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_4_lut_adj_1891 (.I0(n2529), .I1(n36642), .I2(n2530), .I3(n2531), 
            .O(n49761));
    defparam i1_4_lut_adj_1891.LUT_INIT = 16'ha080;
    SB_LUT4 unary_minus_19_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5475));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1892 (.I0(n2519), .I1(n2520), .I2(n2521), .I3(n51532), 
            .O(n51538));
    defparam i1_4_lut_adj_1892.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1893 (.I0(n2517), .I1(n2518), .I2(n51538), .I3(n49761), 
            .O(n51544));
    defparam i1_4_lut_adj_1893.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1894 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n51544), 
            .O(n51550));
    defparam i1_4_lut_adj_1894.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_19_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5474));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i40118_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n51550), 
            .O(n2544));
    defparam i40118_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1646_3_lut (.I0(n2419), 
            .I1(n2486), .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1713_3_lut (.I0(n2518), 
            .I1(n2585), .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1727_3_lut (.I0(n2532), 
            .I1(n2599), .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1726_3_lut (.I0(n2531), 
            .I1(n2598), .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n28664), 
            .I3(rx_data_ready), .O(n48270));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i13_3_lut_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3777[2]), .O(n28664));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13_3_lut_4_lut_4_lut.LUT_INIT = 16'h2505;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1895 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3777[2]), .O(n48565));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut_adj_1895.LUT_INIT = 16'h2000;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1725_3_lut (.I0(n2530), 
            .I1(n2597), .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n56302_bdd_4_lut (.I0(n56302), .I1(duty[0]), .I2(n270), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_11[0]));
    defparam n56302_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1037_3_lut (.I0(n1522), 
            .I1(n1589), .I2(n1554_adj_5610), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1896 (.I0(n2628), .I1(n2622), .I2(GND_net), .I3(GND_net), 
            .O(n51864));
    defparam i1_2_lut_adj_1896.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1897 (.I0(n2624), .I1(n2627), .I2(n2623), .I3(n2625), 
            .O(n51872));
    defparam i1_4_lut_adj_1897.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1104_3_lut (.I0(n1621), 
            .I1(n1688), .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1171_3_lut (.I0(n1720), 
            .I1(n1787), .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1238_3_lut (.I0(n1819), 
            .I1(n1886), .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15345_3_lut (.I0(deadband[19]), .I1(\data_in_frame[14] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29421));   // verilog/coms.v(128[12] 303[6])
    defparam i15345_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i23_3_lut (.I0(encoder0_position_scaled_23__N_327[22]), 
            .I1(n11_adj_5500), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n522));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1898 (.I0(n2621), .I1(n51864), .I2(n2620), .I3(n2626), 
            .O(n51874));
    defparam i1_4_lut_adj_1898.LUT_INIT = 16'hfffe;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 i21994_2_lut_2_lut (.I0(n296), .I1(n356), .I2(GND_net), .I3(GND_net), 
            .O(n4883));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i21994_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i777_3_lut (.I0(n522), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22570_3_lut (.I0(n537), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n36640));
    defparam i22570_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1045_3_lut (.I0(n1530), 
            .I1(n1597), .I2(n1554_adj_5610), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33772_4_lut_4_lut_4_lut (.I0(hall1), .I1(commutation_state[2]), 
            .I2(hall2), .I3(hall3), .O(n49501));
    defparam i33772_4_lut_4_lut_4_lut.LUT_INIT = 16'hd504;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1305_3_lut (.I0(n1918), 
            .I1(n1985), .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5473));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5472));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1112_3_lut (.I0(n1629), 
            .I1(n1696), .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5471));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39476_3_lut (.I0(n1827), .I1(n1894), .I2(n1851), .I3(GND_net), 
            .O(n1926));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam i39476_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1313_3_lut (.I0(n1926), 
            .I1(n1993), .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1380_3_lut (.I0(n2025), 
            .I1(n2092), .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1447_rep_49_3_lut (.I0(n2124), 
            .I1(n2191), .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1447_rep_49_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1514_3_lut (.I0(n2223), 
            .I1(n2290), .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1581_3_lut (.I0(n2322), 
            .I1(n2389), .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1648_3_lut (.I0(n2421), 
            .I1(n2488), .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1715_3_lut (.I0(n2520), 
            .I1(n2587), .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1899 (.I0(n2618), .I1(n51874), .I2(n2619), .I3(n51872), 
            .O(n51880));
    defparam i1_4_lut_adj_1899.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1900 (.I0(n2629), .I1(n36640), .I2(n2630), .I3(n2631), 
            .O(n49802));
    defparam i1_4_lut_adj_1900.LUT_INIT = 16'ha080;
    SB_LUT4 unary_minus_19_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5470));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1782_3_lut (.I0(n2619), 
            .I1(n2686), .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1372_3_lut (.I0(n2017), 
            .I1(n2084), .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1901 (.I0(n2616), .I1(n2617), .I2(n49802), .I3(n51880), 
            .O(n51886));
    defparam i1_4_lut_adj_1901.LUT_INIT = 16'hfffe;
    SB_LUT4 i15184_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position_scaled[10]), 
            .I2(n24373), .I3(GND_net), .O(n29260));   // verilog/coms.v(128[12] 303[6])
    defparam i15184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21952_2_lut (.I0(duty[13]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4916));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21952_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1902 (.I0(n2613), .I1(n2614), .I2(n2615), .I3(n51886), 
            .O(n51892));
    defparam i1_4_lut_adj_1902.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1439_3_lut (.I0(n2116), 
            .I1(n2183), .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40089_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n51892), 
            .O(n2643));
    defparam i40089_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_19_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5469));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1506_3_lut (.I0(n2215), 
            .I1(n2282), .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1573_3_lut (.I0(n2314), 
            .I1(n2381), .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15752_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29828));   // verilog/coms.v(128[12] 303[6])
    defparam i15752_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i20_3_lut (.I0(encoder0_position_scaled_23__N_327[19]), 
            .I1(n14_adj_5497), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n525));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15346_3_lut (.I0(deadband[18]), .I1(\data_in_frame[14] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29422));   // verilog/coms.v(128[12] 303[6])
    defparam i15346_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21951_2_lut (.I0(duty[14]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n4915));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i21951_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i24_3_lut (.I0(encoder0_position_scaled_23__N_327[23]), 
            .I1(n10_adj_5501), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n521));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i709_rep_30_3_lut (.I0(n521), 
            .I1(n1101), .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i709_rep_30_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1712_3_lut (.I0(n2517), 
            .I1(n2584), .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_20_i15_2_lut (.I0(duty[7]), .I1(n339), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5551));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i13_2_lut (.I0(duty[6]), .I1(n340), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5552));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1044_3_lut (.I0(n1529), 
            .I1(n1596), .I2(n1554_adj_5610), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_20_i19_2_lut (.I0(duty[9]), .I1(n337), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5543));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1111_rep_25_3_lut (.I0(n1628), 
            .I1(n1695), .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1111_rep_25_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1178_3_lut (.I0(n1727), 
            .I1(n1794), .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1640_rep_36_3_lut (.I0(n2413), 
            .I1(n2480), .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1640_rep_36_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_20_i17_2_lut (.I0(duty[8]), .I1(n338), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5549));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i7_2_lut (.I0(duty[3]), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5556));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1245_3_lut (.I0(n1826), 
            .I1(n1893), .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_20_i9_2_lut (.I0(duty[4]), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5554));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1779_3_lut (.I0(n2616), 
            .I1(n2683), .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_20_i11_2_lut (.I0(duty[5]), .I1(n341), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5553));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5599));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1312_3_lut (.I0(n1925), 
            .I1(n1992), .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1379_3_lut (.I0(n2024), 
            .I1(n2091_adj_5611), .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1446_3_lut (.I0(n2123), 
            .I1(n2190), .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5601));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5578));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1513_3_lut (.I0(n2222), 
            .I1(n2289), .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1580_3_lut (.I0(n2321), 
            .I1(n2388), .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5577));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1647_3_lut (.I0(n2420), 
            .I1(n2487), .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5574));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i5_2_lut (.I0(duty[2]), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5558));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38536_4_lut (.I0(n11_adj_5553), .I1(n9_adj_5554), .I2(n7_adj_5556), 
            .I3(n5_adj_5558), .O(n54328));
    defparam i38536_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_20_i8_3_lut (.I0(n342), .I1(n338), .I2(n17_adj_5549), 
            .I3(GND_net), .O(n8_adj_5555));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1714_3_lut (.I0(n2519), 
            .I1(n2586), .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1781_3_lut (.I0(n2618), 
            .I1(n2685), .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_20_i6_3_lut (.I0(n344), .I1(n343), .I2(n7_adj_5556), 
            .I3(GND_net), .O(n6_adj_5557));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i21_3_lut (.I0(encoder0_position_scaled_23__N_327[20]), 
            .I1(n13_adj_5498), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n524));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i16_3_lut (.I0(n8_adj_5555), .I1(n337), .I2(n19_adj_5543), 
            .I3(GND_net), .O(n16_adj_5550));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36988_3_lut (.I0(duty[17]), .I1(duty[19]), .I2(n330), .I3(GND_net), 
            .O(n52728));
    defparam i36988_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i36992_3_lut (.I0(duty[21]), .I1(duty[15]), .I2(n330), .I3(GND_net), 
            .O(n52732));
    defparam i36992_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i37063_4_lut (.I0(duty[20]), .I1(n52728), .I2(duty[22]), .I3(n330), 
            .O(n52805));
    defparam i37063_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i913_3_lut (.I0(n524), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1641_3_lut (.I0(n2414), 
            .I1(n2481), .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_20_i4_3_lut (.I0(n54237), .I1(n345), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_5559));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39581_3_lut (.I0(n4_adj_5559), .I1(n341), .I2(n11_adj_5553), 
            .I3(GND_net), .O(n55374));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5588_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_514));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5588_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1780_3_lut (.I0(n2617), 
            .I1(n2684), .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15347_3_lut (.I0(deadband[17]), .I1(\data_in_frame[14] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29423));   // verilog/coms.v(128[12] 303[6])
    defparam i15347_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5590_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_523));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5590_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1708_3_lut (.I0(n2513), 
            .I1(n2580), .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39582_3_lut (.I0(n55374), .I1(n340), .I2(n13_adj_5552), .I3(GND_net), 
            .O(n55375));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38928_4_lut (.I0(n17_adj_5549), .I1(n15_adj_5551), .I2(n13_adj_5552), 
            .I3(n54328), .O(n54721));
    defparam i38928_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39681_4_lut (.I0(n16_adj_5550), .I1(n6_adj_5557), .I2(n19_adj_5543), 
            .I3(n54718), .O(n55474));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39681_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39470_3_lut (.I0(n55375), .I1(n339), .I2(n15_adj_5551), .I3(GND_net), 
            .O(n55263));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1707_3_lut (.I0(n2512), 
            .I1(n2579), .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39739_4_lut (.I0(n55263), .I1(n55474), .I2(n19_adj_5543), 
            .I3(n54721), .O(n55532));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39739_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39740_3_lut (.I0(n55532), .I1(n336), .I2(duty[10]), .I3(GND_net), 
            .O(n55533));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39740_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15348_3_lut (.I0(deadband[16]), .I1(\data_in_frame[14] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29424));   // verilog/coms.v(128[12] 303[6])
    defparam i15348_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i39712_3_lut (.I0(n55533), .I1(n335), .I2(duty[11]), .I3(GND_net), 
            .O(n55505));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i39712_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_20_i26_3_lut (.I0(n55505), .I1(n334), .I2(duty[12]), 
            .I3(GND_net), .O(n26_adj_5542));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7_4_lut_adj_1903 (.I0(duty[18]), .I1(n26_adj_5542), .I2(n330), 
            .I3(duty[23]), .O(n20));
    defparam i7_4_lut_adj_1903.LUT_INIT = 16'h2100;
    SB_LUT4 i11_4_lut (.I0(n330), .I1(n52805), .I2(n52732), .I3(duty[13]), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i38590_4_lut (.I0(duty[16]), .I1(n20), .I2(duty[14]), .I3(n330), 
            .O(n54298));
    defparam i38590_4_lut.LUT_INIT = 16'h8004;
    SB_LUT4 mux_15_i1_3_lut (.I0(current[0]), .I1(n2091), .I2(n209), .I3(GND_net), 
            .O(n270));   // verilog/TinyFPGA_B.v(112[16] 114[10])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut_adj_1904 (.I0(n54298), .I1(pwm_setpoint_23__N_263), 
            .I2(n296), .I3(n24), .O(n10832));
    defparam i14_4_lut_adj_1904.LUT_INIT = 16'hcac0;
    SB_LUT4 i15246_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n24373), .I3(GND_net), .O(n29322));   // verilog/coms.v(128[12] 303[6])
    defparam i15246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15247_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n24373), .I3(GND_net), .O(n29323));   // verilog/coms.v(128[12] 303[6])
    defparam i15247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1310_3_lut (.I0(n1923), 
            .I1(n1990), .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15352_3_lut (.I0(deadband[13]), .I1(\data_in_frame[15] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29428));   // verilog/coms.v(128[12] 303[6])
    defparam i15352_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15353_3_lut (.I0(deadband[12]), .I1(\data_in_frame[15] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29429));   // verilog/coms.v(128[12] 303[6])
    defparam i15353_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15354_3_lut (.I0(deadband[11]), .I1(\data_in_frame[15] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29430));   // verilog/coms.v(128[12] 303[6])
    defparam i15354_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15355_3_lut (.I0(deadband[10]), .I1(\data_in_frame[15] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29431));   // verilog/coms.v(128[12] 303[6])
    defparam i15355_3_lut.LUT_INIT = 16'hacac;
    EEPROM eeprom (.clk16MHz(clk16MHz), .\state[3] (state_adj_5747[3]), 
           .n6(n6_adj_5650), .GND_net(GND_net), .read(read), .\state[0] (state_adj_5716[0]), 
           .enable_slow_N_4393(enable_slow_N_4393), .n6271({n6272}), .\state[1] (state_adj_5716[1]), 
           .n48226(n48226), .VCC_net(VCC_net), .n36101(n36101), .n49533(n49533), 
           .n49611(n49611), .n48264(n48264), .n29303(n29303), .rw(rw), 
           .n48368(n48368), .data_ready(data_ready), .n7354(n7354), .\state[2] (state_adj_5747[2]), 
           .\state_7__N_4290[0] (state_7__N_4290[0]), .n4(n4), .n4_adj_19(n4_adj_5459), 
           .n35819(n35819), .scl_enable(scl_enable), .n26(n26_adj_5594), 
           .\state_7__N_4306[3] (state_7__N_4306[3]), .n7936(n7936), .sda_enable(sda_enable), 
           .n29357(n29357), .\saved_addr[0] (saved_addr[0]), .\state[0]_adj_20 (state_adj_5747[0]), 
           .n29269(n29269), .data({data}), .n29268(n29268), .n29267(n29267), 
           .n29266(n29266), .n29265(n29265), .n29264(n29264), .n29263(n29263), 
           .n10(n10_adj_5536), .n10_adj_21(n10_adj_5617), .n8(n8_adj_5657), 
           .n29727(n29727), .n54311(n54311), .n27267(n27267), .n27262(n27262), 
           .scl(scl), .sda_out(sda_out)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(398[10] 409[6])
    SB_LUT4 i15356_3_lut (.I0(deadband[9]), .I1(\data_in_frame[15] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29432));   // verilog/coms.v(128[12] 303[6])
    defparam i15356_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15248_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5734[1]), .I2(n19731), 
            .I3(n4_adj_5479), .O(n29324));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15248_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i15753_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29829));   // verilog/coms.v(128[12] 303[6])
    defparam i15753_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15357_3_lut (.I0(deadband[8]), .I1(\data_in_frame[15] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29433));   // verilog/coms.v(128[12] 303[6])
    defparam i15357_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15249_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n24373), .I3(GND_net), .O(n29325));   // verilog/coms.v(128[12] 303[6])
    defparam i15249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15358_3_lut (.I0(deadband[7]), .I1(\data_in_frame[16] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29434));   // verilog/coms.v(128[12] 303[6])
    defparam i15358_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15250_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n24373), .I3(GND_net), .O(n29326));   // verilog/coms.v(128[12] 303[6])
    defparam i15250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15361_3_lut (.I0(deadband[6]), .I1(\data_in_frame[16] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29437));   // verilog/coms.v(128[12] 303[6])
    defparam i15361_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15362_3_lut (.I0(deadband[5]), .I1(\data_in_frame[16] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29438));   // verilog/coms.v(128[12] 303[6])
    defparam i15362_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15251_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n24373), .I3(GND_net), .O(n29327));   // verilog/coms.v(128[12] 303[6])
    defparam i15251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15252_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n24373), .I3(GND_net), .O(n29328));   // verilog/coms.v(128[12] 303[6])
    defparam i15252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15253_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n24373), .I3(GND_net), .O(n29329));   // verilog/coms.v(128[12] 303[6])
    defparam i15253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15254_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n24373), .I3(GND_net), .O(n29330));   // verilog/coms.v(128[12] 303[6])
    defparam i15254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15255_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n24373), .I3(GND_net), .O(n29331));   // verilog/coms.v(128[12] 303[6])
    defparam i15255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15363_3_lut (.I0(deadband[4]), .I1(\data_in_frame[16] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29439));   // verilog/coms.v(128[12] 303[6])
    defparam i15363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15256_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n24373), .I3(GND_net), .O(n29332));   // verilog/coms.v(128[12] 303[6])
    defparam i15256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15364_3_lut (.I0(deadband[3]), .I1(\data_in_frame[16] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29440));   // verilog/coms.v(128[12] 303[6])
    defparam i15364_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5468));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15257_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n24373), .I3(GND_net), .O(n29333));   // verilog/coms.v(128[12] 303[6])
    defparam i15257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15258_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n24373), 
            .I3(GND_net), .O(n29334));   // verilog/coms.v(128[12] 303[6])
    defparam i15258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15365_3_lut (.I0(deadband[2]), .I1(\data_in_frame[16] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29441));   // verilog/coms.v(128[12] 303[6])
    defparam i15365_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15366_3_lut (.I0(deadband[1]), .I1(\data_in_frame[16] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29442));   // verilog/coms.v(128[12] 303[6])
    defparam i15366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15259_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n24373), 
            .I3(GND_net), .O(n29335));   // verilog/coms.v(128[12] 303[6])
    defparam i15259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15260_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n24373), 
            .I3(GND_net), .O(n29336));   // verilog/coms.v(128[12] 303[6])
    defparam i15260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15261_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n24373), 
            .I3(GND_net), .O(n29337));   // verilog/coms.v(128[12] 303[6])
    defparam i15261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15262_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n24373), 
            .I3(GND_net), .O(n29338));   // verilog/coms.v(128[12] 303[6])
    defparam i15262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5602));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15263_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n24373), 
            .I3(GND_net), .O(n29339));   // verilog/coms.v(128[12] 303[6])
    defparam i15263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15264_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n24373), 
            .I3(GND_net), .O(n29340));   // verilog/coms.v(128[12] 303[6])
    defparam i15264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15369_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n50602), 
            .I3(GND_net), .O(n29445));   // verilog/coms.v(128[12] 303[6])
    defparam i15369_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15370_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29446));   // verilog/coms.v(128[12] 303[6])
    defparam i15370_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5467));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38909_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n54702));
    defparam i38909_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i15371_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29447));   // verilog/coms.v(128[12] 303[6])
    defparam i15371_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15372_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29448));   // verilog/coms.v(128[12] 303[6])
    defparam i15372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15373_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29449));   // verilog/coms.v(128[12] 303[6])
    defparam i15373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5466));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15374_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29450));   // verilog/coms.v(128[12] 303[6])
    defparam i15374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15754_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29830));   // verilog/coms.v(128[12] 303[6])
    defparam i15754_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5600));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15375_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29451));   // verilog/coms.v(128[12] 303[6])
    defparam i15375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15265_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n24373), 
            .I3(GND_net), .O(n29341));   // verilog/coms.v(128[12] 303[6])
    defparam i15265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15267_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29343));   // verilog/coms.v(128[12] 303[6])
    defparam i15267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22670_4_lut (.I0(n520), .I1(n931), .I2(n932), .I3(n933), 
            .O(n36740));
    defparam i22670_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15376_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29452));   // verilog/coms.v(128[12] 303[6])
    defparam i15376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15377_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29453));   // verilog/coms.v(128[12] 303[6])
    defparam i15377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15269_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29345));   // verilog/coms.v(128[12] 303[6])
    defparam i15269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15270_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29346));   // verilog/coms.v(128[12] 303[6])
    defparam i15270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15271_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29347));   // verilog/coms.v(128[12] 303[6])
    defparam i15271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15378_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29454));   // verilog/coms.v(128[12] 303[6])
    defparam i15378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15379_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29455));   // verilog/coms.v(128[12] 303[6])
    defparam i15379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15273_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29349));   // verilog/coms.v(128[12] 303[6])
    defparam i15273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15380_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29456));   // verilog/coms.v(128[12] 303[6])
    defparam i15380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15755_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29831));   // verilog/coms.v(128[12] 303[6])
    defparam i15755_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15275_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29351));   // verilog/coms.v(128[12] 303[6])
    defparam i15275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15381_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29457));   // verilog/coms.v(128[12] 303[6])
    defparam i15381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15276_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29352));   // verilog/coms.v(128[12] 303[6])
    defparam i15276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15277_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29353));   // verilog/coms.v(128[12] 303[6])
    defparam i15277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15382_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29458));   // verilog/coms.v(128[12] 303[6])
    defparam i15382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15349_3_lut (.I0(deadband[15]), .I1(\data_in_frame[15] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29425));   // verilog/coms.v(128[12] 303[6])
    defparam i15349_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_adj_1905 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5661));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut_adj_1905.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1906 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5660));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut_adj_1906.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1907 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n51630));
    defparam i1_2_lut_adj_1907.LUT_INIT = 16'h8888;
    SB_LUT4 i14_3_lut (.I0(hall2), .I1(hall3), .I2(hall1), .I3(GND_net), 
            .O(n6_adj_5668));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1908 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_264[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_1908.LUT_INIT = 16'h1414;
    SB_LUT4 i15383_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29459));   // verilog/coms.v(128[12] 303[6])
    defparam i15383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut_adj_1909 (.I0(dti_counter[0]), .I1(n14_adj_5660), .I2(n10_adj_5661), 
            .I3(dti_counter[3]), .O(n24565));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut_adj_1909.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1910 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5605));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_1910.LUT_INIT = 16'h7bde;
    SB_LUT4 i15384_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29460));   // verilog/coms.v(128[12] 303[6])
    defparam i15384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i40439_2_lut (.I0(n24565), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_527));
    defparam i40439_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i15385_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n50602), .I3(GND_net), .O(n29461));   // verilog/coms.v(128[12] 303[6])
    defparam i15385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15386_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n50602), .I3(GND_net), .O(n29462));   // verilog/coms.v(128[12] 303[6])
    defparam i15386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1911 (.I0(n927), .I1(n51630), .I2(n928), .I3(n36740), 
            .O(n960));
    defparam i1_4_lut_adj_1911.LUT_INIT = 16'hfefa;
    SB_LUT4 i15387_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n50602), .I3(GND_net), .O(n29463));   // verilog/coms.v(128[12] 303[6])
    defparam i15387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_1_lut_adj_1912 (.I0(current[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut_adj_1912.LUT_INIT = 16'h5555;
    SB_LUT4 i15278_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29354));   // verilog/coms.v(128[12] 303[6])
    defparam i15278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15388_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29464));   // verilog/coms.v(128[12] 303[6])
    defparam i15388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15389_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29465));   // verilog/coms.v(128[12] 303[6])
    defparam i15389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15279_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29355));   // verilog/coms.v(128[12] 303[6])
    defparam i15279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15281_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_4290[0]), 
            .I3(enable_slow_N_4393), .O(n29357));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15281_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_mux_3_i25_3_lut (.I0(encoder0_position_scaled_23__N_327[24]), 
            .I1(n9_adj_5502), .I2(encoder0_position_scaled_23__N_327[31]), 
            .I3(GND_net), .O(n520));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15282_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29358));   // verilog/coms.v(128[12] 303[6])
    defparam i15282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15390_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n50602), .I3(GND_net), .O(n29466));   // verilog/coms.v(128[12] 303[6])
    defparam i15390_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15391_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n50602), .I3(GND_net), .O(n29467));   // verilog/coms.v(128[12] 303[6])
    defparam i15391_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15284_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29360));   // verilog/coms.v(128[12] 303[6])
    defparam i15284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15285_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29361));   // verilog/coms.v(128[12] 303[6])
    defparam i15285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15286_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29362));   // verilog/coms.v(128[12] 303[6])
    defparam i15286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15392_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n50602), .I3(GND_net), .O(n29468));   // verilog/coms.v(128[12] 303[6])
    defparam i15392_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15287_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29363));   // verilog/coms.v(128[12] 303[6])
    defparam i15287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15288_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29364));   // verilog/coms.v(128[12] 303[6])
    defparam i15288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15289_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29365));   // verilog/coms.v(128[12] 303[6])
    defparam i15289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15290_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29366));   // verilog/coms.v(128[12] 303[6])
    defparam i15290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15292_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29368));   // verilog/coms.v(128[12] 303[6])
    defparam i15292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15293_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29369));   // verilog/coms.v(128[12] 303[6])
    defparam i15293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15756_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n50602), .I3(GND_net), .O(n29832));   // verilog/coms.v(128[12] 303[6])
    defparam i15756_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15294_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29370));   // verilog/coms.v(128[12] 303[6])
    defparam i15294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15295_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29371));   // verilog/coms.v(128[12] 303[6])
    defparam i15295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15400_3_lut (.I0(\data_in_frame[20] [7]), .I1(rx_data[7]), 
            .I2(n48646), .I3(GND_net), .O(n29476));   // verilog/coms.v(128[12] 303[6])
    defparam i15400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15401_3_lut (.I0(\data_in_frame[20] [6]), .I1(rx_data[6]), 
            .I2(n48646), .I3(GND_net), .O(n29477));   // verilog/coms.v(128[12] 303[6])
    defparam i15401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15402_3_lut (.I0(\data_in_frame[20] [5]), .I1(rx_data[5]), 
            .I2(n48646), .I3(GND_net), .O(n29478));   // verilog/coms.v(128[12] 303[6])
    defparam i15402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15403_3_lut (.I0(\data_in_frame[20] [4]), .I1(rx_data[4]), 
            .I2(n48646), .I3(GND_net), .O(n29479));   // verilog/coms.v(128[12] 303[6])
    defparam i15403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15404_3_lut (.I0(\data_in_frame[20] [3]), .I1(rx_data[3]), 
            .I2(n48646), .I3(GND_net), .O(n29480));   // verilog/coms.v(128[12] 303[6])
    defparam i15404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15405_3_lut (.I0(\data_in_frame[20] [2]), .I1(rx_data[2]), 
            .I2(n48646), .I3(GND_net), .O(n29481));   // verilog/coms.v(128[12] 303[6])
    defparam i15405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15406_3_lut (.I0(\data_in_frame[20] [1]), .I1(rx_data[1]), 
            .I2(n48646), .I3(GND_net), .O(n29482));   // verilog/coms.v(128[12] 303[6])
    defparam i15406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15296_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29372));   // verilog/coms.v(128[12] 303[6])
    defparam i15296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15407_3_lut (.I0(\data_in_frame[20] [0]), .I1(rx_data[0]), 
            .I2(n48646), .I3(GND_net), .O(n29483));   // verilog/coms.v(128[12] 303[6])
    defparam i15407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15757_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n50602), .I3(GND_net), .O(n29833));   // verilog/coms.v(128[12] 303[6])
    defparam i15757_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15297_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29373));   // verilog/coms.v(128[12] 303[6])
    defparam i15297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15298_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n50602), 
            .I3(GND_net), .O(n29374));   // verilog/coms.v(128[12] 303[6])
    defparam i15298_3_lut.LUT_INIT = 16'hacac;
    coms neopxl_color_23__I_0 (.n29426(n29426), .deadband({deadband}), .clk16MHz(clk16MHz), 
         .n29425(n29425), .n29424(n29424), .n29423(n29423), .n29422(n29422), 
         .GND_net(GND_net), .\data_in_frame[16] ({\data_in_frame[16] }), 
         .rx_data({rx_data}), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n29421(n29421), .\data_in_frame[14] ({\data_in_frame[14] }), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[15] ({\data_in_frame[15] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .n4452(n4452), .\FRAME_MATCHER.i_31__N_2845 (\FRAME_MATCHER.i_31__N_2845 ), 
         .n22902(n22902), .\data_in_frame[3] ({\data_in_frame[3] }), .n29419(n29419), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .\data_in_frame[21] ({\data_in_frame[21] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[22] ({\data_out_frame[22] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[21] ({\data_out_frame[21] }), .n29418(n29418), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .n29417(n29417), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in[1] ({Open_1, Open_2, \data_in[1] [5:4], Open_3, Open_4, 
         Open_5, \data_in[1] [0]}), .\data_in[2] ({Open_6, Open_7, Open_8, 
         \data_in[2] [4], Open_9, \data_in[2] [2], Open_10, Open_11}), 
         .\data_in[3] ({Open_12, Open_13, Open_14, \data_in[3] [4], 
         Open_15, \data_in[3] [2], Open_16, \data_in[3] [0]}), .\data_in[0] ({Open_17, 
         \data_in[0] [6:0]}), .\data_in[1][1] (\data_in[1] [1]), .\data_in[2][5] (\data_in[2] [5]), 
         .\data_in[1][6] (\data_in[1] [6]), .\data_in[1][3] (\data_in[1] [3]), 
         .\data_in[2][0] (\data_in[2] [0]), .\data_in[1][2] (\data_in[1] [2]), 
         .\data_in[2][6] (\data_in[2] [6]), .\data_in[2][3] (\data_in[2] [3]), 
         .\data_in[3][3] (\data_in[3] [3]), .\data_in[3][5] (\data_in[3] [5]), 
         .\data_in[3][6] (\data_in[3] [6]), .\data_in[2][1] (\data_in[2] [1]), 
         .rx_data_ready(rx_data_ready), .n63(n63_adj_5615), .n3303(n3303), 
         .n4599(n4599), .n48672(n48672), .n4(n4_adj_5606), .n48616(n48616), 
         .\data_in_frame[8] ({\data_in_frame[8] }), .n29416(n29416), .n29415(n29415), 
         .\Kp[2] (Kp[2]), .setpoint({setpoint}), .ID({ID}), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .n29411(n29411), .\Kp[3] (Kp[3]), .tx_active(tx_active), .\data_in_frame[20] ({\data_in_frame[20] }), 
         .n29410(n29410), .\Kp[4] (Kp[4]), .\data_in_frame[23] ({\data_in_frame[23] }), 
         .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), .n29409(n29409), 
         .\Kp[5] (Kp[5]), .n29408(n29408), .\Kp[6] (Kp[6]), .n29407(n29407), 
         .\Kp[7] (Kp[7]), .n29406(n29406), .\Kp[8] (Kp[8]), .n29405(n29405), 
         .\Kp[9] (Kp[9]), .n29404(n29404), .\Kp[10] (Kp[10]), .n29403(n29403), 
         .\Kp[11] (Kp[11]), .n29402(n29402), .\Kp[12] (Kp[12]), .n29401(n29401), 
         .\Kp[13] (Kp[13]), .n29400(n29400), .\Kp[14] (Kp[14]), .n29396(n29396), 
         .\Kp[15] (Kp[15]), .n29395(n29395), .\Ki[1] (Ki[1]), .n29394(n29394), 
         .\Ki[2] (Ki[2]), .n29391(n29391), .\Ki[3] (Ki[3]), .n29390(n29390), 
         .\Ki[4] (Ki[4]), .n29389(n29389), .\Ki[5] (Ki[5]), .n29388(n29388), 
         .\Ki[6] (Ki[6]), .n29387(n29387), .\Ki[7] (Ki[7]), .n29386(n29386), 
         .\Ki[8] (Ki[8]), .n29385(n29385), .\Ki[9] (Ki[9]), .n29384(n29384), 
         .\Ki[10] (Ki[10]), .n29378(n29378), .\Ki[11] (Ki[11]), .n29377(n29377), 
         .\Ki[12] (Ki[12]), .n29376(n29376), .\Ki[13] (Ki[13]), .n29375(n29375), 
         .\Ki[14] (Ki[14]), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .n29374(n29374), 
         .\Ki[15] (Ki[15]), .n29373(n29373), .n29372(n29372), .n29371(n29371), 
         .n29370(n29370), .n29369(n29369), .n29368(n29368), .n29366(n29366), 
         .n29365(n29365), .n29364(n29364), .n29363(n29363), .n29362(n29362), 
         .n29361(n29361), .n29360(n29360), .n29358(n29358), .n29355(n29355), 
         .n29354(n29354), .n29353(n29353), .n29352(n29352), .n29351(n29351), 
         .n29349(n29349), .n29347(n29347), .n29346(n29346), .n29345(n29345), 
         .n29343(n29343), .n29341(n29341), .n29340(n29340), .n29339(n29339), 
         .n29338(n29338), .n29337(n29337), .n29336(n29336), .n29335(n29335), 
         .n29334(n29334), .n29333(n29333), .n29332(n29332), .n29331(n29331), 
         .n29330(n29330), .n29329(n29329), .n29328(n29328), .n29327(n29327), 
         .n29326(n29326), .n29325(n29325), .n29323(n29323), .n29322(n29322), 
         .n50602(n50602), .n122(n122), .\FRAME_MATCHER.i_31__N_2843 (\FRAME_MATCHER.i_31__N_2843 ), 
         .n5(n5_adj_5616), .n57092(n57092), .n29321(n29321), .n29957(n29957), 
         .n29956(n29956), .n29955(n29955), .n29954(n29954), .n29953(n29953), 
         .n29952(n29952), .n29951(n29951), .n29950(n29950), .n29949(n29949), 
         .n29948(n29948), .n29947(n29947), .n29946(n29946), .n29945(n29945), 
         .n29944(n29944), .n29943(n29943), .n29942(n29942), .n29941(n29941), 
         .n29940(n29940), .n29939(n29939), .n29938(n29938), .n29937(n29937), 
         .n29936(n29936), .n29935(n29935), .n29934(n29934), .n29933(n29933), 
         .n29932(n29932), .n29931(n29931), .n29930(n29930), .n29929(n29929), 
         .n29928(n29928), .n29927(n29927), .n29926(n29926), .n29925(n29925), 
         .n29924(n29924), .n29923(n29923), .n29922(n29922), .n29921(n29921), 
         .n29920(n29920), .n29919(n29919), .n29918(n29918), .n29917(n29917), 
         .n29916(n29916), .n29915(n29915), .n29914(n29914), .n29913(n29913), 
         .n29912(n29912), .n29911(n29911), .n29910(n29910), .n29909(n29909), 
         .n29908(n29908), .n29907(n29907), .n29906(n29906), .n29905(n29905), 
         .n29904(n29904), .n29903(n29903), .n29902(n29902), .n29901(n29901), 
         .n29900(n29900), .n29899(n29899), .n29898(n29898), .n29897(n29897), 
         .n29896(n29896), .n29895(n29895), .n29894(n29894), .n29893(n29893), 
         .n29892(n29892), .n29891(n29891), .n29890(n29890), .n29889(n29889), 
         .n29888(n29888), .n29887(n29887), .n29886(n29886), .n29885(n29885), 
         .n29884(n29884), .n29883(n29883), .n29882(n29882), .DE_c(DE_c), 
         .LED_c(LED_c), .n29319(n29319), .n29318(n29318), .n29316(n29316), 
         .n29315(n29315), .n29314(n29314), .n29313(n29313), .n29312(n29312), 
         .n29311(n29311), .n29310(n29310), .n29307(n29307), .n29306(n29306), 
         .n29305(n29305), .n29304(n29304), .n29300(n29300), .n29299(n29299), 
         .n29298(n29298), .n29297(n29297), .n29296(n29296), .n29881(n29881), 
         .n29880(n29880), .n29879(n29879), .n29878(n29878), .n29877(n29877), 
         .n29876(n29876), .n29875(n29875), .n29874(n29874), .n29873(n29873), 
         .n29872(n29872), .n29871(n29871), .n29870(n29870), .n29869(n29869), 
         .n29868(n29868), .n29867(n29867), .n29859(n29859), .n29858(n29858), 
         .n29857(n29857), .n29856(n29856), .n29855(n29855), .n29854(n29854), 
         .n29853(n29853), .n29852(n29852), .n29851(n29851), .control_mode({control_mode}), 
         .n29295(n29295), .n29850(n29850), .n29849(n29849), .n29848(n29848), 
         .n29847(n29847), .n29846(n29846), .n29845(n29845), .n29294(n29294), 
         .n29844(n29844), .current_limit({current_limit}), .n29293(n29293), 
         .n29843(n29843), .n29842(n29842), .n29841(n29841), .n29840(n29840), 
         .n29292(n29292), .n29291(n29291), .n29290(n29290), .n29288(n29288), 
         .n29287(n29287), .n29286(n29286), .n48016(n48016), .n29284(n29284), 
         .PWMLimit({PWMLimit}), .n29283(n29283), .n29282(n29282), .n29280(n29280), 
         .neopxl_color({neopxl_color}), .n29279(n29279), .n29278(n29278), 
         .\Ki[0] (Ki[0]), .n29277(n29277), .\Kp[0] (Kp[0]), .n29276(n29276), 
         .IntegralLimit({IntegralLimit}), .n29275(n29275), .n29274(n29274), 
         .n29273(n29273), .n29839(n29839), .n29838(n29838), .n29837(n29837), 
         .n29836(n29836), .n29835(n29835), .n29834(n29834), .n63_adj_6(n63), 
         .n29833(n29833), .n29832(n29832), .n9(n9_adj_5607), .n29831(n29831), 
         .n29830(n29830), .n29829(n29829), .n29828(n29828), .n29260(n29260), 
         .n29259(n29259), .n29827(n29827), .n29826(n29826), .n29825(n29825), 
         .n29824(n29824), .n29823(n29823), .n29822(n29822), .n29821(n29821), 
         .n29820(n29820), .n29256(n29256), .n29819(n29819), .n29818(n29818), 
         .n29817(n29817), .n29816(n29816), .n29815(n29815), .n29814(n29814), 
         .n29813(n29813), .n29812(n29812), .n29811(n29811), .n29810(n29810), 
         .n29809(n29809), .n29808(n29808), .n29807(n29807), .n56702(n56702), 
         .n29762(n29762), .n29761(n29761), .n29760(n29760), .n29759(n29759), 
         .n29758(n29758), .n29757(n29757), .n29756(n29756), .n29755(n29755), 
         .n29754(n29754), .n29753(n29753), .n29752(n29752), .n29751(n29751), 
         .n29726(n29726), .n29725(n29725), .n29724(n29724), .n29723(n29723), 
         .n29722(n29722), .n29721(n29721), .n29720(n29720), .n29719(n29719), 
         .n29718(n29718), .n29717(n29717), .n29716(n29716), .n29707(n29707), 
         .n29706(n29706), .n29705(n29705), .n29704(n29704), .n29703(n29703), 
         .n29702(n29702), .n29701(n29701), .n29687(n29687), .n29686(n29686), 
         .n29685(n29685), .n29666(n29666), .n29665(n29665), .n29664(n29664), 
         .n29663(n29663), .n29662(n29662), .n29661(n29661), .n29660(n29660), 
         .n29659(n29659), .n29658(n29658), .n29657(n29657), .n29656(n29656), 
         .n29655(n29655), .n29654(n29654), .n29653(n29653), .n29652(n29652), 
         .n29651(n29651), .n29650(n29650), .n29649(n29649), .n29648(n29648), 
         .n29646(n29646), .n29645(n29645), .n29644(n29644), .n29643(n29643), 
         .n29483(n29483), .n29482(n29482), .n29481(n29481), .n29480(n29480), 
         .n29479(n29479), .n29478(n29478), .n29477(n29477), .n29476(n29476), 
         .n29468(n29468), .n29467(n29467), .n29466(n29466), .n29465(n29465), 
         .n29464(n29464), .n29463(n29463), .n29462(n29462), .n29461(n29461), 
         .n29460(n29460), .n29459(n29459), .n29458(n29458), .n29457(n29457), 
         .n29456(n29456), .n29455(n29455), .n29454(n29454), .n29453(n29453), 
         .n29452(n29452), .n29451(n29451), .n29450(n29450), .n29449(n29449), 
         .n29448(n29448), .n29447(n29447), .n29446(n29446), .n29445(n29445), 
         .\Kp[1] (Kp[1]), .n29442(n29442), .n29441(n29441), .n29440(n29440), 
         .n29439(n29439), .n29438(n29438), .n29437(n29437), .n29434(n29434), 
         .n29433(n29433), .n29432(n29432), .n29431(n29431), .n29430(n29430), 
         .n29429(n29429), .n29428(n29428), .n5_adj_7(n5_adj_5458), .n50620(n50620), 
         .n24373(n24373), .n48646(n48646), .n48638(n48638), .\state[0] (state_adj_5747[0]), 
         .\state[2] (state_adj_5747[2]), .\state[3] (state_adj_5747[3]), 
         .n7936(n7936), .n28758(n28758), .n29184(n29184), .\r_Bit_Index[0] (r_Bit_Index_adj_5736[0]), 
         .r_SM_Main({r_SM_Main_adj_5734}), .\r_SM_Main_2__N_3848[1] (r_SM_Main_2__N_3848[1]), 
         .VCC_net(VCC_net), .tx_o(tx_o), .n29324(n29324), .n29732(n29732), 
         .n56700(n56700), .n4_adj_8(n4_adj_5479), .tx_enable(tx_enable), 
         .n19731(n19731), .n28762(n28762), .n29186(n29186), .n29420(n29420), 
         .r_SM_Main_adj_16({r_SM_Main}), .r_Rx_Data(r_Rx_Data), .\r_SM_Main_2__N_3777[2] (r_SM_Main_2__N_3777[2]), 
         .n35837(n35837), .RX_N_10(RX_N_10), .n4_adj_12(n4_adj_5595), 
         .n4_adj_13(n4_adj_5539), .n29735(n29735), .\r_Bit_Index[0]_adj_14 (r_Bit_Index[0]), 
         .n48270(n48270), .n29261(n29261), .n4_adj_15(n4_adj_5478), .n29769(n29769), 
         .n29767(n29767), .n29766(n29766), .n48565(n48565), .n29749(n29749), 
         .n29748(n29748), .n29740(n29740), .n27227(n27227), .n27232(n27232)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(254[8] 278[4])
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_5747[0]), .I1(n54311), .I2(n7354), 
            .I3(n10_adj_5536), .O(n8_adj_5657));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_LUT4 i5584_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_500));
    defparam i5584_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i5586_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_509));
    defparam i5586_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i22602_3_lut (.I0(n521), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n36672));
    defparam i22602_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5734[2]), .I1(r_SM_Main_adj_5734[0]), 
            .I2(r_SM_Main_adj_5734[1]), .I3(r_SM_Main_2__N_3848[1]), .O(n56700));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i15317_3_lut_4_lut (.I0(n2233), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_4108), .O(n29393));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15317_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i15316_3_lut_4_lut (.I0(n2274), .I1(b_prev_adj_5545), .I2(a_new_adj_5703[1]), 
            .I3(position_31__N_4108_adj_5546), .O(n29392));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15316_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_4_lut_adj_1913 (.I0(n1029), .I1(n36672), .I2(n1030), .I3(n1031), 
            .O(n49689));
    defparam i1_4_lut_adj_1913.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_227_i1778_3_lut (.I0(n2615), 
            .I1(n2682), .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(322[33:71])
    defparam encoder0_position_scaled_23__I_0_227_i1778_3_lut.LUT_INIT = 16'hacac;
    TLI4970 tli (.\state[0] (state_adj_5724[0]), .\state[1] (state_adj_5724[1]), 
            .state_7__N_4499(state_7__N_4499), .GND_net(GND_net), .\data[12] (data_adj_5722[12]), 
            .clk16MHz(clk16MHz), .VCC_net(VCC_net), .\data[15] (data_adj_5722[15]), 
            .n28640(n28640), .n35803(n35803), .n15(n15_adj_5481), .n35841(n35841), 
            .n6(n6_adj_5537), .n5(n5_adj_5570), .n29966(n29966), .\data[10] (data_adj_5722[10]), 
            .n5_adj_1(n5), .n29965(n29965), .\data[9] (data_adj_5722[9]), 
            .n29959(n29959), .\data[8] (data_adj_5722[8]), .n29958(n29958), 
            .\data[7] (data_adj_5722[7]), .n29320(n29320), .n29317(n29317), 
            .\data[11] (data_adj_5722[11]), .n9(n9_adj_5511), .clk_out(clk_out), 
            .n29308(n29308), .CS_c(CS_c), .n29301(n29301), .\current[0] (current[0]), 
            .n6_adj_2(n6_adj_5571), .n5_adj_3(n5_adj_5538), .n7(n7_adj_5597), 
            .\current[15] (current[15]), .CS_CLK_c(CS_CLK_c), .n29805(n29805), 
            .\data[6] (data_adj_5722[6]), .n29781(n29781), .\data[5] (data_adj_5722[5]), 
            .n29780(n29780), .\current[1] (current[1]), .n29779(n29779), 
            .\current[2] (current[2]), .n29778(n29778), .\current[3] (current[3]), 
            .n29777(n29777), .\current[4] (current[4]), .n29776(n29776), 
            .\current[5] (current[5]), .n29775(n29775), .\current[6] (current[6]), 
            .n29774(n29774), .\current[7] (current[7]), .n29773(n29773), 
            .\current[8] (current[8]), .n29772(n29772), .\current[9] (current[9]), 
            .n29771(n29771), .\current[10] (current[10]), .n29770(n29770), 
            .\current[11] (current[11]), .n29768(n29768), .\data[4] (data_adj_5722[4]), 
            .n29763(n29763), .\data[3] (data_adj_5722[3]), .n29750(n29750), 
            .\data[2] (data_adj_5722[2]), .n29741(n29741), .\data[0] (data_adj_5722[0]), 
            .n29736(n29736), .\data[1] (data_adj_5722[1]), .n29647(n29647), 
            .n27222(n27222), .n27287(n27287), .n27281(n27281), .n27294(n27294), 
            .n27256(n27256)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(411[11] 417[4])
    \quadrature_decoder(1)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .VCC_net(VCC_net), .b_prev(b_prev_adj_5545), 
            .a_new({a_new_adj_5703[1], Open_18}), .position_31__N_4108(position_31__N_4108_adj_5546), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .n2269(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .n29392(n29392), .n2274(n2274)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(310[49] 316[6])
    pwm PWM (.pwm_out(pwm_out), .clk32MHz(clk32MHz), .GND_net(GND_net), 
        .VCC_net(VCC_net), .pwm_setpoint({pwm_setpoint})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(96[6] 101[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, \neo_pixel_transmitter.t0 , 
            GND_net, neopxl_color, \state[1] , \state[0] , n28689, 
            \state_3__N_639[1] , timer, n49594, VCC_net, LED_c, n29258, 
            n29700, n29699, n29698, n29697, n29696, n29695, n29694, 
            n29693, n29692, n29691, n29690, n29689, n29688, n29684, 
            n29683, n29682, n29681, n29680, n29679, n29678, n29677, 
            n29676, n29675, n29674, n29673, n29672, n29671, n29670, 
            n29669, n29668, n29667, NEOPXL_c, n29436) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input GND_net;
    input [23:0]neopxl_color;
    output \state[1] ;
    output \state[0] ;
    output n28689;
    output \state_3__N_639[1] ;
    output [31:0]timer;
    output n49594;
    input VCC_net;
    input LED_c;
    input n29258;
    input n29700;
    input n29699;
    input n29698;
    input n29697;
    input n29696;
    input n29695;
    input n29694;
    input n29693;
    input n29692;
    input n29691;
    input n29690;
    input n29689;
    input n29688;
    input n29684;
    input n29683;
    input n29682;
    input n29681;
    input n29680;
    input n29679;
    input n29678;
    input n29677;
    input n29676;
    input n29675;
    input n29674;
    input n29673;
    input n29672;
    input n29671;
    input n29670;
    input n29669;
    input n29668;
    input n29667;
    output NEOPXL_c;
    input n29436;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire \neo_pixel_transmitter.done_N_847 , n56661, \neo_pixel_transmitter.done , 
        start_N_838, n7, start;
    wire [31:0]n1;
    wire [31:0]n133;
    
    wire n7792;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n29101, n53036, n53037, n53028, n53027, n36592, n51143, 
        n23_adj_5419, n27272, n56371, n56635;
    wire [31:0]color_bit_N_833;
    
    wire n55197, n36459, n45504, n56515, n55259, n56467, n54304;
    wire [3:0]state_3__N_639;
    
    wire n56368;
    wire [31:0]n133_adj_5456;
    
    wire n52931, n52932, n56512, n52926, n52925, n44055, n44054, 
        n44053, n44052, n44051, n27276, n43155, n52408, n44050, 
        n44049, n43154, n52406, n44048, n44047, n43153, n52404, 
        n44046, n44045, n44044, n43152, n52402, n44043, n44042, 
        n44041, n43151, n52400, n43150, n52398, n44040, n29076, 
        n56464, n44039, n44038, n44037, n49519, n44914, n49641, 
        n27135, n43149, n52396, n44036, n44035, n44034, n44033, 
        n44032, n44031, n44030, n44029, n44028, n44027, n44026, 
        n43148, n52394, n43147, n52392, n44025, n44024, n44023, 
        n44022, n43146, n52390, n44021, n44020, n43145, n52388, 
        n44019, n44018, n44017, n43144, n52386, n44016, n44015, 
        n44014, n44013, n43143, n52384, n44012, n44011, n29033, 
        n44010, n43142, n52382, n44009, n44008, n44007, n44006, 
        n46, n44005, n44004, n44003, n44002, n44, n44001, n45, 
        n44000, n43999, n43, n43998, n43997, n43996, n42, n43995, 
        n43994, n40, n43141, n52380, n48, n52, n51, n2586, n10_adj_5453, 
        n7747, n54239, n43140, n52378, n43139, n52376, n43138, 
        n52374, n43137, n52372, n43136;
    wire [31:0]one_wire_N_790;
    
    wire n43135, n43134, n43133, n43132, n43131, n43130, n43129, 
        n43128, n43127, n43126, n43125, n54378, n54379, n54236, 
        n51217, n56632, \neo_pixel_transmitter.done_N_853 , n49637, 
        n52410, n52416, n54242, n49458, n49515, n48656, n103, 
        n16_adj_5454, n6_adj_5455, n49617;
    
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n56661), .D(\neo_pixel_transmitter.done_N_847 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE start_103 (.Q(start), .C(clk16MHz), .E(n7), .D(start_N_838));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_2281__i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n7792), 
            .D(n133[0]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i1 (.Q(bit_ctr[1]), .C(clk16MHz), .E(n7792), 
            .D(n133[1]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i2 (.Q(bit_ctr[2]), .C(clk16MHz), .E(n7792), 
            .D(n133[2]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i3 (.Q(bit_ctr[3]), .C(clk16MHz), .E(n7792), 
            .D(n133[3]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i4 (.Q(bit_ctr[4]), .C(clk16MHz), .E(n7792), 
            .D(n133[4]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i5 (.Q(bit_ctr[5]), .C(clk16MHz), .E(n7792), 
            .D(n133[5]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i6 (.Q(bit_ctr[6]), .C(clk16MHz), .E(n7792), 
            .D(n133[6]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i7 (.Q(bit_ctr[7]), .C(clk16MHz), .E(n7792), 
            .D(n133[7]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i8 (.Q(bit_ctr[8]), .C(clk16MHz), .E(n7792), 
            .D(n133[8]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i9 (.Q(bit_ctr[9]), .C(clk16MHz), .E(n7792), 
            .D(n133[9]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i10 (.Q(bit_ctr[10]), .C(clk16MHz), .E(n7792), 
            .D(n133[10]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i11 (.Q(bit_ctr[11]), .C(clk16MHz), .E(n7792), 
            .D(n133[11]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i12 (.Q(bit_ctr[12]), .C(clk16MHz), .E(n7792), 
            .D(n133[12]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i13 (.Q(bit_ctr[13]), .C(clk16MHz), .E(n7792), 
            .D(n133[13]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i14 (.Q(bit_ctr[14]), .C(clk16MHz), .E(n7792), 
            .D(n133[14]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i15 (.Q(bit_ctr[15]), .C(clk16MHz), .E(n7792), 
            .D(n133[15]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i16 (.Q(bit_ctr[16]), .C(clk16MHz), .E(n7792), 
            .D(n133[16]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i17 (.Q(bit_ctr[17]), .C(clk16MHz), .E(n7792), 
            .D(n133[17]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i18 (.Q(bit_ctr[18]), .C(clk16MHz), .E(n7792), 
            .D(n133[18]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i19 (.Q(bit_ctr[19]), .C(clk16MHz), .E(n7792), 
            .D(n133[19]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i20 (.Q(bit_ctr[20]), .C(clk16MHz), .E(n7792), 
            .D(n133[20]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i21 (.Q(bit_ctr[21]), .C(clk16MHz), .E(n7792), 
            .D(n133[21]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i22 (.Q(bit_ctr[22]), .C(clk16MHz), .E(n7792), 
            .D(n133[22]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i23 (.Q(bit_ctr[23]), .C(clk16MHz), .E(n7792), 
            .D(n133[23]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i24 (.Q(bit_ctr[24]), .C(clk16MHz), .E(n7792), 
            .D(n133[24]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i25 (.Q(bit_ctr[25]), .C(clk16MHz), .E(n7792), 
            .D(n133[25]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i26 (.Q(bit_ctr[26]), .C(clk16MHz), .E(n7792), 
            .D(n133[26]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i27 (.Q(bit_ctr[27]), .C(clk16MHz), .E(n7792), 
            .D(n133[27]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i28 (.Q(bit_ctr[28]), .C(clk16MHz), .E(n7792), 
            .D(n133[28]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i29 (.Q(bit_ctr[29]), .C(clk16MHz), .E(n7792), 
            .D(n133[29]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2281__i30 (.Q(bit_ctr[30]), .C(clk16MHz), .E(n7792), 
            .D(n133[30]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_2281__i31 (.Q(bit_ctr[31]), .C(clk16MHz), .E(n7792), 
            .D(n133[31]), .R(n29101));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 i37244_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n53036));
    defparam i37244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37245_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n53037));
    defparam i37245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37236_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n53028));
    defparam i37236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37235_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n53027));
    defparam i37235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(n36592), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n51143));
    defparam i1_4_lut.LUT_INIT = 16'hf5fd;
    SB_LUT4 i1_4_lut_adj_1721 (.I0(n51143), .I1(n23_adj_5419), .I2(\state[1] ), 
            .I3(n27272), .O(n28689));
    defparam i1_4_lut_adj_1721.LUT_INIT = 16'ha0a8;
    SB_LUT4 i39404_3_lut (.I0(n56371), .I1(n56635), .I2(color_bit_N_833[2]), 
            .I3(GND_net), .O(n55197));
    defparam i39404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[4]), .I1(bit_ctr[3]), .I2(n36459), .I3(GND_net), 
            .O(n45504));
    defparam i1_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i39466_4_lut (.I0(n55197), .I1(n56515), .I2(bit_ctr[3]), .I3(n36459), 
            .O(n55259));   // verilog/neopixel.v(22[26:38])
    defparam i39466_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i38623_3_lut (.I0(n56467), .I1(bit_ctr[3]), .I2(n36459), .I3(GND_net), 
            .O(n54304));
    defparam i38623_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i21666_4_lut (.I0(n54304), .I1(\state_3__N_639[1] ), .I2(n55259), 
            .I3(n45504), .O(state_3__N_639[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i21666_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n56368_bdd_4_lut_4_lut (.I0(color_bit_N_833[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n56368), .O(n56371));   // verilog/neopixel.v(19[6:15])
    defparam n56368_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    SB_DFF timer_2280__i31 (.Q(timer[31]), .C(clk16MHz), .D(n133_adj_5456[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i30 (.Q(timer[30]), .C(clk16MHz), .D(n133_adj_5456[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i29 (.Q(timer[29]), .C(clk16MHz), .D(n133_adj_5456[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i28 (.Q(timer[28]), .C(clk16MHz), .D(n133_adj_5456[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i27 (.Q(timer[27]), .C(clk16MHz), .D(n133_adj_5456[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i26 (.Q(timer[26]), .C(clk16MHz), .D(n133_adj_5456[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i25 (.Q(timer[25]), .C(clk16MHz), .D(n133_adj_5456[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i24 (.Q(timer[24]), .C(clk16MHz), .D(n133_adj_5456[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i23 (.Q(timer[23]), .C(clk16MHz), .D(n133_adj_5456[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i22 (.Q(timer[22]), .C(clk16MHz), .D(n133_adj_5456[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i21 (.Q(timer[21]), .C(clk16MHz), .D(n133_adj_5456[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i20 (.Q(timer[20]), .C(clk16MHz), .D(n133_adj_5456[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i19 (.Q(timer[19]), .C(clk16MHz), .D(n133_adj_5456[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i18 (.Q(timer[18]), .C(clk16MHz), .D(n133_adj_5456[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i17 (.Q(timer[17]), .C(clk16MHz), .D(n133_adj_5456[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i16 (.Q(timer[16]), .C(clk16MHz), .D(n133_adj_5456[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i15 (.Q(timer[15]), .C(clk16MHz), .D(n133_adj_5456[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i14 (.Q(timer[14]), .C(clk16MHz), .D(n133_adj_5456[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i13 (.Q(timer[13]), .C(clk16MHz), .D(n133_adj_5456[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i12 (.Q(timer[12]), .C(clk16MHz), .D(n133_adj_5456[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i11 (.Q(timer[11]), .C(clk16MHz), .D(n133_adj_5456[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i10 (.Q(timer[10]), .C(clk16MHz), .D(n133_adj_5456[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i9 (.Q(timer[9]), .C(clk16MHz), .D(n133_adj_5456[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i8 (.Q(timer[8]), .C(clk16MHz), .D(n133_adj_5456[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i7 (.Q(timer[7]), .C(clk16MHz), .D(n133_adj_5456[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i6 (.Q(timer[6]), .C(clk16MHz), .D(n133_adj_5456[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i5 (.Q(timer[5]), .C(clk16MHz), .D(n133_adj_5456[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i4 (.Q(timer[4]), .C(clk16MHz), .D(n133_adj_5456[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i3 (.Q(timer[3]), .C(clk16MHz), .D(n133_adj_5456[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i2 (.Q(timer[2]), .C(clk16MHz), .D(n133_adj_5456[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2280__i1 (.Q(timer[1]), .C(clk16MHz), .D(n133_adj_5456[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 color_bit_N_833_1__bdd_4_lut (.I0(color_bit_N_833[1]), .I1(n52931), 
            .I2(n52932), .I3(color_bit_N_833[2]), .O(n56512));
    defparam color_bit_N_833_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n56512_bdd_4_lut (.I0(n56512), .I1(n52926), .I2(n52925), .I3(color_bit_N_833[2]), 
            .O(n56515));
    defparam n56512_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2281_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[31]), 
            .I3(n44055), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_2281_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[30]), 
            .I3(n44054), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_32 (.CI(n44054), .I0(GND_net), .I1(bit_ctr[30]), 
            .CO(n44055));
    SB_LUT4 bit_ctr_2281_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[29]), 
            .I3(n44053), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_31 (.CI(n44053), .I0(GND_net), .I1(bit_ctr[29]), 
            .CO(n44054));
    SB_LUT4 bit_ctr_2281_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[28]), 
            .I3(n44052), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_30 (.CI(n44052), .I0(GND_net), .I1(bit_ctr[28]), 
            .CO(n44053));
    SB_LUT4 bit_ctr_2281_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[27]), 
            .I3(n44051), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_33_lut (.I0(n52408), .I1(timer[31]), .I2(n1[31]), 
            .I3(n43155), .O(n27276)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_CARRY bit_ctr_2281_add_4_29 (.CI(n44051), .I0(GND_net), .I1(bit_ctr[27]), 
            .CO(n44052));
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2281_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[26]), 
            .I3(n44050), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_28 (.CI(n44050), .I0(GND_net), .I1(bit_ctr[26]), 
            .CO(n44051));
    SB_LUT4 bit_ctr_2281_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[25]), 
            .I3(n44049), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n52406), .I1(timer[30]), .I2(n1[30]), 
            .I3(n43154), .O(n52408)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY bit_ctr_2281_add_4_27 (.CI(n44049), .I0(GND_net), .I1(bit_ctr[25]), 
            .CO(n44050));
    SB_LUT4 bit_ctr_2281_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[24]), 
            .I3(n44048), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_26 (.CI(n44048), .I0(GND_net), .I1(bit_ctr[24]), 
            .CO(n44049));
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_32 (.CI(n43154), .I0(timer[30]), .I1(n1[30]), 
            .CO(n43155));
    SB_LUT4 bit_ctr_2281_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[23]), 
            .I3(n44047), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_25 (.CI(n44047), .I0(GND_net), .I1(bit_ctr[23]), 
            .CO(n44048));
    SB_LUT4 sub_14_add_2_31_lut (.I0(n52404), .I1(timer[29]), .I2(n1[29]), 
            .I3(n43153), .O(n52406)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2281_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[22]), 
            .I3(n44046), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_24 (.CI(n44046), .I0(GND_net), .I1(bit_ctr[22]), 
            .CO(n44047));
    SB_LUT4 bit_ctr_2281_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[21]), 
            .I3(n44045), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_23 (.CI(n44045), .I0(GND_net), .I1(bit_ctr[21]), 
            .CO(n44046));
    SB_CARRY sub_14_add_2_31 (.CI(n43153), .I0(timer[29]), .I1(n1[29]), 
            .CO(n43154));
    SB_LUT4 bit_ctr_2281_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[20]), 
            .I3(n44044), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_22 (.CI(n44044), .I0(GND_net), .I1(bit_ctr[20]), 
            .CO(n44045));
    SB_LUT4 sub_14_add_2_30_lut (.I0(n52402), .I1(timer[28]), .I2(n1[28]), 
            .I3(n43152), .O(n52404)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_2281_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[19]), 
            .I3(n44043), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY bit_ctr_2281_add_4_21 (.CI(n44043), .I0(GND_net), .I1(bit_ctr[19]), 
            .CO(n44044));
    SB_LUT4 bit_ctr_2281_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[18]), 
            .I3(n44042), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_20 (.CI(n44042), .I0(GND_net), .I1(bit_ctr[18]), 
            .CO(n44043));
    SB_CARRY sub_14_add_2_30 (.CI(n43152), .I0(timer[28]), .I1(n1[28]), 
            .CO(n43153));
    SB_DFF timer_2280__i0 (.Q(timer[0]), .C(clk16MHz), .D(n133_adj_5456[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 bit_ctr_2281_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[17]), 
            .I3(n44041), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_29_lut (.I0(n52400), .I1(timer[27]), .I2(n1[27]), 
            .I3(n43151), .O(n52402)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n43151), .I0(timer[27]), .I1(n1[27]), 
            .CO(n43152));
    SB_CARRY bit_ctr_2281_add_4_19 (.CI(n44041), .I0(GND_net), .I1(bit_ctr[17]), 
            .CO(n44042));
    SB_LUT4 sub_14_add_2_28_lut (.I0(n52398), .I1(timer[26]), .I2(n1[26]), 
            .I3(n43150), .O(n52400)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_2281_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[16]), 
            .I3(n44040), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_18 (.CI(n44040), .I0(GND_net), .I1(bit_ctr[16]), 
            .CO(n44041));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk16MHz), .E(n28689), .D(state_3__N_639[0]), 
            .S(n29076));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 color_bit_N_833_1__bdd_4_lut_40680 (.I0(color_bit_N_833[1]), .I1(n53027), 
            .I2(n53028), .I3(color_bit_N_833[2]), .O(n56464));
    defparam color_bit_N_833_1__bdd_4_lut_40680.LUT_INIT = 16'he4aa;
    SB_LUT4 n56464_bdd_4_lut (.I0(n56464), .I1(n53037), .I2(n53036), .I3(color_bit_N_833[2]), 
            .O(n56467));
    defparam n56464_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2281_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[15]), 
            .I3(n44039), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_17 (.CI(n44039), .I0(GND_net), .I1(bit_ctr[15]), 
            .CO(n44040));
    SB_LUT4 bit_ctr_2281_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[14]), 
            .I3(n44038), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_16 (.CI(n44038), .I0(GND_net), .I1(bit_ctr[14]), 
            .CO(n44039));
    SB_CARRY sub_14_add_2_28 (.CI(n43150), .I0(timer[26]), .I1(n1[26]), 
            .CO(n43151));
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2281_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[13]), 
            .I3(n44037), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_4_lut (.I0(n49519), .I1(n44914), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n49641));
    defparam i22_4_lut.LUT_INIT = 16'hacca;
    SB_CARRY bit_ctr_2281_add_4_15 (.CI(n44037), .I0(GND_net), .I1(bit_ctr[13]), 
            .CO(n44038));
    SB_LUT4 i33859_4_lut (.I0(n49641), .I1(\state[1] ), .I2(n27135), .I3(start), 
            .O(n49594));
    defparam i33859_4_lut.LUT_INIT = 16'hcccd;
    SB_LUT4 sub_14_add_2_27_lut (.I0(n52396), .I1(timer[25]), .I2(n1[25]), 
            .I3(n43149), .O(n52398)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_2281_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[12]), 
            .I3(n44036), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_14 (.CI(n44036), .I0(GND_net), .I1(bit_ctr[12]), 
            .CO(n44037));
    SB_LUT4 bit_ctr_2281_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[11]), 
            .I3(n44035), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_13 (.CI(n44035), .I0(GND_net), .I1(bit_ctr[11]), 
            .CO(n44036));
    SB_LUT4 bit_ctr_2281_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[10]), 
            .I3(n44034), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_12 (.CI(n44034), .I0(GND_net), .I1(bit_ctr[10]), 
            .CO(n44035));
    SB_LUT4 bit_ctr_2281_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[9]), 
            .I3(n44033), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_11 (.CI(n44033), .I0(GND_net), .I1(bit_ctr[9]), 
            .CO(n44034));
    SB_LUT4 bit_ctr_2281_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[8]), 
            .I3(n44032), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_10 (.CI(n44032), .I0(GND_net), .I1(bit_ctr[8]), 
            .CO(n44033));
    SB_LUT4 bit_ctr_2281_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[7]), 
            .I3(n44031), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_9 (.CI(n44031), .I0(GND_net), .I1(bit_ctr[7]), 
            .CO(n44032));
    SB_LUT4 bit_ctr_2281_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[6]), 
            .I3(n44030), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_8 (.CI(n44030), .I0(GND_net), .I1(bit_ctr[6]), 
            .CO(n44031));
    SB_LUT4 bit_ctr_2281_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[5]), 
            .I3(n44029), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_7 (.CI(n44029), .I0(GND_net), .I1(bit_ctr[5]), 
            .CO(n44030));
    SB_CARRY sub_14_add_2_27 (.CI(n43149), .I0(timer[25]), .I1(n1[25]), 
            .CO(n43150));
    SB_LUT4 bit_ctr_2281_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[4]), 
            .I3(n44028), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_6 (.CI(n44028), .I0(GND_net), .I1(bit_ctr[4]), 
            .CO(n44029));
    SB_LUT4 bit_ctr_2281_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[3]), 
            .I3(n44027), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_5 (.CI(n44027), .I0(GND_net), .I1(bit_ctr[3]), 
            .CO(n44028));
    SB_LUT4 bit_ctr_2281_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[2]), 
            .I3(n44026), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_26_lut (.I0(n52394), .I1(timer[24]), .I2(n1[24]), 
            .I3(n43148), .O(n52396)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_26 (.CI(n43148), .I0(timer[24]), .I1(n1[24]), 
            .CO(n43149));
    SB_CARRY bit_ctr_2281_add_4_4 (.CI(n44026), .I0(GND_net), .I1(bit_ctr[2]), 
            .CO(n44027));
    SB_LUT4 sub_14_add_2_25_lut (.I0(n52392), .I1(timer[23]), .I2(n1[23]), 
            .I3(n43147), .O(n52394)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_2281_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[1]), 
            .I3(n44025), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_3 (.CI(n44025), .I0(GND_net), .I1(bit_ctr[1]), 
            .CO(n44026));
    SB_LUT4 bit_ctr_2281_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2281_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2281_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_ctr[0]), 
            .CO(n44025));
    SB_LUT4 timer_2280_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n44024), .O(n133_adj_5456[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2280_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n44023), .O(n133_adj_5456[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_32 (.CI(n44023), .I0(GND_net), .I1(timer[30]), 
            .CO(n44024));
    SB_LUT4 timer_2280_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n44022), .O(n133_adj_5456[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_31 (.CI(n44022), .I0(GND_net), .I1(timer[29]), 
            .CO(n44023));
    SB_CARRY sub_14_add_2_25 (.CI(n43147), .I0(timer[23]), .I1(n1[23]), 
            .CO(n43148));
    SB_LUT4 sub_14_add_2_24_lut (.I0(n52390), .I1(timer[22]), .I2(n1[22]), 
            .I3(n43146), .O(n52392)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 timer_2280_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n44021), .O(n133_adj_5456[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_30 (.CI(n44021), .I0(GND_net), .I1(timer[28]), 
            .CO(n44022));
    SB_CARRY sub_14_add_2_24 (.CI(n43146), .I0(timer[22]), .I1(n1[22]), 
            .CO(n43147));
    SB_LUT4 timer_2280_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n44020), .O(n133_adj_5456[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_23_lut (.I0(n52388), .I1(timer[21]), .I2(n1[21]), 
            .I3(n43145), .O(n52390)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY timer_2280_add_4_29 (.CI(n44020), .I0(GND_net), .I1(timer[27]), 
            .CO(n44021));
    SB_LUT4 timer_2280_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n44019), .O(n133_adj_5456[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_28 (.CI(n44019), .I0(GND_net), .I1(timer[26]), 
            .CO(n44020));
    SB_LUT4 timer_2280_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n44018), .O(n133_adj_5456[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_27 (.CI(n44018), .I0(GND_net), .I1(timer[25]), 
            .CO(n44019));
    SB_LUT4 timer_2280_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n44017), .O(n133_adj_5456[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_23 (.CI(n43145), .I0(timer[21]), .I1(n1[21]), 
            .CO(n43146));
    SB_LUT4 sub_14_add_2_22_lut (.I0(n52386), .I1(timer[20]), .I2(n1[20]), 
            .I3(n43144), .O(n52388)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY timer_2280_add_4_26 (.CI(n44017), .I0(GND_net), .I1(timer[24]), 
            .CO(n44018));
    SB_LUT4 timer_2280_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n44016), .O(n133_adj_5456[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_25 (.CI(n44016), .I0(GND_net), .I1(timer[23]), 
            .CO(n44017));
    SB_LUT4 timer_2280_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n44015), .O(n133_adj_5456[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37133_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n52925));
    defparam i37133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37134_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n52926));
    defparam i37134_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2280_add_4_24 (.CI(n44015), .I0(GND_net), .I1(timer[22]), 
            .CO(n44016));
    SB_LUT4 timer_2280_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n44014), .O(n133_adj_5456[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_22 (.CI(n43144), .I0(timer[20]), .I1(n1[20]), 
            .CO(n43145));
    SB_CARRY timer_2280_add_4_23 (.CI(n44014), .I0(GND_net), .I1(timer[21]), 
            .CO(n44015));
    SB_LUT4 i37140_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n52932));
    defparam i37140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37139_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n52931));
    defparam i37139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2280_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n44013), .O(n133_adj_5456[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_21_lut (.I0(n52384), .I1(timer[19]), .I2(n1[19]), 
            .I3(n43143), .O(n52386)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_833[1]));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY timer_2280_add_4_22 (.CI(n44013), .I0(GND_net), .I1(timer[20]), 
            .CO(n44014));
    SB_LUT4 timer_2280_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n44012), .O(n133_adj_5456[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_21 (.CI(n44012), .I0(GND_net), .I1(timer[19]), 
            .CO(n44013));
    SB_CARRY sub_14_add_2_21 (.CI(n43143), .I0(timer[19]), .I1(n1[19]), 
            .CO(n43144));
    SB_LUT4 timer_2280_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n44011), .O(n133_adj_5456[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_20 (.CI(n44011), .I0(GND_net), .I1(timer[18]), 
            .CO(n44012));
    SB_LUT4 i14958_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n29033));   // verilog/neopixel.v(36[4] 116[11])
    defparam i14958_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 timer_2280_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n44010), .O(n133_adj_5456[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_19 (.CI(n44010), .I0(GND_net), .I1(timer[17]), 
            .CO(n44011));
    SB_LUT4 sub_14_add_2_20_lut (.I0(n52382), .I1(timer[18]), .I2(n1[18]), 
            .I3(n43142), .O(n52384)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 timer_2280_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n44009), .O(n133_adj_5456[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_18 (.CI(n44009), .I0(GND_net), .I1(timer[16]), 
            .CO(n44010));
    SB_LUT4 timer_2280_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n44008), .O(n133_adj_5456[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_17 (.CI(n44008), .I0(GND_net), .I1(timer[15]), 
            .CO(n44009));
    SB_LUT4 timer_2280_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n44007), .O(n133_adj_5456[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_16 (.CI(n44007), .I0(GND_net), .I1(timer[14]), 
            .CO(n44008));
    SB_LUT4 timer_2280_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n44006), .O(n133_adj_5456[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_15 (.CI(n44006), .I0(GND_net), .I1(timer[13]), 
            .CO(n44007));
    SB_LUT4 i19_4_lut (.I0(bit_ctr[23]), .I1(bit_ctr[16]), .I2(bit_ctr[20]), 
            .I3(bit_ctr[7]), .O(n46));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_2280_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n44005), .O(n133_adj_5456[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_14 (.CI(n44005), .I0(GND_net), .I1(timer[12]), 
            .CO(n44006));
    SB_LUT4 timer_2280_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n44004), .O(n133_adj_5456[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_13 (.CI(n44004), .I0(GND_net), .I1(timer[11]), 
            .CO(n44005));
    SB_LUT4 timer_2280_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n44003), .O(n133_adj_5456[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_12 (.CI(n44003), .I0(GND_net), .I1(timer[10]), 
            .CO(n44004));
    SB_LUT4 timer_2280_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n44002), .O(n133_adj_5456[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut (.I0(bit_ctr[14]), .I1(bit_ctr[9]), .I2(bit_ctr[25]), 
            .I3(bit_ctr[10]), .O(n44));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_2280_add_4_11 (.CI(n44002), .I0(GND_net), .I1(timer[9]), 
            .CO(n44003));
    SB_LUT4 timer_2280_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n44001), .O(n133_adj_5456[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18_4_lut (.I0(bit_ctr[27]), .I1(bit_ctr[12]), .I2(bit_ctr[15]), 
            .I3(bit_ctr[29]), .O(n45));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_2280_add_4_10 (.CI(n44001), .I0(GND_net), .I1(timer[8]), 
            .CO(n44002));
    SB_LUT4 timer_2280_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n44000), .O(n133_adj_5456[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n43142), .I0(timer[18]), .I1(n1[18]), 
            .CO(n43143));
    SB_CARRY timer_2280_add_4_9 (.CI(n44000), .I0(GND_net), .I1(timer[7]), 
            .CO(n44001));
    SB_LUT4 timer_2280_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n43999), .O(n133_adj_5456[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut (.I0(bit_ctr[6]), .I1(bit_ctr[31]), .I2(bit_ctr[19]), 
            .I3(bit_ctr[21]), .O(n43));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_2280_add_4_8 (.CI(n43999), .I0(GND_net), .I1(timer[6]), 
            .CO(n44000));
    SB_LUT4 timer_2280_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n43998), .O(n133_adj_5456[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_7 (.CI(n43998), .I0(GND_net), .I1(timer[5]), 
            .CO(n43999));
    SB_LUT4 timer_2280_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n43997), .O(n133_adj_5456[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_6 (.CI(n43997), .I0(GND_net), .I1(timer[4]), 
            .CO(n43998));
    SB_LUT4 timer_2280_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n43996), .O(n133_adj_5456[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut (.I0(bit_ctr[17]), .I1(bit_ctr[28]), .I2(bit_ctr[11]), 
            .I3(bit_ctr[5]), .O(n42));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_2280_add_4_5 (.CI(n43996), .I0(GND_net), .I1(timer[3]), 
            .CO(n43997));
    SB_LUT4 timer_2280_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n43995), .O(n133_adj_5456[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_4 (.CI(n43995), .I0(GND_net), .I1(timer[2]), 
            .CO(n43996));
    SB_LUT4 timer_2280_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n43994), .O(n133_adj_5456[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_3 (.CI(n43994), .I0(GND_net), .I1(timer[1]), 
            .CO(n43995));
    SB_LUT4 timer_2280_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133_adj_5456[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2280_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2280_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n43994));
    SB_LUT4 i13_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(GND_net), .O(n40));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 sub_14_add_2_19_lut (.I0(n52380), .I1(timer[17]), .I2(n1[17]), 
            .I3(n43141), .O(n52382)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i21_4_lut (.I0(bit_ctr[26]), .I1(n42), .I2(bit_ctr[13]), .I3(bit_ctr[22]), 
            .O(n48));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n43), .I1(n45), .I2(n44), .I3(n46), .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(bit_ctr[30]), .I1(n48), .I2(n40), .I3(bit_ctr[24]), 
            .O(n51));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_19 (.CI(n43141), .I0(timer[17]), .I1(n1[17]), 
            .CO(n43142));
    SB_LUT4 i1_4_lut_adj_1722 (.I0(bit_ctr[3]), .I1(n51), .I2(bit_ctr[4]), 
            .I3(n52), .O(\state_3__N_639[1] ));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'hffec;
    SB_LUT4 i1_2_lut_adj_1723 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n27272));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_2_lut_adj_1723.LUT_INIT = 16'hbbbb;
    SB_LUT4 i547_2_lut (.I0(LED_c), .I1(\state_3__N_639[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n2586));   // verilog/neopixel.v(40[18] 45[12])
    defparam i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4695_4_lut (.I0(n10_adj_5453), .I1(n2586), .I2(\state[1] ), 
            .I3(n27272), .O(n7747));
    defparam i4695_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i3_4_lut (.I0(n7792), .I1(n7747), .I2(n2586), .I3(n29033), 
            .O(n29101));
    defparam i3_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i26_4_lut (.I0(n27272), .I1(n54239), .I2(\state[1] ), .I3(n23_adj_5419), 
            .O(n7792));
    defparam i26_4_lut.LUT_INIT = 16'hc5c0;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk16MHz), .D(n29258));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_18_lut (.I0(n52378), .I1(timer[16]), .I2(n1[16]), 
            .I3(n43140), .O(n52380)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_18 (.CI(n43140), .I0(timer[16]), .I1(n1[16]), 
            .CO(n43141));
    SB_LUT4 sub_14_add_2_17_lut (.I0(n52376), .I1(timer[15]), .I2(n1[15]), 
            .I3(n43139), .O(n52378)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_17 (.CI(n43139), .I0(timer[15]), .I1(n1[15]), 
            .CO(n43140));
    SB_LUT4 sub_14_add_2_16_lut (.I0(n52374), .I1(timer[14]), .I2(n1[14]), 
            .I3(n43138), .O(n52376)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_16 (.CI(n43138), .I0(timer[14]), .I1(n1[14]), 
            .CO(n43139));
    SB_LUT4 sub_14_add_2_15_lut (.I0(n52372), .I1(timer[13]), .I2(n1[13]), 
            .I3(n43137), .O(n52374)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_15 (.CI(n43137), .I0(timer[13]), .I1(n1[13]), 
            .CO(n43138));
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_790[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n43136), .O(n52372)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_14 (.CI(n43136), .I0(timer[12]), .I1(n1[12]), 
            .CO(n43137));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n43135), .O(one_wire_N_790[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n43135), .I0(timer[11]), .I1(n1[11]), 
            .CO(n43136));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n43134), .O(one_wire_N_790[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n43134), .I0(timer[10]), .I1(n1[10]), 
            .CO(n43135));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n43133), .O(one_wire_N_790[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n43133), .I0(timer[9]), .I1(n1[9]), 
            .CO(n43134));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n43132), .O(one_wire_N_790[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n43132), .I0(timer[8]), .I1(n1[8]), 
            .CO(n43133));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n43131), .O(one_wire_N_790[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n43131), .I0(timer[7]), .I1(n1[7]), .CO(n43132));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n43130), .O(one_wire_N_790[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n43130), .I0(timer[6]), .I1(n1[6]), .CO(n43131));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n43129), .O(one_wire_N_790[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n43129), .I0(timer[5]), .I1(n1[5]), .CO(n43130));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n43128), .O(one_wire_N_790[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n43128), .I0(timer[4]), .I1(n1[4]), .CO(n43129));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n43127), .O(one_wire_N_790[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n43127), .I0(timer[3]), .I1(n1[3]), .CO(n43128));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n43126), .O(one_wire_N_790[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n43126), .I0(timer[2]), .I1(n1[2]), .CO(n43127));
    SB_LUT4 sub_14_add_2_3_lut (.I0(GND_net), .I1(timer[1]), .I2(n1[1]), 
            .I3(n43125), .O(one_wire_N_790[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_3 (.CI(n43125), .I0(timer[1]), .I1(n1[1]), .CO(n43126));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n43125));
    SB_LUT4 i38586_3_lut_4_lut (.I0(n27135), .I1(n54378), .I2(start), 
            .I3(\state[1] ), .O(n54379));
    defparam i38586_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i38724_2_lut_3_lut (.I0(one_wire_N_790[3]), .I1(one_wire_N_790[2]), 
            .I2(start), .I3(GND_net), .O(n54236));
    defparam i38724_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n36592), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n51217));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk16MHz), .D(n29700));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk16MHz), .D(n29699));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk16MHz), .D(n29698));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk16MHz), .D(n29697));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk16MHz), .D(n29696));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk16MHz), .D(n29695));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk16MHz), .D(n29694));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk16MHz), .D(n29693));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk16MHz), .D(n29692));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk16MHz), .D(n29691));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk16MHz), .D(n29690));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk16MHz), .D(n29689));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk16MHz), .D(n29688));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk16MHz), .D(n29684));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk16MHz), .D(n29683));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk16MHz), .D(n29682));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk16MHz), .D(n29681));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk16MHz), .D(n29680));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk16MHz), .D(n29679));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk16MHz), .D(n29678));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk16MHz), .D(n29677));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk16MHz), .D(n29676));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk16MHz), .D(n29675));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk16MHz), .D(n29674));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk16MHz), .D(n29673));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk16MHz), .D(n29672));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk16MHz), .D(n29671));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk16MHz), .D(n29670));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk16MHz), .D(n29669));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk16MHz), .D(n29668));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk16MHz), .D(n29667));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n56632));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk16MHz), .E(n49637), .D(\neo_pixel_transmitter.done_N_853 ), 
            .R(n51217));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk16MHz), .E(VCC_net), .D(n29436));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22397_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(n36459));
    defparam i22397_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(color_bit_N_833[2]));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1e1e;
    SB_LUT4 i38602_2_lut_3_lut (.I0(LED_c), .I1(\state_3__N_639[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n54239));
    defparam i38602_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_2_lut_3_lut (.I0(n27135), .I1(one_wire_N_790[3]), .I2(one_wire_N_790[2]), 
            .I3(GND_net), .O(n10_adj_5453));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i22526_4_lut (.I0(one_wire_N_790[8]), .I1(n27276), .I2(one_wire_N_790[10]), 
            .I3(one_wire_N_790[9]), .O(n36592));
    defparam i22526_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i33789_2_lut (.I0(one_wire_N_790[3]), .I1(one_wire_N_790[2]), 
            .I2(GND_net), .I3(GND_net), .O(n49519));
    defparam i33789_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(one_wire_N_790[3]), .I1(one_wire_N_790[2]), .I2(one_wire_N_790[1]), 
            .I3(GND_net), .O(n44914));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1724 (.I0(one_wire_N_790[5]), .I1(one_wire_N_790[4]), 
            .I2(GND_net), .I3(GND_net), .O(n52410));   // verilog/neopixel.v(62[15:42])
    defparam i1_2_lut_adj_1724.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(one_wire_N_790[8]), .I1(one_wire_N_790[7]), 
            .I2(one_wire_N_790[6]), .I3(n52410), .O(n52416));   // verilog/neopixel.v(62[15:42])
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(one_wire_N_790[10]), .I1(n27276), .I2(one_wire_N_790[9]), 
            .I3(n52416), .O(n27135));   // verilog/neopixel.v(62[15:42])
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 i33851_4_lut (.I0(n27135), .I1(n44914), .I2(n49519), .I3(\state[0] ), 
            .O(n23_adj_5419));
    defparam i33851_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i38712_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n54242));
    defparam i38712_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i33731_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n23_adj_5419), .I3(GND_net), .O(n49458));
    defparam i33731_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1727 (.I0(n49458), .I1(n54242), .I2(\state[1] ), 
            .I3(n36592), .O(n7));
    defparam i15_4_lut_adj_1727.LUT_INIT = 16'h3a0a;
    SB_LUT4 i40435_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(start_N_838));   // verilog/neopixel.v(36[4] 116[11])
    defparam i40435_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i33785_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n49515));
    defparam i33785_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39784_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n48656));
    defparam i39784_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1728 (.I0(one_wire_N_790[2]), .I1(n48656), .I2(one_wire_N_790[3]), 
            .I3(one_wire_N_790[1]), .O(n103));
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'h4dcd;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_790[7]), .I1(one_wire_N_790[9]), .I2(n49515), 
            .I3(n103), .O(n16_adj_5454));
    defparam i6_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(one_wire_N_790[8]), .I1(one_wire_N_790[4]), 
            .I2(n16_adj_5454), .I3(n27276), .O(n6_adj_5455));
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut (.I0(one_wire_N_790[10]), .I1(one_wire_N_790[6]), .I2(one_wire_N_790[5]), 
            .I3(n6_adj_5455), .O(n56661));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1370_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_847 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_1370_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n56632_bdd_4_lut (.I0(n56632), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_833[1]), .O(n56635));
    defparam n56632_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38974_4_lut (.I0(n44914), .I1(n49519), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n54378));
    defparam i38974_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53_4_lut (.I0(n54236), .I1(n36592), .I2(\state[1] ), .I3(n27135), 
            .O(n49617));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n49617), .I1(n54379), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n49637));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_853 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_0__bdd_4_lut_40779_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n56368));   // verilog/neopixel.v(19[6:15])
    defparam bit_ctr_0__bdd_4_lut_40779_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15000_2_lut_3_lut (.I0(n28689), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(GND_net), .O(n29076));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15000_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1)_U0 
//

module \quadrature_decoder(1)_U0  (b_prev, n2269, GND_net, a_new, position_31__N_4108, 
            ENCODER0_B_N_keep, ENCODER0_A_N_keep, n29393, n2233, encoder0_position, 
            VCC_net) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input n2269;
    input GND_net;
    output [1:0]a_new;
    output position_31__N_4108;
    input ENCODER0_B_N_keep;
    input ENCODER0_A_N_keep;
    input n29393;
    output n2233;
    output [31:0]encoder0_position;
    input VCC_net;
    
    
    wire n29427;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire position_31__N_4111, debounce_cnt, a_prev, direction_N_4113;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_4116, n29412;
    wire [31:0]n133;
    
    wire n44140, n44139, n44138, n44137, n44136, n44135, n44134, 
        n44133, n44132, n44131, n44130, n44129, n44128, n44127, 
        n44126, n44125, n44124, n44123, n44122, n44121, n44120, 
        n44119, n44118, n44117, n44116, n44115, n44114, n44113, 
        n44112, n44111, n44110;
    
    SB_DFF b_prev_39 (.Q(b_prev), .C(n2269), .D(n29427));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_4111));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_4111), 
            .I3(a_new[1]), .O(position_31__N_4108));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_4113));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n2269), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n2269), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n2269), .D(a_prev_N_4116));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_38 (.Q(a_prev), .C(n2269), .D(n29412));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n2233), .C(n2269), .D(n29393));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2284_add_4_33_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[31]), .I3(n44140), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2284_add_4_32_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[30]), .I3(n44139), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_32 (.CI(n44139), .I0(direction_N_4113), 
            .I1(encoder0_position[30]), .CO(n44140));
    SB_LUT4 position_2284_add_4_31_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[29]), .I3(n44138), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_31 (.CI(n44138), .I0(direction_N_4113), 
            .I1(encoder0_position[29]), .CO(n44139));
    SB_LUT4 position_2284_add_4_30_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[28]), .I3(n44137), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_30 (.CI(n44137), .I0(direction_N_4113), 
            .I1(encoder0_position[28]), .CO(n44138));
    SB_LUT4 position_2284_add_4_29_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[27]), .I3(n44136), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_29 (.CI(n44136), .I0(direction_N_4113), 
            .I1(encoder0_position[27]), .CO(n44137));
    SB_LUT4 position_2284_add_4_28_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[26]), .I3(n44135), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_28 (.CI(n44135), .I0(direction_N_4113), 
            .I1(encoder0_position[26]), .CO(n44136));
    SB_LUT4 position_2284_add_4_27_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[25]), .I3(n44134), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_27 (.CI(n44134), .I0(direction_N_4113), 
            .I1(encoder0_position[25]), .CO(n44135));
    SB_LUT4 position_2284_add_4_26_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[24]), .I3(n44133), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_26 (.CI(n44133), .I0(direction_N_4113), 
            .I1(encoder0_position[24]), .CO(n44134));
    SB_LUT4 position_2284_add_4_25_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[23]), .I3(n44132), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_25 (.CI(n44132), .I0(direction_N_4113), 
            .I1(encoder0_position[23]), .CO(n44133));
    SB_LUT4 position_2284_add_4_24_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[22]), .I3(n44131), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_24 (.CI(n44131), .I0(direction_N_4113), 
            .I1(encoder0_position[22]), .CO(n44132));
    SB_LUT4 position_2284_add_4_23_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[21]), .I3(n44130), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_23 (.CI(n44130), .I0(direction_N_4113), 
            .I1(encoder0_position[21]), .CO(n44131));
    SB_LUT4 position_2284_add_4_22_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[20]), .I3(n44129), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_22 (.CI(n44129), .I0(direction_N_4113), 
            .I1(encoder0_position[20]), .CO(n44130));
    SB_LUT4 position_2284_add_4_21_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[19]), .I3(n44128), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_21 (.CI(n44128), .I0(direction_N_4113), 
            .I1(encoder0_position[19]), .CO(n44129));
    SB_LUT4 position_2284_add_4_20_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[18]), .I3(n44127), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_20 (.CI(n44127), .I0(direction_N_4113), 
            .I1(encoder0_position[18]), .CO(n44128));
    SB_LUT4 position_2284_add_4_19_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[17]), .I3(n44126), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_19 (.CI(n44126), .I0(direction_N_4113), 
            .I1(encoder0_position[17]), .CO(n44127));
    SB_LUT4 position_2284_add_4_18_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[16]), .I3(n44125), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_18 (.CI(n44125), .I0(direction_N_4113), 
            .I1(encoder0_position[16]), .CO(n44126));
    SB_LUT4 position_2284_add_4_17_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[15]), .I3(n44124), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_17 (.CI(n44124), .I0(direction_N_4113), 
            .I1(encoder0_position[15]), .CO(n44125));
    SB_LUT4 position_2284_add_4_16_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[14]), .I3(n44123), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_16 (.CI(n44123), .I0(direction_N_4113), 
            .I1(encoder0_position[14]), .CO(n44124));
    SB_LUT4 position_2284_add_4_15_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[13]), .I3(n44122), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_15 (.CI(n44122), .I0(direction_N_4113), 
            .I1(encoder0_position[13]), .CO(n44123));
    SB_LUT4 position_2284_add_4_14_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[12]), .I3(n44121), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_14 (.CI(n44121), .I0(direction_N_4113), 
            .I1(encoder0_position[12]), .CO(n44122));
    SB_LUT4 position_2284_add_4_13_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[11]), .I3(n44120), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_13 (.CI(n44120), .I0(direction_N_4113), 
            .I1(encoder0_position[11]), .CO(n44121));
    SB_LUT4 position_2284_add_4_12_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[10]), .I3(n44119), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_12 (.CI(n44119), .I0(direction_N_4113), 
            .I1(encoder0_position[10]), .CO(n44120));
    SB_LUT4 position_2284_add_4_11_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[9]), .I3(n44118), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_11 (.CI(n44118), .I0(direction_N_4113), 
            .I1(encoder0_position[9]), .CO(n44119));
    SB_LUT4 position_2284_add_4_10_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[8]), .I3(n44117), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_10 (.CI(n44117), .I0(direction_N_4113), 
            .I1(encoder0_position[8]), .CO(n44118));
    SB_LUT4 position_2284_add_4_9_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[7]), .I3(n44116), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_9 (.CI(n44116), .I0(direction_N_4113), 
            .I1(encoder0_position[7]), .CO(n44117));
    SB_LUT4 position_2284_add_4_8_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[6]), .I3(n44115), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_8 (.CI(n44115), .I0(direction_N_4113), 
            .I1(encoder0_position[6]), .CO(n44116));
    SB_LUT4 position_2284_add_4_7_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[5]), .I3(n44114), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_7 (.CI(n44114), .I0(direction_N_4113), 
            .I1(encoder0_position[5]), .CO(n44115));
    SB_LUT4 position_2284_add_4_6_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[4]), .I3(n44113), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_6 (.CI(n44113), .I0(direction_N_4113), 
            .I1(encoder0_position[4]), .CO(n44114));
    SB_LUT4 position_2284_add_4_5_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[3]), .I3(n44112), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_5 (.CI(n44112), .I0(direction_N_4113), 
            .I1(encoder0_position[3]), .CO(n44113));
    SB_LUT4 position_2284_add_4_4_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[2]), .I3(n44111), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_4 (.CI(n44111), .I0(direction_N_4113), 
            .I1(encoder0_position[2]), .CO(n44112));
    SB_LUT4 position_2284_add_4_3_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder0_position[1]), .I3(n44110), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_3 (.CI(n44110), .I0(direction_N_4113), 
            .I1(encoder0_position[1]), .CO(n44111));
    SB_LUT4 position_2284_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2284_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2284_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n44110));
    SB_DFFE position_2284__i31 (.Q(encoder0_position[31]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i30 (.Q(encoder0_position[30]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i29 (.Q(encoder0_position[29]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i28 (.Q(encoder0_position[28]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i27 (.Q(encoder0_position[27]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i26 (.Q(encoder0_position[26]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i25 (.Q(encoder0_position[25]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i24 (.Q(encoder0_position[24]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i23 (.Q(encoder0_position[23]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i22 (.Q(encoder0_position[22]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i21 (.Q(encoder0_position[21]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i20 (.Q(encoder0_position[20]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i19 (.Q(encoder0_position[19]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i18 (.Q(encoder0_position[18]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i17 (.Q(encoder0_position[17]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i16 (.Q(encoder0_position[16]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i15 (.Q(encoder0_position[15]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i14 (.Q(encoder0_position[14]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i13 (.Q(encoder0_position[13]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i12 (.Q(encoder0_position[12]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i11 (.Q(encoder0_position[11]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i10 (.Q(encoder0_position[10]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i9 (.Q(encoder0_position[9]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i8 (.Q(encoder0_position[8]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i7 (.Q(encoder0_position[7]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i6 (.Q(encoder0_position[6]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i5 (.Q(encoder0_position[5]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i4 (.Q(encoder0_position[4]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i3 (.Q(encoder0_position[3]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i2 (.Q(encoder0_position[2]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2284__i1 (.Q(encoder0_position[1]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 i39793_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_4116));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i39793_4_lut.LUT_INIT = 16'h8421;
    SB_DFFE position_2284__i0 (.Q(encoder0_position[0]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n2269), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n2269), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i15351_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4116), .I2(b_new[1]), 
            .I3(b_prev), .O(n29427));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15351_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15336_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4116), .I2(a_new[1]), 
            .I3(a_prev), .O(n29412));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15336_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Kp[8] , \Ki[1] , \PID_CONTROLLER.integral_23__N_3996 , 
            \Ki[0] , \Ki[11] , \Ki[12] , \Ki[2] , \Ki[13] , \Ki[14] , 
            \Ki[3] , \Kp[9] , \Ki[15] , \Kp[10] , \Ki[4] , \Kp[11] , 
            \Ki[5] , IntegralLimit, \Ki[6] , \Ki[7] , \Kp[12] , \Kp[3] , 
            \Ki[9] , PWMLimit, \Kp[4] , \Kp[14] , \Kp[5] , \Kp[1] , 
            \Kp[2] , \Kp[0] , \Kp[13] , \Ki[8] , \Ki[10] , \Kp[15] , 
            \Kp[6] , \Kp[7] , duty, clk16MHz, control_update, deadband, 
            VCC_net, \PID_CONTROLLER.integral , n29289, setpoint, motor_state, 
            n29804, n29803, n29802, n29801, n29800, n29799, n29798, 
            n29797, n29796, n29795, n29794, n29793, n29792, n29791, 
            n29790, n29789, n29788, n29787, n29786, n29785, n29784, 
            n29783, n29782) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \Kp[8] ;
    input \Ki[1] ;
    output [23:0]\PID_CONTROLLER.integral_23__N_3996 ;
    input \Ki[0] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[2] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[3] ;
    input \Kp[9] ;
    input \Ki[15] ;
    input \Kp[10] ;
    input \Ki[4] ;
    input \Kp[11] ;
    input \Ki[5] ;
    input [23:0]IntegralLimit;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Kp[12] ;
    input \Kp[3] ;
    input \Ki[9] ;
    input [23:0]PWMLimit;
    input \Kp[4] ;
    input \Kp[14] ;
    input \Kp[5] ;
    input \Kp[1] ;
    input \Kp[2] ;
    input \Kp[0] ;
    input \Kp[13] ;
    input \Ki[8] ;
    input \Ki[10] ;
    input \Kp[15] ;
    input \Kp[6] ;
    input \Kp[7] ;
    output [23:0]duty;
    input clk16MHz;
    output control_update;
    input [23:0]deadband;
    input VCC_net;
    output [23:0]\PID_CONTROLLER.integral ;
    input n29289;
    input [23:0]setpoint;
    input [23:0]motor_state;
    input n29804;
    input n29803;
    input n29802;
    input n29801;
    input n29800;
    input n29799;
    input n29798;
    input n29797;
    input n29796;
    input n29795;
    input n29794;
    input n29793;
    input n29792;
    input n29791;
    input n29790;
    input n29789;
    input n29788;
    input n29787;
    input n29786;
    input n29785;
    input n29784;
    input n29783;
    input n29782;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [19:0]n13789;
    wire [18:0]n14588;
    
    wire n44656, n44449;
    wire [20:0]n12425;
    
    wire n296, n44450;
    wire [23:0]n1;
    
    wire n597;
    wire [47:0]n257;
    wire [21:0]n11938;
    
    wire n512, n44707, n44657, n1105, n44655;
    wire [7:0]n19029;
    wire [6:0]n19173;
    
    wire n484, n44580;
    wire [21:0]n11407;
    
    wire n223, n44448, n44581, n131, n62, n44708, n819, n892, 
        n195, n965, n204, n1038, n411, n44579, n268, n670, n150, 
        n44447, n661, n1111, n743, n734, n8, n77, n341, n807, 
        n414;
    wire [23:0]n130;
    wire [23:0]n182;
    
    wire n181;
    wire [23:0]n207;
    wire [19:0]n13349;
    
    wire n44446, n338, n44578, n44445, n155, n86;
    wire [1:0]n19493;
    
    wire n42826;
    wire [2:0]n19469;
    
    wire n1032, n44654, n44444, n17, n487, n159, n439, n44706, 
        n959, n44653, n816, n232, n560, n265, n44577, n44443, 
        n192, n44576, n44442, n889, n44441, n305, n271, n661_adj_4878, 
        n1102, n44440, n1029, n44439, n50, n119, n956, n44438, 
        n883, n44437;
    wire [15:0]n16533;
    wire [14:0]n17044;
    
    wire n44575, n1117, n44574, n810, n44436, n737, n44435, n1044, 
        n44573, n880, n664, n44434, n591, n44433, n518, n44432, 
        n886, n44652, n445, n44431, n971, n44572, n813, n44651;
    wire [23:0]n1_adj_5416;
    
    wire n344, n1023, n1041, n417, n490, n52010;
    wire [3:0]n19453;
    
    wire n6;
    wire [4:0]n19404;
    
    wire n52014, n378, n98, n1096, n52012, n204_adj_4880, n29, 
        n43024, n52020, n953, n4;
    wire [3:0]n19429;
    
    wire n6_adj_4882, n8_adj_4883, n451, n6_adj_4884, n51035, n524, 
        n962, n597_adj_4885, n171, n244, n670_adj_4886, n1035;
    wire [1:0]n19501;
    
    wire n743_adj_4887, n317, n816_adj_4888, n889_adj_4889, n131_adj_4890, 
        n62_adj_4891, n411_adj_4892, n551, n624, n697, n390, n1108, 
        n1026, n962_adj_4893, n1035_adj_4894, n1108_adj_4895, n463, 
        n536, n609, n1099, n682, n113_adj_4896, n44, n366, n44705, 
        n755, n186_adj_4897, n259, n734_adj_4898, n332, n828, n658, 
        n405, n478, n901, n83, n14, n551_adj_4899, n28939, n28830, 
        n29234, n624_adj_4900, n974, n898, n44571, n372, n44430, 
        n299_adj_4901, n44429, n28934, n28929, n28924, n28919, n28914, 
        n28909, n28904, n28899, n28894, n28889, n28884, n28879, 
        n28874, n28869, n697_adj_4902, n770, n28864, n28859, n28854, 
        n28849, n28844, n28839, n28834, n226_adj_4903, n44428, n740, 
        n44650, n490_adj_4904, n28829, n52050, n52052, n210_adj_4905, 
        n52056, n42851, n825, n44570, n52060, n8_adj_4906, n770_adj_4907, 
        n6_adj_4908, n4_adj_4909, n50780, n667, n44649, n293, n44704, 
        n220, n44703, n1114, n116, n47, n484_adj_4910, n107_adj_4911, 
        n38, n180, n253, n104, n35, n557, n630, n83_adj_4915, 
        n326, n14_adj_4917, n92, n95, n23, n26, n399, n1047, 
        n472, n147, n44702, n156, n594, n44648, n229, n5_adj_4918, 
        n74, n545, n445_adj_4919, n1120, n618, n877, n691, n89, 
        n20, n95_adj_4921, n518_adj_4922, n26_adj_4923, n156_adj_4924, 
        n229_adj_4925, n302_adj_4926, n807_adj_4927, n752, n44569, 
        n153, n44427, n764, n837, n910, n375, n168, n448, n521, 
        n302_adj_4930, n104_adj_4931, n35_adj_4932, n241, n594_adj_4933, 
        n177, n667_adj_4934, n314, n375_adj_4935, n740_adj_4936, n250, 
        n162, n323, n110_adj_4938, n41, n396, n469, n235, n183_adj_4939, 
        n950, n542, n615, n256, n688, n761, n880_adj_4940, n165, 
        n813_adj_4941, n953_adj_4942, n387, n886_adj_4943, n460, n959_adj_4944, 
        n238, n1032_adj_4945, n448_adj_4946, n1105_adj_4947, n533, 
        n834, n1026_adj_4948;
    wire [23:0]n356;
    wire [0:0]n11431;
    wire [0:0]n10900;
    
    wire n43317, n11_adj_4949, n80;
    wire [47:0]n306;
    
    wire n43316, n43315;
    wire [18:0]n14189;
    
    wire n44426, n679, n44568, n44425, n521_adj_4951, n44647, n44424, 
        n43314;
    wire [31:0]counter;   // verilog/motorControl.v(23[11:18])
    
    wire n18, n44423, n43313, n606, n44567, n12;
    wire [20:0]n12908;
    
    wire n44701, counter_31__N_3995, n50434, n30, n43312, n44422, 
        n44566, n44421, n44700, n44646, n43311, n44420, n43310, 
        n28, n29_adj_4953, n27, n10_adj_4954, n9_adj_4955, n50533, 
        n44419, n44565, n44418, n44564, n43309, n44417, n44699, 
        n1099_adj_4956, n329, n907, n43308, n43307, n43306, n44416, 
        n44645, n44563, n44415, n168_adj_4960, n44414, n44562, n311, 
        n43305, n44698, n44644, n44413, n44412, n44561, n43304, 
        n44411, n177_adj_4962, n43303, n44410, n44643, n44697, n44642;
    wire [13:0]n17493;
    
    wire n44560, n44409, n44408, n44559;
    wire [9:0]n18749;
    wire [8:0]n18948;
    
    wire n44407, n44406, n241_adj_4964;
    wire [23:0]n436;
    
    wire n10863, n28828, n28833, n980, n28838, n28843, n28848, 
        n28853, n28858, n28863, n4_adj_4966, n28868, n28873, n28878, 
        n44558, n44405, n43302, n44404, n28883, n44557, n44403, 
        n28888, n44696, n28893, n44402, n28898, n28903, n28908, 
        n44556, n44401, n28913, n44400, n43301, n28918, n28923;
    wire [23:0]n1_adj_5417;
    wire [17:0]n15309;
    
    wire n44641, n44640, n28928, n44399, n44555, n44695, n43300;
    wire [17:0]n14949;
    
    wire n44398, n28933, n44554, n39, n44397, n44694, n44396, 
        n44639, n44553, n44395, n41_adj_4974, n44638, n44552, n44551, 
        n44394, n45, n44393, n44392, n44693, n43, n44637, n44550, 
        n29_adj_4975, n31, n37, n23_adj_4976, n25_adj_4977, n35_adj_4978, 
        n44391, n44390, n44549, n44389, n44636, n44388, n44548, 
        n44547, n44387, n44635, n44386, n44385, n44692, n44384, 
        n44691, n44383, n44634, n28621;
    wire [5:0]n19285;
    
    wire n44546, n44382, n44633, n384, n44381, n44545, n11_adj_4980;
    wire [16:0]n15633;
    
    wire n44380, n13, n15, n44544, n44379, n122_adj_4981, n44378, 
        n53, n44690, n314_adj_4982, n27_adj_4983, n33, n9_adj_4984, 
        n17_adj_4985, n19, n21_adj_4986, n457_adj_4987, n54467, n54438, 
        n44543, n44689, n44632, n44377, n44688, n44631, n44542;
    wire [31:0]n34;
    
    wire n44109, n44108, n308, n387_adj_4992, n12_adj_4993, n10_adj_4994, 
        n30_adj_4995, n44376, n44107, n44375, n44541, n54484, n54881, 
        n44374, n54877, n55414, n44106, n44373, n44105, n44630, 
        n55151, n55480, n53_adj_5001, n122_adj_5002, n16_adj_5003, 
        n746, n44372, n44104, n44103, n6_adj_5006, n55286, n55287, 
        n8_adj_5007, n673, n44371, n24_adj_5008, n54405, n54400, 
        n55147, n54868, n74_adj_5009, n4_adj_5010, n5_adj_5011, n530, 
        n80_adj_5012, n44102, n55360, n11_adj_5014, n731, n55361, 
        n54428, n54426, n55500, n55277, n524_adj_5018, n44629, n55572, 
        n600, n44370;
    wire [12:0]n17884;
    
    wire n1050, n44540, n977, n44539, n55573, n55553, n54407, 
        n153_adj_5020, n55402, n40, n55404, n409, n147_adj_5024, 
        n527, n44369, n44101, n41_adj_5026, n39_adj_5028, n45_adj_5029, 
        n250_adj_5031, n460_adj_5033, n36533, n43_adj_5034, n37_adj_5035;
    wire [23:0]n1_adj_5418;
    
    wire n189, n262, n44100, n29_adj_5038, n454_adj_5039, n44368, 
        n220_adj_5040, n44099, n43299, n44098, n44097, n381, n44367, 
        n904, n44538, n44096, n293_adj_5044, n603, n31_adj_5045, 
        n308_adj_5046, n44366, n43298, n831, n44537, n235_adj_5047, 
        n44365, n23_adj_5048, n44095, n44094, n162_adj_5051, n44364, 
        n25_adj_5052, n44093, n366_adj_5054, n758, n44536, n20_adj_5055, 
        n89_adj_5056, n588, n44687, n44092, n676, n35_adj_5059, 
        n33_adj_5061, n11_adj_5062, n13_adj_5063, n15_adj_5064, n27_adj_5065, 
        n9_adj_5066, n17_adj_5067, n226_adj_5068, n19_adj_5069, n21_adj_5070, 
        n54380, n54371, n12_adj_5072, n10_adj_5078, n30_adj_5079, 
        n54398, n54781, n54774, n55380, n55119, n55476, n6_adj_5084, 
        n55370, n16_adj_5085, n44091, n451_adj_5086, n44628;
    wire [7:0]n19109;
    
    wire n700, n44363, n8_adj_5087, n515, n44686, n627, n44362, 
        n24_adj_5088, n55371, n54353, n685, n44535, n533_adj_5089, 
        n54351, n55149, n55281, n44090, n378_adj_5090, n44627, n4_adj_5091, 
        n554, n44361, n612, n44534, n481, n44360, n43297, n44089, 
        n55368, n44088, n55369, n44087, n54367, n323_adj_5093, n44086, 
        n408, n44359, n44085, n335_adj_5094, n44358, n305_adj_5095, 
        n44626, n539, n44533, n466, n44532, n54365, n55502, n262_adj_5096, 
        n44357, n55283, n189_adj_5097, n44356, n44084, n44083, n44082, 
        n43296, n393, n44531, n44081, n47_adj_5098, n116_adj_5099, 
        n43295;
    wire [15:0]n16245;
    
    wire n44355, n44354, n44080, n442_adj_5100, n44685, n232_adj_5101, 
        n44625, n44079, n320, n44530, n1114_adj_5103, n44353, n1041_adj_5105, 
        n44352, n159_adj_5106, n44624, n968, n44351, n55574, n55575, 
        n55551, n54355, n43294, n43293, n247, n44529, n55408, 
        n895, n44350, n40_adj_5110, n55410, n439_adj_5111, n55411, 
        n822, n44349, n512_adj_5112, n369_adj_5113, n44684, n17_adj_5114, 
        n86_adj_5115, n749, n44348, n174, n44528;
    wire [8:0]n18849;
    
    wire n700_adj_5116, n44623, n32, n101, n676_adj_5117, n44347, 
        n603_adj_5118, n44346, n43292, n627_adj_5119, n44622, n530_adj_5120, 
        n44345;
    wire [11:0]n18221;
    
    wire n980_adj_5121, n44527, n907_adj_5122, n44526, n457_adj_5123, 
        n44344, n43291, n43290, n749_adj_5124, n41_adj_5125, n384_adj_5126, 
        n44343, n39_adj_5127, n33_adj_5128, n35_adj_5129, n37_adj_5130, 
        n29_adj_5131, n43289, n43288, n43287, n31_adj_5134, n23_adj_5135, 
        n43286, n43285, n43284, n804, n585, n43283, n25_adj_5141, 
        n45_adj_5142, n299_adj_5143, n43_adj_5144, n311_adj_5145, n44342, 
        n296_adj_5146, n44683, n554_adj_5147, n44621, n238_adj_5148, 
        n44341, n834_adj_5150, n44525, n165_adj_5151, n44340, n43282, 
        n110_adj_5153, n43281, n9_adj_5155, n41_adj_5156, n17_adj_5157, 
        n223_adj_5158, n44682, n19_adj_5160, n23_adj_5161, n92_adj_5162, 
        n183_adj_5163, n21_adj_5164, n43280, n761_adj_5166, n44524, 
        n481_adj_5167, n44620, n43279;
    wire [14:0]n16789;
    
    wire n44339, n11_adj_5168, n13_adj_5169, n15_adj_5170, n27_adj_5171;
    wire [23:0]n382;
    
    wire n54521, n54907, n56813, n54905, n56808, n1117_adj_5174, 
        n44338, n43278, n150_adj_5176, n44681, n688_adj_5177, n44523, 
        n1044_adj_5178, n44337, n615_adj_5179, n44522, n971_adj_5180, 
        n44336, n43277, n898_adj_5182, n44335, n408_adj_5183, n44619, 
        n825_adj_5184, n44334, n542_adj_5185, n44521, n42958;
    wire [2:0]n19484;
    
    wire n658_adj_5186, n54553, n54560, n16_adj_5187, n256_adj_5188, 
        n822_adj_5189, n8_adj_5191, n24_adj_5192, n54571, n54947, 
        n329_adj_5194, n402_adj_5195, n335_adj_5196, n54943, n43276, 
        n55434, n55183, n55492, n195_adj_5198, n752_adj_5199, n44333, 
        n402_adj_5200, n43275, n469_adj_5201, n44520, n731_adj_5202, 
        n54525, n54911, n396_adj_5204, n606_adj_5205, n56801, n54899, 
        n56795, n12_adj_5208, n54501, n56819, n10_adj_5210, n30_adj_5211, 
        n895_adj_5212, n54529, n56839, n77_adj_5213, n8_adj_5214, 
        n54527, n679_adj_5216, n44332, n56832, n804_adj_5218, n55173, 
        n56835, n43274, n475, n548, n54909, n55318, n44331, n591_adj_5222, 
        n621, n268_adj_5223, n44519, n54513, n56799, n694, n55167, 
        n43273, n56824, n55422, n475_adj_5227, n44618, n56790, n55524, 
        n56787, n6_adj_5229, n55294, n44518, n44330, n16_adj_5231, 
        n877_adj_5232, n381_adj_5233, n968_adj_5234, n54487, n43272, 
        n44680, n44617, n44616, n8_adj_5238, n372_adj_5239, n44329, 
        n44517, n44328, n24_adj_5241, n44327, n767, n44679, n341_adj_5242, 
        n414_adj_5243, n44678, n28622, n55295, n548_adj_5244, n487_adj_5245, 
        n54490, n840, n560_adj_5246, n56785, n55145, n44723, n101_adj_5247, 
        n44722, n950_adj_5248, n54858, n12_adj_5249, n4_adj_5250, 
        n55298, n55299, n44326, n44516, n44325, n10_adj_5251, n32_adj_5252, 
        n30_adj_5253, n54549, n54547, n55462, n54850, n621_adj_5255, 
        n55546, n174_adj_5256, n55547, n125_adj_5257, n56, n6_adj_5258, 
        n55300, n55301, n54533, n247_adj_5259, n198_adj_5261, n454_adj_5264, 
        n54531, n55143, n320_adj_5265, n54848, n55521, n54535, n694_adj_5266, 
        n55396, n54856, n54263, n4_adj_5268, n55292, n55293, n54503, 
        n55464, n54860, n55548, n55549, n55519, n54492, n44677;
    wire [6:0]n19236;
    
    wire n44324, n44323, n44676, n55398, n54866, n44322, n55488, 
        n55486, n47_adj_5269, n52036, n44721;
    wire [9:0]n18629;
    
    wire n43477, n43476, n43475, n44720, n43474;
    wire [16:0]n15956;
    
    wire n44615, n44321, n44515, n44614;
    wire [4:0]n19369;
    
    wire n417_adj_5270, n44514, n338_adj_5271, n44320, n265_adj_5272, 
        n44319, n478_adj_5273, n43473, n44675, n405_adj_5274, n43472, 
        n332_adj_5275, n43471, n192_adj_5276, n44318, n344_adj_5277, 
        n44513, n259_adj_5278, n43470, n186_adj_5279, n43469, n44_adj_5280, 
        n113_adj_5281, n50_adj_5282, n119_adj_5283, n271_adj_5285, n44512;
    wire [13:0]n17269;
    
    wire n1120_adj_5286, n44317, n1047_adj_5287, n44316, n44719, n44613, 
        n198_adj_5288, n44511, n974_adj_5289, n44315, n56_adj_5290, 
        n125_adj_5291, n1111_adj_5292, n44612, n1102_adj_5293, n44674, 
        n44718;
    wire [10:0]n18508;
    
    wire n910_adj_5294, n44510, n44717, n1038_adj_5295, n44611, n837_adj_5296, 
        n44509, n901_adj_5297, n44314, n965_adj_5298, n44610, n1029_adj_5299, 
        n44673, n764_adj_5300, n44508, n828_adj_5301, n44313, n956_adj_5302, 
        n44672, n755_adj_5303, n44312, n682_adj_5304, n44311, n28938, 
        n44716, n691_adj_5305, n44507, n1096_adj_5306, n44715, n883_adj_5307, 
        n44671, n892_adj_5308, n44609, n609_adj_5309, n44310, n618_adj_5310, 
        n44506, n536_adj_5311, n44309, n819_adj_5312, n44608, n463_adj_5313, 
        n44308, n545_adj_5314, n44505, n390_adj_5315, n44307, n317_adj_5316, 
        n44306, n472_adj_5317, n44504, n244_adj_5318, n44305, n171_adj_5319, 
        n44304, n746_adj_5320, n44607, n810_adj_5321, n44670, n399_adj_5322, 
        n44503, n29_adj_5323, n98_adj_5324;
    wire [12:0]n17689;
    
    wire n1050_adj_5325, n44303, n326_adj_5326, n44502, n977_adj_5327, 
        n44302, n737_adj_5328, n44669, n673_adj_5329, n44606, n904_adj_5330, 
        n44301, n831_adj_5331, n44300, n253_adj_5332, n44501, n180_adj_5333, 
        n44500, n758_adj_5334, n44299, n685_adj_5335, n44298, n1023_adj_5336, 
        n44714, n600_adj_5337, n44605, n38_adj_5338, n107_adj_5339, 
        n612_adj_5340, n44297, n539_adj_5341, n44296, n664_adj_5342, 
        n44668, n840_adj_5343, n44499, n466_adj_5344, n44295, n767_adj_5345, 
        n44498, n393_adj_5346, n44294, n527_adj_5347, n44604, n44497, 
        n44293, n44603, n44292, n44291, n44496;
    wire [5:0]n19333;
    
    wire n44290, n44289, n44495, n44288, n44287, n44602, n44494, 
        n44286, n44667, n44493, n44285, n44601;
    wire [11:0]n18053;
    
    wire n44284, n44283, n44492, n44282, n44281, n44280, n42908, 
        n44491, n44279, n44278, n44713, n44490, n44600, n44277, 
        n44276, n44489, n44275, n44599, n44274, n44488, n44273, 
        n44487;
    wire [10:0]n18365;
    
    wire n44272, n44271, n44270, n44666, n44269, n44712, n44486, 
        n44268, n43424, n43423, n43422, n44665, n44267, n43421, 
        n4_adj_5348, n44598, n44485, n44266, n44484, n44265, n44264, 
        n44597, n43420, n43419, n44263, n44483, n43418, n44262, 
        n43417, n44482, n44596, n44261, n44481, n44260, n44595, 
        n43416, n44480, n44259, n43415, n44258, n43233, n43232, 
        n43231, n43414, n43413, n44257, n43412, n43230, n43411, 
        n43229, n43228, n44479, n43227, n44256, n44255, n44664, 
        n43410, n44594, n44478, n43409, n43226, n43225, n43408, 
        n43224, n44254, n43407, n44253, n44252, n43406, n44251, 
        n43405, n43404, n43223, n44477, n43403, n43402, n44593, 
        n43222, n43221, n44476, n43220, n43401, n43219, n44250, 
        n44249, n43400, n43399, n44592, n44248, n43218, n44475, 
        n43217, n43398, n43216, n44247, n43397, n43396, n43215, 
        n43395, n44663, n43214, n43394, n44474, n43393, n44711, 
        n43213, n43392, n44591, n44473, n44472, n43391, n43212, 
        n43390, n43389, n43211, n43388, n43387, n43386, n43385, 
        n43384, n43383, n44662, n43382, n44590, n43381, n44471, 
        n43380, n44589, n44470, n43379, n44469, n54573, n54583, 
        n43378, n43377, n43376, n44468, n43375, n43374, n43373, 
        n44661, n43372, n43371, n43370, n43369, n44710, n44588, 
        n44467, n43368, n43367, n43366, n43365, n43364, n43363, 
        n44466, n43362, n44465, n43361, n43360, n44660, n44587, 
        n44464, n54607, n44586, n44463, n43359, n43358, n43357, 
        n43356, n54617, n44462, n44461, n44659, n44585, n44460, 
        n44459, n44584, n44458, n44583, n44457, n44658, n54605, 
        n44456, n6_adj_5351, n44709, n44455, n44454, n54640, n630_adj_5352, 
        n44582, n588_adj_5353, n44453, n6_adj_5354, n515_adj_5355, 
        n44452, n557_adj_5356, n442_adj_5357, n44451, n585_adj_5358, 
        n369_adj_5359, n4_adj_5360, n43040, n201_adj_5362, n9_adj_5363, 
        n11_adj_5364, n13_adj_5365, n4_adj_5366, n15_adj_5367, n21_adj_5368, 
        n9_adj_5369, n11_adj_5370, n13_adj_5371, n15_adj_5372, n21_adj_5373, 
        n39_adj_5374, n41_adj_5375, n37_adj_5376, n35_adj_5377, n31_adj_5378, 
        n33_adj_5379, n27_adj_5380, n29_adj_5381, n45_adj_5382, n25_adj_5383, 
        n23_adj_5384, n17_adj_5385, n19_adj_5386, n43_adj_5387, n54630, 
        n54623, n12_adj_5388, n10_adj_5389, n30_adj_5390, n55027, 
        n55023, n55446, n55217, n55496, n16_adj_5391, n55316, n55317, 
        n8_adj_5392, n24_adj_5393, n54609, n55139, n54828, n4_adj_5394, 
        n55314, n55315, n54619, n55458, n54830, n55542, n55543, 
        n55527, n54611, n55392, n54836, n55482, n41_adj_5395, n37_adj_5396, 
        n39_adj_5397, n35_adj_5398, n19_adj_5399, n31_adj_5400, n33_adj_5401, 
        n29_adj_5402, n27_adj_5403, n23_adj_5404, n25_adj_5405, n43_adj_5406, 
        n45_adj_5407, n17_adj_5408, n54595, n54589, n12_adj_5409, 
        n10_adj_5410, n30_adj_5411, n54991, n54987, n55440, n55201, 
        n55494, n16_adj_5412, n55308, n55309, n8_adj_5413, n24_adj_5414, 
        n54575, n55141, n54838, n4_adj_5415, n55306, n55307, n54585, 
        n55460, n54840, n55544, n55545, n55523, n54577, n55394, 
        n54846, n55484;
    
    SB_LUT4 add_5179_17_lut (.I0(GND_net), .I1(n14588[14]), .I2(GND_net), 
            .I3(n44656), .O(n13789[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_5 (.CI(n44449), .I0(n12425[2]), .I1(n296), .CO(n44450));
    SB_LUT4 mult_16_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_8_lut (.I0(GND_net), .I1(n11938[5]), .I2(n512), 
            .I3(n44707), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_17 (.CI(n44656), .I0(n14588[14]), .I1(GND_net), 
            .CO(n44657));
    SB_LUT4 add_5179_16_lut (.I0(GND_net), .I1(n14588[13]), .I2(n1105), 
            .I3(n44655), .O(n13789[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5495_7_lut (.I0(GND_net), .I1(n19173[4]), .I2(n484), .I3(n44580), 
            .O(n19029[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5073_4_lut (.I0(GND_net), .I1(n12425[1]), .I2(n223), .I3(n44448), 
            .O(n11407[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5495_7 (.CI(n44580), .I0(n19173[4]), .I1(n484), .CO(n44581));
    SB_LUT4 mult_17_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i89_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5073_4 (.CI(n44448), .I0(n12425[1]), .I1(n223), .CO(n44449));
    SB_LUT4 mult_17_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i42_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_8 (.CI(n44707), .I0(n11938[5]), .I1(n512), 
            .CO(n44708));
    SB_LUT4 mult_17_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i600_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5179_16 (.CI(n44655), .I0(n14588[13]), .I1(n1105), .CO(n44656));
    SB_LUT4 mult_17_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5495_6_lut (.I0(GND_net), .I1(n19173[3]), .I2(n411), .I3(n44579), 
            .O(n19029[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5073_3_lut (.I0(GND_net), .I1(n12425[0]), .I2(n150), .I3(n44447), 
            .O(n11407[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i445_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5495_6 (.CI(n44579), .I0(n19173[3]), .I1(n411), .CO(n44580));
    SB_CARRY add_5073_3 (.CI(n44447), .I0(n12425[0]), .I1(n150), .CO(n44448));
    SB_LUT4 mult_17_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5073_2_lut (.I0(GND_net), .I1(n8), .I2(n77), .I3(GND_net), 
            .O(n11407[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i230_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5073_2 (.CI(GND_net), .I0(n8), .I1(n77), .CO(n44447));
    SB_LUT4 mult_16_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i6_3_lut (.I0(n130[5]), .I1(n182[5]), .I2(n181), .I3(GND_net), 
            .O(n207[5]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5118_22_lut (.I0(GND_net), .I1(n13349[19]), .I2(GND_net), 
            .I3(n44446), .O(n12425[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5495_5_lut (.I0(GND_net), .I1(n19173[2]), .I2(n338), .I3(n44578), 
            .O(n19029[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_21_lut (.I0(GND_net), .I1(n13349[18]), .I2(GND_net), 
            .I3(n44445), .O(n12425[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i6_3_lut (.I0(n207[5]), .I1(IntegralLimit[5]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [5]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i59_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5118_21 (.CI(n44445), .I0(n13349[18]), .I1(GND_net), 
            .CO(n44446));
    SB_LUT4 i1_4_lut (.I0(n19493[0]), .I1(n42826), .I2(\Ki[2] ), .I3(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .O(n19469[1]));   // verilog/motorControl.v(52[27:38])
    defparam i1_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 add_5179_15_lut (.I0(GND_net), .I1(n14588[12]), .I2(n1032), 
            .I3(n44654), .O(n13789[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_20_lut (.I0(GND_net), .I1(n13349[17]), .I2(GND_net), 
            .I3(n44444), .O(n12425[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_7_lut (.I0(GND_net), .I1(n11938[4]), .I2(n439), 
            .I3(n44706), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_15 (.CI(n44654), .I0(n14588[12]), .I1(n1032), .CO(n44655));
    SB_CARRY add_5118_20 (.CI(n44444), .I0(n13349[17]), .I1(GND_net), 
            .CO(n44445));
    SB_LUT4 add_5179_14_lut (.I0(GND_net), .I1(n14588[11]), .I2(n959), 
            .I3(n44653), .O(n13789[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i549_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5495_5 (.CI(n44578), .I0(n19173[2]), .I1(n338), .CO(n44579));
    SB_LUT4 mult_17_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i21_3_lut (.I0(n130[20]), .I1(n182[20]), .I2(n181), 
            .I3(GND_net), .O(n207[20]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i21_3_lut (.I0(n207[20]), .I1(IntegralLimit[20]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [20]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5495_4_lut (.I0(GND_net), .I1(n19173[1]), .I2(n265), .I3(n44577), 
            .O(n19029[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5495_4 (.CI(n44577), .I0(n19173[1]), .I1(n265), .CO(n44578));
    SB_LUT4 add_5118_19_lut (.I0(GND_net), .I1(n13349[16]), .I2(GND_net), 
            .I3(n44443), .O(n12425[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5495_3_lut (.I0(GND_net), .I1(n19173[0]), .I2(n192), .I3(n44576), 
            .O(n19029[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_19 (.CI(n44443), .I0(n13349[16]), .I1(GND_net), 
            .CO(n44444));
    SB_LUT4 add_5118_18_lut (.I0(GND_net), .I1(n13349[15]), .I2(GND_net), 
            .I3(n44442), .O(n12425[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i598_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5118_18 (.CI(n44442), .I0(n13349[15]), .I1(GND_net), 
            .CO(n44443));
    SB_LUT4 add_5118_17_lut (.I0(GND_net), .I1(n13349[14]), .I2(GND_net), 
            .I3(n44441), .O(n12425[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_17 (.CI(n44441), .I0(n13349[14]), .I1(GND_net), 
            .CO(n44442));
    SB_LUT4 mult_17_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4878));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i22_3_lut (.I0(n130[21]), .I1(n182[21]), .I2(n181), 
            .I3(GND_net), .O(n207[21]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5118_16_lut (.I0(GND_net), .I1(n13349[13]), .I2(n1102), 
            .I3(n44440), .O(n12425[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_16 (.CI(n44440), .I0(n13349[13]), .I1(n1102), .CO(n44441));
    SB_CARRY add_5495_3 (.CI(n44576), .I0(n19173[0]), .I1(n192), .CO(n44577));
    SB_LUT4 add_5118_15_lut (.I0(GND_net), .I1(n13349[12]), .I2(n1029), 
            .I3(n44439), .O(n12425[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5495_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n19029[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_15 (.CI(n44439), .I0(n13349[12]), .I1(n1029), .CO(n44440));
    SB_CARRY add_5179_14 (.CI(n44653), .I0(n14588[11]), .I1(n959), .CO(n44654));
    SB_CARRY add_5495_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n44576));
    SB_LUT4 add_5118_14_lut (.I0(GND_net), .I1(n13349[11]), .I2(n956), 
            .I3(n44438), .O(n12425[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_14 (.CI(n44438), .I0(n13349[11]), .I1(n956), .CO(n44439));
    SB_LUT4 add_5118_13_lut (.I0(GND_net), .I1(n13349[10]), .I2(n883), 
            .I3(n44437), .O(n12425[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5319_17_lut (.I0(GND_net), .I1(n17044[14]), .I2(GND_net), 
            .I3(n44575), .O(n16533[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_13 (.CI(n44437), .I0(n13349[10]), .I1(n883), .CO(n44438));
    SB_LUT4 add_5319_16_lut (.I0(GND_net), .I1(n17044[13]), .I2(n1117), 
            .I3(n44574), .O(n16533[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_16 (.CI(n44574), .I0(n17044[13]), .I1(n1117), .CO(n44575));
    SB_LUT4 add_5118_12_lut (.I0(GND_net), .I1(n13349[9]), .I2(n810), 
            .I3(n44436), .O(n12425[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_12 (.CI(n44436), .I0(n13349[9]), .I1(n810), .CO(n44437));
    SB_LUT4 add_5118_11_lut (.I0(GND_net), .I1(n13349[8]), .I2(n737), 
            .I3(n44435), .O(n12425[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5319_15_lut (.I0(GND_net), .I1(n17044[12]), .I2(n1044), 
            .I3(n44573), .O(n16533[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_15 (.CI(n44573), .I0(n17044[12]), .I1(n1044), .CO(n44574));
    SB_CARRY add_5118_11 (.CI(n44435), .I0(n13349[8]), .I1(n737), .CO(n44436));
    SB_LUT4 mux_15_i22_3_lut (.I0(n207[21]), .I1(IntegralLimit[21]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [21]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5118_10_lut (.I0(GND_net), .I1(n13349[7]), .I2(n664), 
            .I3(n44434), .O(n12425[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_10 (.CI(n44434), .I0(n13349[7]), .I1(n664), .CO(n44435));
    SB_LUT4 add_5118_9_lut (.I0(GND_net), .I1(n13349[6]), .I2(n591), .I3(n44433), 
            .O(n12425[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_9 (.CI(n44433), .I0(n13349[6]), .I1(n591), .CO(n44434));
    SB_LUT4 add_5118_8_lut (.I0(GND_net), .I1(n13349[5]), .I2(n518), .I3(n44432), 
            .O(n12425[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_8 (.CI(n44432), .I0(n13349[5]), .I1(n518), .CO(n44433));
    SB_LUT4 add_5179_13_lut (.I0(GND_net), .I1(n14588[10]), .I2(n886), 
            .I3(n44652), .O(n13789[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_7_lut (.I0(GND_net), .I1(n13349[4]), .I2(n445), .I3(n44431), 
            .O(n12425[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_7 (.CI(n44706), .I0(n11938[4]), .I1(n439), 
            .CO(n44707));
    SB_CARRY add_5179_13 (.CI(n44652), .I0(n14588[10]), .I1(n886), .CO(n44653));
    SB_LUT4 add_5319_14_lut (.I0(GND_net), .I1(n17044[11]), .I2(n971), 
            .I3(n44572), .O(n16533[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_14 (.CI(n44572), .I0(n17044[11]), .I1(n971), .CO(n44573));
    SB_CARRY add_5118_7 (.CI(n44431), .I0(n13349[4]), .I1(n445), .CO(n44432));
    SB_LUT4 add_5179_12_lut (.I0(GND_net), .I1(n14588[9]), .I2(n813), 
            .I3(n44651), .O(n13789[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[14]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i20_3_lut (.I0(n130[19]), .I1(n182[19]), .I2(n181), 
            .I3(GND_net), .O(n207[19]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i20_3_lut (.I0(n207[19]), .I1(IntegralLimit[19]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [19]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i19_3_lut (.I0(n130[18]), .I1(n182[18]), .I2(n181), 
            .I3(GND_net), .O(n207[18]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i19_3_lut (.I0(n207[18]), .I1(IntegralLimit[18]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [18]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i24_3_lut (.I0(n130[23]), .I1(n182[23]), .I2(n181), 
            .I3(GND_net), .O(n207[23]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i24_3_lut (.I0(n207[23]), .I1(IntegralLimit[23]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [23]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_26_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[15]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i23_3_lut (.I0(n130[22]), .I1(n182[22]), .I2(n181), 
            .I3(GND_net), .O(n207[22]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i23_3_lut (.I0(n207[22]), .I1(IntegralLimit[22]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [22]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(\PID_CONTROLLER.integral_23__N_3996 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [23]), .O(n52010));   // verilog/motorControl.v(52[27:38])
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'h93a0;
    SB_LUT4 i1_4_lut_adj_1701 (.I0(n19453[2]), .I1(n6), .I2(\Kp[4] ), 
            .I3(n1[18]), .O(n19404[3]));   // verilog/motorControl.v(52[18:24])
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'h9666;
    SB_LUT4 i1_4_lut_adj_1702 (.I0(\Ki[5] ), .I1(\Ki[4] ), .I2(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [19]), .O(n52014));   // verilog/motorControl.v(52[27:38])
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_17_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [21]), .O(n52012));   // verilog/motorControl.v(52[27:38])
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_16_i138_2_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204_adj_4880));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n52012), .I1(n43024), .I2(n52014), 
            .I3(n52010), .O(n52020));   // verilog/motorControl.v(52[27:38])
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'h6996;
    SB_LUT4 mult_16_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28775_4_lut (.I0(n19493[0]), .I1(\Ki[2] ), .I2(n42826), .I3(\PID_CONTROLLER.integral_23__N_3996 [20]), 
            .O(n4));   // verilog/motorControl.v(52[27:38])
    defparam i28775_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i28867_4_lut (.I0(n19429[2]), .I1(\Ki[4] ), .I2(n6_adj_4882), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [18]), .O(n8_adj_4883));   // verilog/motorControl.v(52[27:38])
    defparam i28867_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_17_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n6_adj_4884), .I1(n8_adj_4883), .I2(n4), 
            .I3(n52020), .O(n51035));   // verilog/motorControl.v(52[27:38])
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4885));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4886));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28785_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n19501[0]));   // verilog/motorControl.v(52[18:24])
    defparam i28785_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_17_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4887));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4888));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4889));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i89_2_lut (.I0(\Kp[1] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131_adj_4890));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i42_2_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_4891));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4892));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4893));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4894));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4895));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4896));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_6_lut (.I0(GND_net), .I1(n11938[3]), .I2(n366), 
            .I3(n44705), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4897));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4898));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4899));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i371_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR result__i1 (.Q(duty[1]), .C(clk16MHz), .E(n28830), .D(n28939), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 mult_16_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4900));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5319_13_lut (.I0(GND_net), .I1(n17044[10]), .I2(n898), 
            .I3(n44571), .O(n16533[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_6_lut (.I0(GND_net), .I1(n13349[3]), .I2(n372), .I3(n44430), 
            .O(n12425[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_6 (.CI(n44430), .I0(n13349[3]), .I1(n372), .CO(n44431));
    SB_CARRY add_5319_13 (.CI(n44571), .I0(n17044[10]), .I1(n898), .CO(n44572));
    SB_LUT4 add_5118_5_lut (.I0(GND_net), .I1(n13349[2]), .I2(n299_adj_4901), 
            .I3(n44429), .O(n12425[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR result__i2 (.Q(duty[2]), .C(clk16MHz), .E(n28830), .D(n28934), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i3 (.Q(duty[3]), .C(clk16MHz), .E(n28830), .D(n28929), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i4 (.Q(duty[4]), .C(clk16MHz), .E(n28830), .D(n28924), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i5 (.Q(duty[5]), .C(clk16MHz), .E(n28830), .D(n28919), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i6 (.Q(duty[6]), .C(clk16MHz), .E(n28830), .D(n28914), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i7 (.Q(duty[7]), .C(clk16MHz), .E(n28830), .D(n28909), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i8 (.Q(duty[8]), .C(clk16MHz), .E(n28830), .D(n28904), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i9 (.Q(duty[9]), .C(clk16MHz), .E(n28830), .D(n28899), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i10 (.Q(duty[10]), .C(clk16MHz), .E(n28830), .D(n28894), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i11 (.Q(duty[11]), .C(clk16MHz), .E(n28830), .D(n28889), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i12 (.Q(duty[12]), .C(clk16MHz), .E(n28830), .D(n28884), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i13 (.Q(duty[13]), .C(clk16MHz), .E(n28830), .D(n28879), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i14 (.Q(duty[14]), .C(clk16MHz), .E(n28830), .D(n28874), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i15 (.Q(duty[15]), .C(clk16MHz), .E(n28830), .D(n28869), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 mult_16_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4902));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i518_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR result__i16 (.Q(duty[16]), .C(clk16MHz), .E(n28830), .D(n28864), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i17 (.Q(duty[17]), .C(clk16MHz), .E(n28830), .D(n28859), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i18 (.Q(duty[18]), .C(clk16MHz), .E(n28830), .D(n28854), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i19 (.Q(duty[19]), .C(clk16MHz), .E(n28830), .D(n28849), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i20 (.Q(duty[20]), .C(clk16MHz), .E(n28830), .D(n28844), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i21 (.Q(duty[21]), .C(clk16MHz), .E(n28830), .D(n28839), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFFESR result__i22 (.Q(duty[22]), .C(clk16MHz), .E(n28830), .D(n28834), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_CARRY mult_16_add_1225_6 (.CI(n44705), .I0(n11938[3]), .I1(n366), 
            .CO(n44706));
    SB_CARRY add_5179_12 (.CI(n44651), .I0(n14588[9]), .I1(n813), .CO(n44652));
    SB_CARRY add_5118_5 (.CI(n44429), .I0(n13349[2]), .I1(n299_adj_4901), 
            .CO(n44430));
    SB_LUT4 add_5118_4_lut (.I0(GND_net), .I1(n13349[1]), .I2(n226_adj_4903), 
            .I3(n44428), .O(n12425[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5179_11_lut (.I0(GND_net), .I1(n14588[8]), .I2(n740), 
            .I3(n44650), .O(n13789[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4904));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i330_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR result__i23 (.Q(duty[23]), .C(clk16MHz), .E(n28830), .D(n28829), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 i1_4_lut_adj_1706 (.I0(\Kp[4] ), .I1(\Kp[5] ), .I2(n1[19]), 
            .I3(n1[18]), .O(n52050));   // verilog/motorControl.v(52[18:24])
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_3_lut (.I0(\Kp[3] ), .I1(n52050), .I2(n1[20]), .I3(GND_net), 
            .O(n52052));   // verilog/motorControl.v(52[18:24])
    defparam i1_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_16_i142_2_lut (.I0(\Kp[2] ), .I1(n1[21]), .I2(GND_net), 
            .I3(GND_net), .O(n210_adj_4905));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1707 (.I0(\Kp[1] ), .I1(n210_adj_4905), .I2(n1[22]), 
            .I3(n52052), .O(n52056));   // verilog/motorControl.v(52[18:24])
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'h936c;
    SB_LUT4 i28787_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n42851));   // verilog/motorControl.v(52[18:24])
    defparam i28787_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_5319_12_lut (.I0(GND_net), .I1(n17044[9]), .I2(n825), 
            .I3(n44570), .O(n16533[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1708 (.I0(n42851), .I1(\Kp[0] ), .I2(n52056), 
            .I3(n1[23]), .O(n52060));   // verilog/motorControl.v(52[18:24])
    defparam i1_4_lut_adj_1708.LUT_INIT = 16'h695a;
    SB_LUT4 mux_14_i14_3_lut (.I0(n130[13]), .I1(n182[13]), .I2(n181), 
            .I3(GND_net), .O(n207[13]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i14_3_lut (.I0(n207[13]), .I1(IntegralLimit[13]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [13]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28989_4_lut (.I0(n19453[2]), .I1(\Kp[4] ), .I2(n6), .I3(n1[18]), 
            .O(n8_adj_4906));   // verilog/motorControl.v(52[18:24])
    defparam i28989_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_17_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4907));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n6_adj_4908), .I1(n8_adj_4906), .I2(n4_adj_4909), 
            .I3(n52060), .O(n50780));   // verilog/motorControl.v(52[18:24])
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'h6996;
    SB_CARRY add_5179_11 (.CI(n44650), .I0(n14588[8]), .I1(n740), .CO(n44651));
    SB_LUT4 add_5179_10_lut (.I0(GND_net), .I1(n14588[7]), .I2(n667), 
            .I3(n44649), .O(n13789[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_5_lut (.I0(GND_net), .I1(n11938[2]), .I2(n293), 
            .I3(n44704), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_5 (.CI(n44704), .I0(n11938[2]), .I1(n293), 
            .CO(n44705));
    SB_CARRY add_5179_10 (.CI(n44649), .I0(n14588[7]), .I1(n667), .CO(n44650));
    SB_LUT4 mult_16_add_1225_4_lut (.I0(GND_net), .I1(n11938[1]), .I2(n220), 
            .I3(n44703), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4910));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[16]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i13_3_lut (.I0(n130[12]), .I1(n182[12]), .I2(n181), 
            .I3(GND_net), .O(n207[12]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i13_3_lut (.I0(n207[12]), .I1(IntegralLimit[12]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [12]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4911));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[17]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[18]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[19]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i5_3_lut (.I0(n130[4]), .I1(n182[4]), .I2(n181), .I3(GND_net), 
            .O(n207[4]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i5_3_lut (.I0(n207[4]), .I1(IntegralLimit[4]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [4]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4915));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i9_3_lut (.I0(n130[8]), .I1(n182[8]), .I2(n181), .I3(GND_net), 
            .O(n207[8]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4917));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i9_3_lut (.I0(n207[8]), .I1(IntegralLimit[8]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [8]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i318_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5319_12 (.CI(n44570), .I0(n17044[9]), .I1(n825), .CO(n44571));
    SB_CARRY mult_16_add_1225_4 (.CI(n44703), .I0(n11938[1]), .I1(n220), 
            .CO(n44704));
    SB_LUT4 mult_16_add_1225_3_lut (.I0(GND_net), .I1(n11938[0]), .I2(n147), 
            .I3(n44702), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5179_9_lut (.I0(GND_net), .I1(n14588[6]), .I2(n594), .I3(n44648), 
            .O(n13789[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_3 (.CI(n44702), .I0(n11938[0]), .I1(n147), 
            .CO(n44703));
    SB_LUT4 mult_17_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[20]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4918), .I2(n74), 
            .I3(GND_net), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4919));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[21]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[22]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[23]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4921));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4922));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4923));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4924));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4925));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4926));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4927));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i543_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5118_4 (.CI(n44428), .I0(n13349[1]), .I1(n226_adj_4903), 
            .CO(n44429));
    SB_LUT4 add_5319_11_lut (.I0(GND_net), .I1(n17044[8]), .I2(n752), 
            .I3(n44569), .O(n16533[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_9 (.CI(n44648), .I0(n14588[6]), .I1(n594), .CO(n44649));
    SB_LUT4 add_5118_3_lut (.I0(GND_net), .I1(n13349[0]), .I2(n153), .I3(n44427), 
            .O(n12425[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i12_3_lut (.I0(n130[11]), .I1(n182[11]), .I2(n181), 
            .I3(GND_net), .O(n207[11]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i12_3_lut (.I0(n207[11]), .I1(IntegralLimit[11]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [11]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4930));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4931));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4932));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4933));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4934));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4935));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4936));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4938));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4939));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4940));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4941));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4942));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4943));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4944));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4945));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4946));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4947));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4948));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i690_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5319_11 (.CI(n44569), .I0(n17044[8]), .I1(n752), .CO(n44570));
    SB_LUT4 add_18_25_lut (.I0(GND_net), .I1(n11431[0]), .I2(n10900[0]), 
            .I3(n43317), .O(n356[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_3 (.CI(n44427), .I0(n13349[0]), .I1(n153), .CO(n44428));
    SB_LUT4 add_5118_2_lut (.I0(GND_net), .I1(n11_adj_4949), .I2(n80), 
            .I3(GND_net), .O(n12425[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_2 (.CI(GND_net), .I0(n11_adj_4949), .I1(n80), .CO(n44427));
    SB_LUT4 add_18_24_lut (.I0(GND_net), .I1(n257[22]), .I2(n306[22]), 
            .I3(n43316), .O(n356[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_24 (.CI(n43316), .I0(n257[22]), .I1(n306[22]), .CO(n43317));
    SB_LUT4 add_18_23_lut (.I0(GND_net), .I1(n257[21]), .I2(n306[21]), 
            .I3(n43315), .O(n356[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_2 (.CI(GND_net), .I0(n5_adj_4918), .I1(n74), 
            .CO(n44702));
    SB_LUT4 add_5159_21_lut (.I0(GND_net), .I1(n14189[18]), .I2(GND_net), 
            .I3(n44426), .O(n13349[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5319_10_lut (.I0(GND_net), .I1(n17044[7]), .I2(n679), 
            .I3(n44568), .O(n16533[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_20_lut (.I0(GND_net), .I1(n14189[17]), .I2(GND_net), 
            .I3(n44425), .O(n13349[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5179_8_lut (.I0(GND_net), .I1(n14588[5]), .I2(n521_adj_4951), 
            .I3(n44647), .O(n13789[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_10 (.CI(n44568), .I0(n17044[7]), .I1(n679), .CO(n44569));
    SB_CARRY add_5159_20 (.CI(n44425), .I0(n14189[17]), .I1(GND_net), 
            .CO(n44426));
    SB_CARRY add_18_23 (.CI(n43315), .I0(n257[21]), .I1(n306[21]), .CO(n43316));
    SB_LUT4 add_5159_19_lut (.I0(GND_net), .I1(n14189[16]), .I2(GND_net), 
            .I3(n44424), .O(n13349[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_22_lut (.I0(GND_net), .I1(n257[20]), .I2(n306[20]), 
            .I3(n43314), .O(n356[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_19 (.CI(n44424), .I0(n14189[16]), .I1(GND_net), 
            .CO(n44425));
    SB_LUT4 i1_2_lut (.I0(counter[23]), .I1(counter[24]), .I2(GND_net), 
            .I3(GND_net), .O(n18));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_18_22 (.CI(n43314), .I0(n257[20]), .I1(n306[20]), .CO(n43315));
    SB_LUT4 add_5159_18_lut (.I0(GND_net), .I1(n14189[15]), .I2(GND_net), 
            .I3(n44423), .O(n13349[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_21_lut (.I0(GND_net), .I1(n257[19]), .I2(n306[19]), 
            .I3(n43313), .O(n356[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5319_9_lut (.I0(GND_net), .I1(n17044[6]), .I2(n606), .I3(n44567), 
            .O(n16533[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[1]), 
            .I3(counter[3]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_5096_23_lut (.I0(GND_net), .I1(n12908[20]), .I2(GND_net), 
            .I3(n44701), .O(n11938[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_21 (.CI(n43313), .I0(n257[19]), .I1(n306[19]), .CO(n43314));
    SB_DFF control_update_37 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3995));   // verilog/motorControl.v(25[10] 32[6])
    SB_CARRY add_5159_18 (.CI(n44423), .I0(n14189[15]), .I1(GND_net), 
            .CO(n44424));
    SB_CARRY add_5319_9 (.CI(n44567), .I0(n17044[6]), .I1(n606), .CO(n44568));
    SB_LUT4 i6_4_lut (.I0(counter[5]), .I1(n12), .I2(counter[2]), .I3(counter[0]), 
            .O(n50434));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(counter[15]), .I1(counter[19]), .I2(counter[25]), 
            .I3(n18), .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_18_20_lut (.I0(GND_net), .I1(n257[18]), .I2(n306[18]), 
            .I3(n43312), .O(n356[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_17_lut (.I0(GND_net), .I1(n14189[14]), .I2(GND_net), 
            .I3(n44422), .O(n13349[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_8 (.CI(n44647), .I0(n14588[5]), .I1(n521_adj_4951), 
            .CO(n44648));
    SB_LUT4 add_5319_8_lut (.I0(GND_net), .I1(n17044[5]), .I2(n533), .I3(n44566), 
            .O(n16533[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_17 (.CI(n44422), .I0(n14189[14]), .I1(GND_net), 
            .CO(n44423));
    SB_LUT4 add_5159_16_lut (.I0(GND_net), .I1(n14189[13]), .I2(n1105_adj_4947), 
            .I3(n44421), .O(n13349[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_20 (.CI(n43312), .I0(n257[18]), .I1(n306[18]), .CO(n43313));
    SB_LUT4 add_5096_22_lut (.I0(GND_net), .I1(n12908[19]), .I2(GND_net), 
            .I3(n44700), .O(n11938[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5179_7_lut (.I0(GND_net), .I1(n14588[4]), .I2(n448_adj_4946), 
            .I3(n44646), .O(n13789[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_19_lut (.I0(GND_net), .I1(n257[17]), .I2(n306[17]), 
            .I3(n43311), .O(n356[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_16 (.CI(n44421), .I0(n14189[13]), .I1(n1105_adj_4947), 
            .CO(n44422));
    SB_LUT4 add_5159_15_lut (.I0(GND_net), .I1(n14189[12]), .I2(n1032_adj_4945), 
            .I3(n44420), .O(n13349[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_19 (.CI(n43311), .I0(n257[17]), .I1(n306[17]), .CO(n43312));
    SB_LUT4 add_18_18_lut (.I0(GND_net), .I1(n257[16]), .I2(n306[16]), 
            .I3(n43310), .O(n356[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_8 (.CI(n44566), .I0(n17044[5]), .I1(n533), .CO(n44567));
    SB_CARRY add_5159_15 (.CI(n44420), .I0(n14189[12]), .I1(n1032_adj_4945), 
            .CO(n44421));
    SB_LUT4 i11_4_lut (.I0(counter[21]), .I1(counter[27]), .I2(counter[26]), 
            .I3(counter[30]), .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(counter[20]), .I1(counter[22]), .I2(counter[14]), 
            .I3(counter[18]), .O(n29_adj_4953));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(counter[29]), .I1(counter[28]), .I2(counter[17]), 
            .I3(counter[16]), .O(n27));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_5096_22 (.CI(n44700), .I0(n12908[19]), .I1(GND_net), 
            .CO(n44701));
    SB_LUT4 i4_4_lut (.I0(counter[13]), .I1(counter[9]), .I2(counter[10]), 
            .I3(counter[11]), .O(n10_adj_4954));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i3_4_lut (.I0(counter[12]), .I1(n50434), .I2(counter[8]), 
            .I3(counter[7]), .O(n9_adj_4955));
    defparam i3_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29_adj_4953), .I2(n28), .I3(n30), 
            .O(n50533));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_18_18 (.CI(n43310), .I0(n257[16]), .I1(n306[16]), .CO(n43311));
    SB_LUT4 add_5159_14_lut (.I0(GND_net), .I1(n14189[11]), .I2(n959_adj_4944), 
            .I3(n44419), .O(n13349[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_14 (.CI(n44419), .I0(n14189[11]), .I1(n959_adj_4944), 
            .CO(n44420));
    SB_LUT4 add_5319_7_lut (.I0(GND_net), .I1(n17044[4]), .I2(n460), .I3(n44565), 
            .O(n16533[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21899_4_lut (.I0(n50533), .I1(counter[31]), .I2(n9_adj_4955), 
            .I3(n10_adj_4954), .O(counter_31__N_3995));   // verilog/motorControl.v(28[8:41])
    defparam i21899_4_lut.LUT_INIT = 16'h3222;
    SB_CARRY add_5319_7 (.CI(n44565), .I0(n17044[4]), .I1(n460), .CO(n44566));
    SB_LUT4 add_5159_13_lut (.I0(GND_net), .I1(n14189[10]), .I2(n886_adj_4943), 
            .I3(n44418), .O(n13349[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5319_6_lut (.I0(GND_net), .I1(n17044[3]), .I2(n387), .I3(n44564), 
            .O(n16533[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5159_13 (.CI(n44418), .I0(n14189[10]), .I1(n886_adj_4943), 
            .CO(n44419));
    SB_LUT4 add_18_17_lut (.I0(GND_net), .I1(n257[15]), .I2(n306[15]), 
            .I3(n43309), .O(n356[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_12_lut (.I0(GND_net), .I1(n14189[9]), .I2(n813_adj_4941), 
            .I3(n44417), .O(n13349[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_17 (.CI(n43309), .I0(n257[15]), .I1(n306[15]), .CO(n43310));
    SB_LUT4 mult_16_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4951));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5096_21_lut (.I0(GND_net), .I1(n12908[18]), .I2(GND_net), 
            .I3(n44699), .O(n11938[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_6 (.CI(n44564), .I0(n17044[3]), .I1(n387), .CO(n44565));
    SB_LUT4 mult_16_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i4_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n181), .I3(GND_net), 
            .O(n207[3]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4956));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i4_3_lut (.I0(n207[3]), .I1(IntegralLimit[3]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [3]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_18_16_lut (.I0(GND_net), .I1(n257[14]), .I2(n306[14]), 
            .I3(n43308), .O(n356[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_16 (.CI(n43308), .I0(n257[14]), .I1(n306[14]), .CO(n43309));
    SB_LUT4 mult_17_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4949));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i8_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5179_7 (.CI(n44646), .I0(n14588[4]), .I1(n448_adj_4946), 
            .CO(n44647));
    SB_CARRY add_5096_21 (.CI(n44699), .I0(n12908[18]), .I1(GND_net), 
            .CO(n44700));
    SB_LUT4 add_18_15_lut (.I0(GND_net), .I1(n257[13]), .I2(n306[13]), 
            .I3(n43307), .O(n356[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_12 (.CI(n44417), .I0(n14189[9]), .I1(n813_adj_4941), 
            .CO(n44418));
    SB_CARRY add_18_15 (.CI(n43307), .I0(n257[13]), .I1(n306[13]), .CO(n43308));
    SB_LUT4 add_18_14_lut (.I0(GND_net), .I1(n257[12]), .I2(n306[12]), 
            .I3(n43306), .O(n356[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_11_lut (.I0(GND_net), .I1(n14189[8]), .I2(n740_adj_4936), 
            .I3(n44416), .O(n13349[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_11 (.CI(n44416), .I0(n14189[8]), .I1(n740_adj_4936), 
            .CO(n44417));
    SB_LUT4 add_5179_6_lut (.I0(GND_net), .I1(n14588[3]), .I2(n375_adj_4935), 
            .I3(n44645), .O(n13789[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_6 (.CI(n44645), .I0(n14588[3]), .I1(n375_adj_4935), 
            .CO(n44646));
    SB_LUT4 add_5319_5_lut (.I0(GND_net), .I1(n17044[2]), .I2(n314), .I3(n44563), 
            .O(n16533[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_5 (.CI(n44563), .I0(n17044[2]), .I1(n314), .CO(n44564));
    SB_LUT4 add_5159_10_lut (.I0(GND_net), .I1(n14189[7]), .I2(n667_adj_4934), 
            .I3(n44415), .O(n13349[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_14 (.CI(n43306), .I0(n257[12]), .I1(n306[12]), .CO(n43307));
    SB_LUT4 mult_17_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4960));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i114_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5159_10 (.CI(n44415), .I0(n14189[7]), .I1(n667_adj_4934), 
            .CO(n44416));
    SB_LUT4 add_5159_9_lut (.I0(GND_net), .I1(n14189[6]), .I2(n594_adj_4933), 
            .I3(n44414), .O(n13349[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5319_4_lut (.I0(GND_net), .I1(n17044[1]), .I2(n241), .I3(n44562), 
            .O(n16533[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5159_9 (.CI(n44414), .I0(n14189[6]), .I1(n594_adj_4933), 
            .CO(n44415));
    SB_LUT4 add_18_13_lut (.I0(GND_net), .I1(n257[11]), .I2(n306[11]), 
            .I3(n43305), .O(n356[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_13 (.CI(n43305), .I0(n257[11]), .I1(n306[11]), .CO(n43306));
    SB_LUT4 add_5096_20_lut (.I0(GND_net), .I1(n12908[17]), .I2(GND_net), 
            .I3(n44698), .O(n11938[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5179_5_lut (.I0(GND_net), .I1(n14588[2]), .I2(n302_adj_4930), 
            .I3(n44644), .O(n13789[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_4 (.CI(n44562), .I0(n17044[1]), .I1(n241), .CO(n44563));
    SB_LUT4 add_5159_8_lut (.I0(GND_net), .I1(n14189[5]), .I2(n521), .I3(n44413), 
            .O(n13349[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_8 (.CI(n44413), .I0(n14189[5]), .I1(n521), .CO(n44414));
    SB_LUT4 add_5159_7_lut (.I0(GND_net), .I1(n14189[4]), .I2(n448), .I3(n44412), 
            .O(n13349[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_5 (.CI(n44644), .I0(n14588[2]), .I1(n302_adj_4930), 
            .CO(n44645));
    SB_LUT4 add_5319_3_lut (.I0(GND_net), .I1(n17044[0]), .I2(n168), .I3(n44561), 
            .O(n16533[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_7 (.CI(n44412), .I0(n14189[4]), .I1(n448), .CO(n44413));
    SB_LUT4 mult_17_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_18_12_lut (.I0(GND_net), .I1(n257[10]), .I2(n306[10]), 
            .I3(n43304), .O(n356[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i506_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_12 (.CI(n43304), .I0(n257[10]), .I1(n306[10]), .CO(n43305));
    SB_LUT4 add_5159_6_lut (.I0(GND_net), .I1(n14189[3]), .I2(n375), .I3(n44411), 
            .O(n13349[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4962));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i120_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5159_6 (.CI(n44411), .I0(n14189[3]), .I1(n375), .CO(n44412));
    SB_LUT4 add_18_11_lut (.I0(GND_net), .I1(n257[9]), .I2(n306[9]), .I3(n43303), 
            .O(n356[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_20 (.CI(n44698), .I0(n12908[17]), .I1(GND_net), 
            .CO(n44699));
    SB_LUT4 add_5159_5_lut (.I0(GND_net), .I1(n14189[2]), .I2(n302_adj_4926), 
            .I3(n44410), .O(n13349[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5179_4_lut (.I0(GND_net), .I1(n14588[1]), .I2(n229_adj_4925), 
            .I3(n44643), .O(n13789[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5096_19_lut (.I0(GND_net), .I1(n12908[16]), .I2(GND_net), 
            .I3(n44697), .O(n11938[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_3 (.CI(n44561), .I0(n17044[0]), .I1(n168), .CO(n44562));
    SB_CARRY add_5179_4 (.CI(n44643), .I0(n14588[1]), .I1(n229_adj_4925), 
            .CO(n44644));
    SB_LUT4 add_5179_3_lut (.I0(GND_net), .I1(n14588[0]), .I2(n156_adj_4924), 
            .I3(n44642), .O(n13789[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5319_2_lut (.I0(GND_net), .I1(n26_adj_4923), .I2(n95_adj_4921), 
            .I3(GND_net), .O(n16533[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5319_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5319_2 (.CI(GND_net), .I0(n26_adj_4923), .I1(n95_adj_4921), 
            .CO(n44561));
    SB_LUT4 add_5349_16_lut (.I0(GND_net), .I1(n17493[13]), .I2(n1120), 
            .I3(n44560), .O(n17044[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_5 (.CI(n44410), .I0(n14189[2]), .I1(n302_adj_4926), 
            .CO(n44411));
    SB_LUT4 add_5159_4_lut (.I0(GND_net), .I1(n14189[1]), .I2(n229), .I3(n44409), 
            .O(n13349[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_4 (.CI(n44409), .I0(n14189[1]), .I1(n229), .CO(n44410));
    SB_CARRY add_18_11 (.CI(n43303), .I0(n257[9]), .I1(n306[9]), .CO(n43304));
    SB_LUT4 add_5159_3_lut (.I0(GND_net), .I1(n14189[0]), .I2(n156), .I3(n44408), 
            .O(n13349[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5349_15_lut (.I0(GND_net), .I1(n17493[12]), .I2(n1047), 
            .I3(n44559), .O(n17044[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i51_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5159_3 (.CI(n44408), .I0(n14189[0]), .I1(n156), .CO(n44409));
    SB_LUT4 add_5159_2_lut (.I0(GND_net), .I1(n14_adj_4917), .I2(n83_adj_4915), 
            .I3(GND_net), .O(n13349[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_2 (.CI(GND_net), .I0(n14_adj_4917), .I1(n83_adj_4915), 
            .CO(n44408));
    SB_LUT4 mult_16_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4918));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5096_19 (.CI(n44697), .I0(n12908[16]), .I1(GND_net), 
            .CO(n44698));
    SB_CARRY add_5179_3 (.CI(n44642), .I0(n14588[0]), .I1(n156_adj_4924), 
            .CO(n44643));
    SB_CARRY add_5349_15 (.CI(n44559), .I0(n17493[12]), .I1(n1047), .CO(n44560));
    SB_LUT4 add_5469_11_lut (.I0(GND_net), .I1(n18948[8]), .I2(n770), 
            .I3(n44407), .O(n18749[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5469_10_lut (.I0(GND_net), .I1(n18948[7]), .I2(n697_adj_4902), 
            .I3(n44406), .O(n18749[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4964));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14757_3_lut (.I0(n356[23]), .I1(n436[23]), .I2(n10863), .I3(GND_net), 
            .O(n28828));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4903));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14762_3_lut (.I0(n356[22]), .I1(n436[22]), .I2(n10863), .I3(GND_net), 
            .O(n28833));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14767_3_lut (.I0(n356[21]), .I1(n436[21]), .I2(n10863), .I3(GND_net), 
            .O(n28838));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14772_3_lut (.I0(n356[20]), .I1(n436[20]), .I2(n10863), .I3(GND_net), 
            .O(n28843));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14777_3_lut (.I0(n356[19]), .I1(n436[19]), .I2(n10863), .I3(GND_net), 
            .O(n28848));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14782_3_lut (.I0(n356[18]), .I1(n436[18]), .I2(n10863), .I3(GND_net), 
            .O(n28853));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14787_3_lut (.I0(n356[17]), .I1(n436[17]), .I2(n10863), .I3(GND_net), 
            .O(n28858));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14792_3_lut (.I0(n356[16]), .I1(n436[16]), .I2(n10863), .I3(GND_net), 
            .O(n28863));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14792_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5469_10 (.CI(n44406), .I0(n18948[7]), .I1(n697_adj_4902), 
            .CO(n44407));
    SB_LUT4 i28813_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n19469[0]), 
            .O(n4_adj_4966));   // verilog/motorControl.v(52[27:38])
    defparam i28813_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i14797_3_lut (.I0(n356[15]), .I1(n436[15]), .I2(n10863), .I3(GND_net), 
            .O(n28868));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14802_3_lut (.I0(n356[14]), .I1(n436[14]), .I2(n10863), .I3(GND_net), 
            .O(n28873));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14807_3_lut (.I0(n356[13]), .I1(n436[13]), .I2(n10863), .I3(GND_net), 
            .O(n28878));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5349_14_lut (.I0(GND_net), .I1(n17493[11]), .I2(n974), 
            .I3(n44558), .O(n17044[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5469_9_lut (.I0(GND_net), .I1(n18948[6]), .I2(n624_adj_4900), 
            .I3(n44405), .O(n18749[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_10_lut (.I0(GND_net), .I1(n257[8]), .I2(n306[8]), .I3(n43302), 
            .O(n356[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5469_9 (.CI(n44405), .I0(n18948[6]), .I1(n624_adj_4900), 
            .CO(n44406));
    SB_CARRY add_5349_14 (.CI(n44558), .I0(n17493[11]), .I1(n974), .CO(n44559));
    SB_LUT4 add_5469_8_lut (.I0(GND_net), .I1(n18948[5]), .I2(n551_adj_4899), 
            .I3(n44404), .O(n18749[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5469_8 (.CI(n44404), .I0(n18948[5]), .I1(n551_adj_4899), 
            .CO(n44405));
    SB_CARRY add_18_10 (.CI(n43302), .I0(n257[8]), .I1(n306[8]), .CO(n43303));
    SB_LUT4 add_5179_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n13789[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14812_3_lut (.I0(n356[12]), .I1(n436[12]), .I2(n10863), .I3(GND_net), 
            .O(n28883));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5349_13_lut (.I0(GND_net), .I1(n17493[10]), .I2(n901), 
            .I3(n44557), .O(n17044[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5469_7_lut (.I0(GND_net), .I1(n18948[4]), .I2(n478), .I3(n44403), 
            .O(n18749[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5469_7 (.CI(n44403), .I0(n18948[4]), .I1(n478), .CO(n44404));
    SB_LUT4 i14817_3_lut (.I0(n356[11]), .I1(n436[11]), .I2(n10863), .I3(GND_net), 
            .O(n28888));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5096_18_lut (.I0(GND_net), .I1(n12908[15]), .I2(GND_net), 
            .I3(n44696), .O(n11938[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14822_3_lut (.I0(n356[10]), .I1(n436[10]), .I2(n10863), .I3(GND_net), 
            .O(n28893));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5469_6_lut (.I0(GND_net), .I1(n18948[3]), .I2(n405), .I3(n44402), 
            .O(n18749[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14827_3_lut (.I0(n356[9]), .I1(n436[9]), .I2(n10863), .I3(GND_net), 
            .O(n28898));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14827_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5179_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n44642));
    SB_LUT4 i14832_3_lut (.I0(n356[8]), .I1(n436[8]), .I2(n10863), .I3(GND_net), 
            .O(n28903));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14832_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5349_13 (.CI(n44557), .I0(n17493[10]), .I1(n901), .CO(n44558));
    SB_LUT4 i14837_3_lut (.I0(n356[7]), .I1(n436[7]), .I2(n10863), .I3(GND_net), 
            .O(n28908));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5349_12_lut (.I0(GND_net), .I1(n17493[9]), .I2(n828), 
            .I3(n44556), .O(n17044[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5469_6 (.CI(n44402), .I0(n18948[3]), .I1(n405), .CO(n44403));
    SB_LUT4 add_5469_5_lut (.I0(GND_net), .I1(n18948[2]), .I2(n332), .I3(n44401), 
            .O(n18749[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5469_5 (.CI(n44401), .I0(n18948[2]), .I1(n332), .CO(n44402));
    SB_LUT4 i14842_3_lut (.I0(n356[6]), .I1(n436[6]), .I2(n10863), .I3(GND_net), 
            .O(n28913));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5469_4_lut (.I0(GND_net), .I1(n18948[1]), .I2(n259), .I3(n44400), 
            .O(n18749[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_9_lut (.I0(GND_net), .I1(n257[7]), .I2(n306[7]), .I3(n43301), 
            .O(n356[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_18 (.CI(n44696), .I0(n12908[15]), .I1(GND_net), 
            .CO(n44697));
    SB_CARRY add_5469_4 (.CI(n44400), .I0(n18948[1]), .I1(n259), .CO(n44401));
    SB_LUT4 i14847_3_lut (.I0(n356[5]), .I1(n436[5]), .I2(n10863), .I3(GND_net), 
            .O(n28918));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14847_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_18_9 (.CI(n43301), .I0(n257[7]), .I1(n306[7]), .CO(n43302));
    SB_LUT4 i14852_3_lut (.I0(n356[4]), .I1(n436[4]), .I2(n10863), .I3(GND_net), 
            .O(n28923));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[0]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5217_20_lut (.I0(GND_net), .I1(n15309[17]), .I2(GND_net), 
            .I3(n44641), .O(n14588[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5217_19_lut (.I0(GND_net), .I1(n15309[16]), .I2(GND_net), 
            .I3(n44640), .O(n14588[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[1]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14857_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n10863), .I3(GND_net), 
            .O(n28928));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14857_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5349_12 (.CI(n44556), .I0(n17493[9]), .I1(n828), .CO(n44557));
    SB_LUT4 add_5469_3_lut (.I0(GND_net), .I1(n18948[0]), .I2(n186_adj_4897), 
            .I3(n44399), .O(n18749[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5469_3 (.CI(n44399), .I0(n18948[0]), .I1(n186_adj_4897), 
            .CO(n44400));
    SB_LUT4 add_5349_11_lut (.I0(GND_net), .I1(n17493[8]), .I2(n755), 
            .I3(n44555), .O(n17044[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5096_17_lut (.I0(GND_net), .I1(n12908[14]), .I2(GND_net), 
            .I3(n44695), .O(n11938[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_8_lut (.I0(GND_net), .I1(n257[6]), .I2(n306[6]), .I3(n43300), 
            .O(n356[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5469_2_lut (.I0(GND_net), .I1(n44), .I2(n113_adj_4896), 
            .I3(GND_net), .O(n18749[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5469_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_11 (.CI(n44555), .I0(n17493[8]), .I1(n755), .CO(n44556));
    SB_CARRY add_5469_2 (.CI(GND_net), .I0(n44), .I1(n113_adj_4896), .CO(n44399));
    SB_LUT4 add_5198_20_lut (.I0(GND_net), .I1(n14949[17]), .I2(GND_net), 
            .I3(n44398), .O(n14189[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14862_3_lut (.I0(n356[2]), .I1(n436[2]), .I2(n10863), .I3(GND_net), 
            .O(n28933));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[2]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5349_10_lut (.I0(GND_net), .I1(n17493[7]), .I2(n682), 
            .I3(n44554), .O(n17044[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4901));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i202_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5349_10 (.CI(n44554), .I0(n17493[7]), .I1(n682), .CO(n44555));
    SB_LUT4 mult_17_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i39_2_lut (.I0(PWMLimit[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5096_17 (.CI(n44695), .I0(n12908[14]), .I1(GND_net), 
            .CO(n44696));
    SB_LUT4 add_5198_19_lut (.I0(GND_net), .I1(n14949[16]), .I2(GND_net), 
            .I3(n44397), .O(n14189[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_19 (.CI(n44397), .I0(n14949[16]), .I1(GND_net), 
            .CO(n44398));
    SB_LUT4 add_5096_16_lut (.I0(GND_net), .I1(n12908[13]), .I2(n1099), 
            .I3(n44694), .O(n11938[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5198_18_lut (.I0(GND_net), .I1(n14949[15]), .I2(GND_net), 
            .I3(n44396), .O(n14189[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_19 (.CI(n44640), .I0(n15309[16]), .I1(GND_net), 
            .CO(n44641));
    SB_LUT4 add_5217_18_lut (.I0(GND_net), .I1(n15309[15]), .I2(GND_net), 
            .I3(n44639), .O(n14588[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_18 (.CI(n44639), .I0(n15309[15]), .I1(GND_net), 
            .CO(n44640));
    SB_LUT4 add_5349_9_lut (.I0(GND_net), .I1(n17493[6]), .I2(n609), .I3(n44553), 
            .O(n17044[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_18 (.CI(n44396), .I0(n14949[15]), .I1(GND_net), 
            .CO(n44397));
    SB_LUT4 unary_minus_13_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[3]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5198_17_lut (.I0(GND_net), .I1(n14949[14]), .I2(GND_net), 
            .I3(n44395), .O(n14189[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_9 (.CI(n44553), .I0(n17493[6]), .I1(n609), .CO(n44554));
    SB_LUT4 LessThan_23_i41_2_lut (.I0(PWMLimit[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4974));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5198_17 (.CI(n44395), .I0(n14949[14]), .I1(GND_net), 
            .CO(n44396));
    SB_LUT4 add_5217_17_lut (.I0(GND_net), .I1(n15309[14]), .I2(GND_net), 
            .I3(n44638), .O(n14588[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5349_8_lut (.I0(GND_net), .I1(n17493[5]), .I2(n536), .I3(n44552), 
            .O(n17044[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_8 (.CI(n44552), .I0(n17493[5]), .I1(n536), .CO(n44553));
    SB_LUT4 add_5349_7_lut (.I0(GND_net), .I1(n17493[4]), .I2(n463), .I3(n44551), 
            .O(n17044[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5198_16_lut (.I0(GND_net), .I1(n14949[13]), .I2(n1108_adj_4895), 
            .I3(n44394), .O(n14189[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_16 (.CI(n44394), .I0(n14949[13]), .I1(n1108_adj_4895), 
            .CO(n44395));
    SB_CARRY add_5096_16 (.CI(n44694), .I0(n12908[13]), .I1(n1099), .CO(n44695));
    SB_LUT4 LessThan_23_i45_2_lut (.I0(PWMLimit[22]), .I1(n356[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5217_17 (.CI(n44638), .I0(n15309[14]), .I1(GND_net), 
            .CO(n44639));
    SB_CARRY add_5349_7 (.CI(n44551), .I0(n17493[4]), .I1(n463), .CO(n44552));
    SB_LUT4 add_5198_15_lut (.I0(GND_net), .I1(n14949[12]), .I2(n1035_adj_4894), 
            .I3(n44393), .O(n14189[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_15 (.CI(n44393), .I0(n14949[12]), .I1(n1035_adj_4894), 
            .CO(n44394));
    SB_LUT4 add_5198_14_lut (.I0(GND_net), .I1(n14949[11]), .I2(n962_adj_4893), 
            .I3(n44392), .O(n14189[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_14 (.CI(n44392), .I0(n14949[11]), .I1(n962_adj_4893), 
            .CO(n44393));
    SB_LUT4 add_5096_15_lut (.I0(GND_net), .I1(n12908[12]), .I2(n1026), 
            .I3(n44693), .O(n11938[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i43_2_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5217_16_lut (.I0(GND_net), .I1(n15309[13]), .I2(n1108), 
            .I3(n44637), .O(n14588[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_16 (.CI(n44637), .I0(n15309[13]), .I1(n1108), .CO(n44638));
    SB_LUT4 add_5349_6_lut (.I0(GND_net), .I1(n17493[3]), .I2(n390), .I3(n44550), 
            .O(n17044[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i29_2_lut (.I0(PWMLimit[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4975));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i31_2_lut (.I0(PWMLimit[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_13_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[4]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_23_i37_2_lut (.I0(PWMLimit[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i23_2_lut (.I0(PWMLimit[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4976));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i25_2_lut (.I0(PWMLimit[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4977));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i35_2_lut (.I0(PWMLimit[17]), .I1(n356[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4978));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5349_6 (.CI(n44550), .I0(n17493[3]), .I1(n390), .CO(n44551));
    SB_LUT4 add_5198_13_lut (.I0(GND_net), .I1(n14949[10]), .I2(n889_adj_4889), 
            .I3(n44391), .O(n14189[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_13 (.CI(n44391), .I0(n14949[10]), .I1(n889_adj_4889), 
            .CO(n44392));
    SB_LUT4 add_5198_12_lut (.I0(GND_net), .I1(n14949[9]), .I2(n816_adj_4888), 
            .I3(n44390), .O(n14189[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5349_5_lut (.I0(GND_net), .I1(n17493[2]), .I2(n317), .I3(n44549), 
            .O(n17044[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_12 (.CI(n44390), .I0(n14949[9]), .I1(n816_adj_4888), 
            .CO(n44391));
    SB_LUT4 add_5198_11_lut (.I0(GND_net), .I1(n14949[8]), .I2(n743_adj_4887), 
            .I3(n44389), .O(n14189[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_5 (.CI(n44549), .I0(n17493[2]), .I1(n317), .CO(n44550));
    SB_CARRY add_5198_11 (.CI(n44389), .I0(n14949[8]), .I1(n743_adj_4887), 
            .CO(n44390));
    SB_LUT4 add_5217_15_lut (.I0(GND_net), .I1(n15309[12]), .I2(n1035), 
            .I3(n44636), .O(n14588[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_15 (.CI(n44693), .I0(n12908[12]), .I1(n1026), .CO(n44694));
    SB_LUT4 add_5198_10_lut (.I0(GND_net), .I1(n14949[7]), .I2(n670_adj_4886), 
            .I3(n44388), .O(n14189[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5349_4_lut (.I0(GND_net), .I1(n17493[1]), .I2(n244), .I3(n44548), 
            .O(n17044[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_10 (.CI(n44388), .I0(n14949[7]), .I1(n670_adj_4886), 
            .CO(n44389));
    SB_CARRY add_5349_4 (.CI(n44548), .I0(n17493[1]), .I1(n244), .CO(n44549));
    SB_LUT4 add_5349_3_lut (.I0(GND_net), .I1(n17493[0]), .I2(n171), .I3(n44547), 
            .O(n17044[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5198_9_lut (.I0(GND_net), .I1(n14949[6]), .I2(n597_adj_4885), 
            .I3(n44387), .O(n14189[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_9 (.CI(n44387), .I0(n14949[6]), .I1(n597_adj_4885), 
            .CO(n44388));
    SB_CARRY add_5217_15 (.CI(n44636), .I0(n15309[12]), .I1(n1035), .CO(n44637));
    SB_LUT4 add_5217_14_lut (.I0(GND_net), .I1(n15309[11]), .I2(n962), 
            .I3(n44635), .O(n14588[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_3 (.CI(n44547), .I0(n17493[0]), .I1(n171), .CO(n44548));
    SB_LUT4 add_5198_8_lut (.I0(GND_net), .I1(n14949[5]), .I2(n524), .I3(n44386), 
            .O(n14189[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_8 (.CI(n44386), .I0(n14949[5]), .I1(n524), .CO(n44387));
    SB_LUT4 add_5198_7_lut (.I0(GND_net), .I1(n14949[4]), .I2(n451), .I3(n44385), 
            .O(n14189[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_7 (.CI(n44385), .I0(n14949[4]), .I1(n451), .CO(n44386));
    SB_LUT4 add_5096_14_lut (.I0(GND_net), .I1(n12908[11]), .I2(n953), 
            .I3(n44692), .O(n11938[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_14 (.CI(n44635), .I0(n15309[11]), .I1(n962), .CO(n44636));
    SB_CARRY add_5096_14 (.CI(n44692), .I0(n12908[11]), .I1(n953), .CO(n44693));
    SB_LUT4 add_5349_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n17044[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5198_6_lut (.I0(GND_net), .I1(n14949[3]), .I2(n378), .I3(n44384), 
            .O(n14189[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_6 (.CI(n44384), .I0(n14949[3]), .I1(n378), .CO(n44385));
    SB_CARRY add_5349_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n44547));
    SB_LUT4 add_5096_13_lut (.I0(GND_net), .I1(n12908[10]), .I2(n880), 
            .I3(n44691), .O(n11938[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5198_5_lut (.I0(GND_net), .I1(n14949[2]), .I2(n305), .I3(n44383), 
            .O(n14189[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_13 (.CI(n44691), .I0(n12908[10]), .I1(n880), .CO(n44692));
    SB_LUT4 add_5217_13_lut (.I0(GND_net), .I1(n15309[10]), .I2(n889), 
            .I3(n44634), .O(n14588[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_5 (.CI(n44383), .I0(n14949[2]), .I1(n305), .CO(n44384));
    SB_CARRY add_5217_13 (.CI(n44634), .I0(n15309[10]), .I1(n889), .CO(n44635));
    SB_LUT4 i14550_3_lut (.I0(n356[0]), .I1(n436[0]), .I2(n10863), .I3(GND_net), 
            .O(n28621));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5510_8_lut (.I0(GND_net), .I1(n19285[5]), .I2(n560), .I3(n44546), 
            .O(n19173[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5510_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5198_4_lut (.I0(GND_net), .I1(n14949[1]), .I2(n232), .I3(n44382), 
            .O(n14189[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_4 (.CI(n44382), .I0(n14949[1]), .I1(n232), .CO(n44383));
    SB_LUT4 add_5217_12_lut (.I0(GND_net), .I1(n15309[9]), .I2(n816), 
            .I3(n44633), .O(n14588[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5198_3_lut (.I0(GND_net), .I1(n14949[0]), .I2(n159), .I3(n44381), 
            .O(n14189[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5510_7_lut (.I0(GND_net), .I1(n19285[4]), .I2(n487), .I3(n44545), 
            .O(n19173[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5510_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_3 (.CI(n44381), .I0(n14949[0]), .I1(n159), .CO(n44382));
    SB_LUT4 add_5198_2_lut (.I0(GND_net), .I1(n17), .I2(n86), .I3(GND_net), 
            .O(n14189[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_2 (.CI(GND_net), .I0(n17), .I1(n86), .CO(n44381));
    SB_CARRY add_5510_7 (.CI(n44545), .I0(n19285[4]), .I1(n487), .CO(n44546));
    SB_LUT4 LessThan_23_i11_2_lut (.I0(PWMLimit[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4980));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5235_19_lut (.I0(GND_net), .I1(n15633[16]), .I2(GND_net), 
            .I3(n44380), .O(n14949[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i13_2_lut (.I0(PWMLimit[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i15_2_lut (.I0(PWMLimit[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5510_6_lut (.I0(GND_net), .I1(n19285[3]), .I2(n414), .I3(n44544), 
            .O(n19173[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5510_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5235_18_lut (.I0(GND_net), .I1(n15633[15]), .I2(GND_net), 
            .I3(n44379), .O(n14949[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_18 (.CI(n44379), .I0(n15633[15]), .I1(GND_net), 
            .CO(n44380));
    SB_LUT4 mult_16_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4981));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5235_17_lut (.I0(GND_net), .I1(n15633[14]), .I2(GND_net), 
            .I3(n44378), .O(n14949[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5096_12_lut (.I0(GND_net), .I1(n12908[9]), .I2(n807), 
            .I3(n44690), .O(n11938[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n19469[0]), 
            .O(n19429[1]));   // verilog/motorControl.v(52[27:38])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_17_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4982));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5510_6 (.CI(n44544), .I0(n19285[3]), .I1(n414), .CO(n44545));
    SB_LUT4 LessThan_23_i27_2_lut (.I0(PWMLimit[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4983));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i33_2_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i9_2_lut (.I0(PWMLimit[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4984));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i17_2_lut (.I0(PWMLimit[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4985));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i19_2_lut (.I0(PWMLimit[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i21_2_lut (.I0(PWMLimit[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4986));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5235_17 (.CI(n44378), .I0(n15633[14]), .I1(GND_net), 
            .CO(n44379));
    SB_LUT4 mult_16_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4987));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38674_4_lut (.I0(n21_adj_4986), .I1(n19), .I2(n17_adj_4985), 
            .I3(n9_adj_4984), .O(n54467));
    defparam i38674_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_13_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[5]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5217_12 (.CI(n44633), .I0(n15309[9]), .I1(n816), .CO(n44634));
    SB_LUT4 i38645_4_lut (.I0(n27_adj_4983), .I1(n15), .I2(n13), .I3(n11_adj_4980), 
            .O(n54438));
    defparam i38645_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5510_5_lut (.I0(GND_net), .I1(n19285[2]), .I2(n341), .I3(n44543), 
            .O(n19173[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5510_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_12 (.CI(n44690), .I0(n12908[9]), .I1(n807), .CO(n44691));
    SB_LUT4 add_5096_11_lut (.I0(GND_net), .I1(n12908[8]), .I2(n734), 
            .I3(n44689), .O(n11938[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5217_11_lut (.I0(GND_net), .I1(n15309[8]), .I2(n743), 
            .I3(n44632), .O(n14588[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_11 (.CI(n44632), .I0(n15309[8]), .I1(n743), .CO(n44633));
    SB_LUT4 add_5235_16_lut (.I0(GND_net), .I1(n15633[13]), .I2(n1111), 
            .I3(n44377), .O(n14949[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_11 (.CI(n44689), .I0(n12908[8]), .I1(n734), .CO(n44690));
    SB_LUT4 unary_minus_13_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[6]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5096_10_lut (.I0(GND_net), .I1(n12908[7]), .I2(n661), 
            .I3(n44688), .O(n11938[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5217_10_lut (.I0(GND_net), .I1(n15309[7]), .I2(n670), 
            .I3(n44631), .O(n14588[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5510_5 (.CI(n44543), .I0(n19285[2]), .I1(n341), .CO(n44544));
    SB_LUT4 add_5510_4_lut (.I0(GND_net), .I1(n19285[1]), .I2(n268), .I3(n44542), 
            .O(n19173[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5510_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(counter[31]), 
            .I3(n44109), .O(n34[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(counter[30]), 
            .I3(n44108), .O(n34[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5510_4 (.CI(n44542), .I0(n19285[1]), .I1(n268), .CO(n44543));
    SB_CARRY counter_2283_add_4_32 (.CI(n44108), .I0(GND_net), .I1(counter[30]), 
            .CO(n44109));
    SB_LUT4 mult_16_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4992));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i12_3_lut (.I0(n356[7]), .I1(n356[16]), .I2(n33), 
            .I3(GND_net), .O(n12_adj_4993));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5217_10 (.CI(n44631), .I0(n15309[7]), .I1(n670), .CO(n44632));
    SB_CARRY add_5235_16 (.CI(n44377), .I0(n15633[13]), .I1(n1111), .CO(n44378));
    SB_LUT4 LessThan_23_i10_3_lut (.I0(n356[5]), .I1(n356[6]), .I2(n13), 
            .I3(GND_net), .O(n10_adj_4994));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i30_3_lut (.I0(n12_adj_4993), .I1(n356[17]), .I2(n35_adj_4978), 
            .I3(GND_net), .O(n30_adj_4995));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5235_15_lut (.I0(GND_net), .I1(n15633[12]), .I2(n1038), 
            .I3(n44376), .O(n14949[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(counter[29]), 
            .I3(n44107), .O(n34[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_15 (.CI(n44376), .I0(n15633[12]), .I1(n1038), .CO(n44377));
    SB_LUT4 add_5235_14_lut (.I0(GND_net), .I1(n15633[11]), .I2(n965), 
            .I3(n44375), .O(n14949[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5510_3_lut (.I0(GND_net), .I1(n19285[0]), .I2(n195), .I3(n44541), 
            .O(n19173[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5510_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_14 (.CI(n44375), .I0(n15633[11]), .I1(n965), .CO(n44376));
    SB_CARRY add_5510_3 (.CI(n44541), .I0(n19285[0]), .I1(n195), .CO(n44542));
    SB_LUT4 i39088_4_lut (.I0(n13), .I1(n11_adj_4980), .I2(n9_adj_4984), 
            .I3(n54484), .O(n54881));
    defparam i39088_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY counter_2283_add_4_31 (.CI(n44107), .I0(GND_net), .I1(counter[29]), 
            .CO(n44108));
    SB_LUT4 add_5235_13_lut (.I0(GND_net), .I1(n15633[10]), .I2(n892), 
            .I3(n44374), .O(n14949[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[7]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39084_4_lut (.I0(n19), .I1(n17_adj_4985), .I2(n15), .I3(n54881), 
            .O(n54877));
    defparam i39084_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39621_4_lut (.I0(n25_adj_4977), .I1(n23_adj_4976), .I2(n21_adj_4986), 
            .I3(n54877), .O(n55414));
    defparam i39621_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_5235_13 (.CI(n44374), .I0(n15633[10]), .I1(n892), .CO(n44375));
    SB_LUT4 counter_2283_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(counter[28]), 
            .I3(n44106), .O(n34[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5235_12_lut (.I0(GND_net), .I1(n15633[9]), .I2(n819), 
            .I3(n44373), .O(n14949[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_30 (.CI(n44106), .I0(GND_net), .I1(counter[28]), 
            .CO(n44107));
    SB_LUT4 counter_2283_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(counter[27]), 
            .I3(n44105), .O(n34[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[8]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5217_9_lut (.I0(GND_net), .I1(n15309[6]), .I2(n597), .I3(n44630), 
            .O(n14588[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_9 (.CI(n44630), .I0(n15309[6]), .I1(n597), .CO(n44631));
    SB_CARRY add_5235_12 (.CI(n44373), .I0(n15633[9]), .I1(n819), .CO(n44374));
    SB_LUT4 unary_minus_13_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[9]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY counter_2283_add_4_29 (.CI(n44105), .I0(GND_net), .I1(counter[27]), 
            .CO(n44106));
    SB_LUT4 unary_minus_13_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[10]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39358_4_lut (.I0(n31), .I1(n29_adj_4975), .I2(n27_adj_4983), 
            .I3(n55414), .O(n55151));
    defparam i39358_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39687_4_lut (.I0(n37), .I1(n35_adj_4978), .I2(n33), .I3(n55151), 
            .O(n55480));
    defparam i39687_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_13_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[11]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5510_2_lut (.I0(GND_net), .I1(n53_adj_5001), .I2(n122_adj_5002), 
            .I3(GND_net), .O(n19173[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5510_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i16_3_lut (.I0(n356[9]), .I1(n356[21]), .I2(n43), 
            .I3(GND_net), .O(n16_adj_5003));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[12]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5510_2 (.CI(GND_net), .I0(n53_adj_5001), .I1(n122_adj_5002), 
            .CO(n44541));
    SB_LUT4 add_5235_11_lut (.I0(GND_net), .I1(n15633[8]), .I2(n746), 
            .I3(n44372), .O(n14949[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(counter[26]), 
            .I3(n44104), .O(n34[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_11 (.CI(n44372), .I0(n15633[8]), .I1(n746), .CO(n44373));
    SB_CARRY counter_2283_add_4_28 (.CI(n44104), .I0(GND_net), .I1(counter[26]), 
            .CO(n44105));
    SB_LUT4 counter_2283_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(counter[25]), 
            .I3(n44103), .O(n34[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[13]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39493_3_lut (.I0(n6_adj_5006), .I1(n356[10]), .I2(n21_adj_4986), 
            .I3(GND_net), .O(n55286));   // verilog/motorControl.v(54[14:29])
    defparam i39493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39494_3_lut (.I0(n55286), .I1(n356[11]), .I2(n23_adj_4976), 
            .I3(GND_net), .O(n55287));   // verilog/motorControl.v(54[14:29])
    defparam i39494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17_adj_4985), 
            .I3(GND_net), .O(n8_adj_5007));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5235_10_lut (.I0(GND_net), .I1(n15633[7]), .I2(n673), 
            .I3(n44371), .O(n14949[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_27 (.CI(n44103), .I0(GND_net), .I1(counter[25]), 
            .CO(n44104));
    SB_LUT4 LessThan_23_i24_3_lut (.I0(n16_adj_5003), .I1(n356[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_5008));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38612_4_lut (.I0(n43), .I1(n25_adj_4977), .I2(n23_adj_4976), 
            .I3(n54467), .O(n54405));
    defparam i38612_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39354_4_lut (.I0(n24_adj_5008), .I1(n8_adj_5007), .I2(n45), 
            .I3(n54400), .O(n55147));   // verilog/motorControl.v(54[14:29])
    defparam i39354_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39075_3_lut (.I0(n55287), .I1(n356[12]), .I2(n25_adj_4977), 
            .I3(GND_net), .O(n54868));   // verilog/motorControl.v(54[14:29])
    defparam i39075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_5009));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i4_4_lut (.I0(PWMLimit[0]), .I1(n356[1]), .I2(PWMLimit[1]), 
            .I3(n356[0]), .O(n4_adj_5010));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_17_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5011));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_5012));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2283_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(counter[24]), 
            .I3(n44102), .O(n34[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39567_3_lut (.I0(n4_adj_5010), .I1(n356[13]), .I2(n27_adj_4983), 
            .I3(GND_net), .O(n55360));   // verilog/motorControl.v(54[14:29])
    defparam i39567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5014));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[14]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[15]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39568_3_lut (.I0(n55360), .I1(n356[14]), .I2(n29_adj_4975), 
            .I3(GND_net), .O(n55361));   // verilog/motorControl.v(54[14:29])
    defparam i39568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38635_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4975), .I3(n54438), 
            .O(n54428));
    defparam i38635_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39707_4_lut (.I0(n30_adj_4995), .I1(n10_adj_4994), .I2(n35_adj_4978), 
            .I3(n54426), .O(n55500));   // verilog/motorControl.v(54[14:29])
    defparam i39707_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39484_3_lut (.I0(n55361), .I1(n356[15]), .I2(n31), .I3(GND_net), 
            .O(n55277));   // verilog/motorControl.v(54[14:29])
    defparam i39484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[16]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5217_8_lut (.I0(GND_net), .I1(n15309[5]), .I2(n524_adj_5018), 
            .I3(n44629), .O(n14588[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_10 (.CI(n44371), .I0(n15633[7]), .I1(n673), .CO(n44372));
    SB_LUT4 i39779_4_lut (.I0(n55277), .I1(n55500), .I2(n35_adj_4978), 
            .I3(n54428), .O(n55572));   // verilog/motorControl.v(54[14:29])
    defparam i39779_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5235_9_lut (.I0(GND_net), .I1(n15633[6]), .I2(n600), .I3(n44370), 
            .O(n14949[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5377_15_lut (.I0(GND_net), .I1(n17884[12]), .I2(n1050), 
            .I3(n44540), .O(n17493[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_9 (.CI(n44370), .I0(n15633[6]), .I1(n600), .CO(n44371));
    SB_LUT4 add_5377_14_lut (.I0(GND_net), .I1(n17884[11]), .I2(n977), 
            .I3(n44539), .O(n17493[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39780_3_lut (.I0(n55572), .I1(n356[18]), .I2(n37), .I3(GND_net), 
            .O(n55573));   // verilog/motorControl.v(54[14:29])
    defparam i39780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39760_3_lut (.I0(n55573), .I1(n356[19]), .I2(n39), .I3(GND_net), 
            .O(n55553));   // verilog/motorControl.v(54[14:29])
    defparam i39760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[17]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38614_4_lut (.I0(n43), .I1(n41_adj_4974), .I2(n39), .I3(n55480), 
            .O(n54407));
    defparam i38614_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_5020));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39609_4_lut (.I0(n54868), .I1(n55147), .I2(n45), .I3(n54405), 
            .O(n55402));   // verilog/motorControl.v(54[14:29])
    defparam i39609_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39722_3_lut (.I0(n55553), .I1(n356[20]), .I2(n41_adj_4974), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(54[14:29])
    defparam i39722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39611_4_lut (.I0(n40), .I1(n55402), .I2(n45), .I3(n54407), 
            .O(n55404));   // verilog/motorControl.v(54[14:29])
    defparam i39611_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39612_3_lut (.I0(n55404), .I1(PWMLimit[23]), .I2(n356[23]), 
            .I3(GND_net), .O(n409));   // verilog/motorControl.v(54[14:29])
    defparam i39612_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_13_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[18]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[19]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[20]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_5024));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i100_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_2283_add_4_26 (.CI(n44102), .I0(GND_net), .I1(counter[24]), 
            .CO(n44103));
    SB_LUT4 add_5235_8_lut (.I0(GND_net), .I1(n15633[5]), .I2(n527), .I3(n44369), 
            .O(n14949[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(counter[23]), 
            .I3(n44101), .O(n34[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_8 (.CI(n44369), .I0(n15633[5]), .I1(n527), .CO(n44370));
    SB_CARRY counter_2283_add_4_25 (.CI(n44101), .I0(GND_net), .I1(counter[23]), 
            .CO(n44102));
    SB_LUT4 LessThan_25_i41_2_lut (.I0(n356[20]), .I1(n436[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5026));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_13_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[21]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_25_i39_2_lut (.I0(n356[19]), .I1(n436[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5028));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i45_2_lut (.I0(n356[22]), .I1(n436[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5029));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_13_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[22]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_5031));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5417[23]));   // verilog/motorControl.v(50[22:36])
    defparam unary_minus_13_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_5033));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22469_1_lut (.I0(n356[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36533));   // verilog/motorControl.v(52[18:38])
    defparam i22469_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_25_i43_2_lut (.I0(n356[21]), .I1(n436[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5034));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i37_2_lut (.I0(n356[18]), .I1(n436[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5035));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[0]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i128_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_8 (.CI(n43300), .I0(n257[6]), .I1(n306[6]), .CO(n43301));
    SB_LUT4 mult_17_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i177_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5377_14 (.CI(n44539), .I0(n17884[11]), .I1(n977), .CO(n44540));
    SB_LUT4 counter_2283_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(counter[22]), 
            .I3(n44100), .O(n34[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_24 (.CI(n44100), .I0(GND_net), .I1(counter[22]), 
            .CO(n44101));
    SB_LUT4 LessThan_25_i29_2_lut (.I0(n356[14]), .I1(n436[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5038));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5235_7_lut (.I0(GND_net), .I1(n15633[4]), .I2(n454_adj_5039), 
            .I3(n44368), .O(n14949[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_7 (.CI(n44368), .I0(n15633[4]), .I1(n454_adj_5039), 
            .CO(n44369));
    SB_LUT4 mult_17_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_5040));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2283_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(counter[21]), 
            .I3(n44099), .O(n34[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_7_lut (.I0(GND_net), .I1(n257[5]), .I2(n306[5]), .I3(n43299), 
            .O(n356[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_23 (.CI(n44099), .I0(GND_net), .I1(counter[21]), 
            .CO(n44100));
    SB_LUT4 counter_2283_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(counter[20]), 
            .I3(n44098), .O(n34[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_10 (.CI(n44688), .I0(n12908[7]), .I1(n661), .CO(n44689));
    SB_CARRY counter_2283_add_4_22 (.CI(n44098), .I0(GND_net), .I1(counter[20]), 
            .CO(n44099));
    SB_LUT4 counter_2283_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(counter[19]), 
            .I3(n44097), .O(n34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_21 (.CI(n44097), .I0(GND_net), .I1(counter[19]), 
            .CO(n44098));
    SB_CARRY add_5217_8 (.CI(n44629), .I0(n15309[5]), .I1(n524_adj_5018), 
            .CO(n44630));
    SB_LUT4 add_5235_6_lut (.I0(GND_net), .I1(n15633[3]), .I2(n381), .I3(n44367), 
            .O(n14949[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5377_13_lut (.I0(GND_net), .I1(n17884[10]), .I2(n904), 
            .I3(n44538), .O(n17493[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[1]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 counter_2283_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(counter[18]), 
            .I3(n44096), .O(n34[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_5044));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i31_2_lut (.I0(n356[15]), .I1(n436[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5045));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5235_6 (.CI(n44367), .I0(n15633[3]), .I1(n381), .CO(n44368));
    SB_LUT4 add_5235_5_lut (.I0(GND_net), .I1(n15633[2]), .I2(n308_adj_5046), 
            .I3(n44366), .O(n14949[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_5 (.CI(n44366), .I0(n15633[2]), .I1(n308_adj_5046), 
            .CO(n44367));
    SB_CARRY add_18_7 (.CI(n43299), .I0(n257[5]), .I1(n306[5]), .CO(n43300));
    SB_CARRY counter_2283_add_4_20 (.CI(n44096), .I0(GND_net), .I1(counter[18]), 
            .CO(n44097));
    SB_LUT4 add_18_6_lut (.I0(GND_net), .I1(n257[4]), .I2(n306[4]), .I3(n43298), 
            .O(n356[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_13 (.CI(n44538), .I0(n17884[10]), .I1(n904), .CO(n44539));
    SB_LUT4 add_5377_12_lut (.I0(GND_net), .I1(n17884[9]), .I2(n831), 
            .I3(n44537), .O(n17493[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_12 (.CI(n44537), .I0(n17884[9]), .I1(n831), .CO(n44538));
    SB_LUT4 add_5235_4_lut (.I0(GND_net), .I1(n15633[1]), .I2(n235_adj_5047), 
            .I3(n44365), .O(n14949[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_4 (.CI(n44365), .I0(n15633[1]), .I1(n235_adj_5047), 
            .CO(n44366));
    SB_LUT4 LessThan_25_i23_2_lut (.I0(n356[11]), .I1(n436[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5048));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 counter_2283_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(counter[17]), 
            .I3(n44095), .O(n34[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_19 (.CI(n44095), .I0(GND_net), .I1(counter[17]), 
            .CO(n44096));
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[2]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 counter_2283_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(counter[16]), 
            .I3(n44094), .O(n34[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5235_3_lut (.I0(GND_net), .I1(n15633[0]), .I2(n162_adj_5051), 
            .I3(n44364), .O(n14949[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i25_2_lut (.I0(n356[12]), .I1(n436[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5052));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY counter_2283_add_4_18 (.CI(n44094), .I0(GND_net), .I1(counter[16]), 
            .CO(n44095));
    SB_CARRY add_18_6 (.CI(n43298), .I0(n257[4]), .I1(n306[4]), .CO(n43299));
    SB_CARRY add_5235_3 (.CI(n44364), .I0(n15633[0]), .I1(n162_adj_5051), 
            .CO(n44365));
    SB_LUT4 counter_2283_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(counter[15]), 
            .I3(n44093), .O(n34[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_5054));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i247_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_2283_add_4_17 (.CI(n44093), .I0(GND_net), .I1(counter[15]), 
            .CO(n44094));
    SB_LUT4 add_5377_11_lut (.I0(GND_net), .I1(n17884[8]), .I2(n758), 
            .I3(n44536), .O(n17493[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5235_2_lut (.I0(GND_net), .I1(n20_adj_5055), .I2(n89_adj_5056), 
            .I3(GND_net), .O(n14949[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5096_9_lut (.I0(GND_net), .I1(n12908[6]), .I2(n588), .I3(n44687), 
            .O(n11938[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(counter[14]), 
            .I3(n44092), .O(n34[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[3]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i35_2_lut (.I0(n356[17]), .I1(n436[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5059));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[4]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_25_i33_2_lut (.I0(n356[16]), .I1(n436[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5061));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i11_2_lut (.I0(n356[5]), .I1(n436[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5062));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i13_2_lut (.I0(n356[6]), .I1(n436[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5063));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i15_2_lut (.I0(n356[7]), .I1(n436[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5064));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i27_2_lut (.I0(n356[13]), .I1(n436[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5065));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i9_2_lut (.I0(n356[4]), .I1(n436[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5066));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i17_2_lut (.I0(n356[8]), .I1(n436[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5067));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_5068));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i153_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter_2283__i31 (.Q(counter[31]), .C(clk16MHz), .D(n34[31]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i30 (.Q(counter[30]), .C(clk16MHz), .D(n34[30]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_LUT4 LessThan_25_i19_2_lut (.I0(n356[9]), .I1(n436[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5069));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i21_2_lut (.I0(n356[10]), .I1(n436[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5070));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38587_4_lut (.I0(n21_adj_5070), .I1(n19_adj_5069), .I2(n17_adj_5067), 
            .I3(n9_adj_5066), .O(n54380));
    defparam i38587_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i38579_4_lut (.I0(n27_adj_5065), .I1(n15_adj_5064), .I2(n13_adj_5063), 
            .I3(n11_adj_5062), .O(n54371));
    defparam i38579_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[5]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_25_i12_3_lut (.I0(n436[7]), .I1(n436[16]), .I2(n33_adj_5061), 
            .I3(GND_net), .O(n12_adj_5072));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR counter_2283__i29 (.Q(counter[29]), .C(clk16MHz), .D(n34[29]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i28 (.Q(counter[28]), .C(clk16MHz), .D(n34[28]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i27 (.Q(counter[27]), .C(clk16MHz), .D(n34[27]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i26 (.Q(counter[26]), .C(clk16MHz), .D(n34[26]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i25 (.Q(counter[25]), .C(clk16MHz), .D(n34[25]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i24 (.Q(counter[24]), .C(clk16MHz), .D(n34[24]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i23 (.Q(counter[23]), .C(clk16MHz), .D(n34[23]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i22 (.Q(counter[22]), .C(clk16MHz), .D(n34[22]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i21 (.Q(counter[21]), .C(clk16MHz), .D(n34[21]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i20 (.Q(counter[20]), .C(clk16MHz), .D(n34[20]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i19 (.Q(counter[19]), .C(clk16MHz), .D(n34[19]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i18 (.Q(counter[18]), .C(clk16MHz), .D(n34[18]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i17 (.Q(counter[17]), .C(clk16MHz), .D(n34[17]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i16 (.Q(counter[16]), .C(clk16MHz), .D(n34[16]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i15 (.Q(counter[15]), .C(clk16MHz), .D(n34[15]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i14 (.Q(counter[14]), .C(clk16MHz), .D(n34[14]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i13 (.Q(counter[13]), .C(clk16MHz), .D(n34[13]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i12 (.Q(counter[12]), .C(clk16MHz), .D(n34[12]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i11 (.Q(counter[11]), .C(clk16MHz), .D(n34[11]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i10 (.Q(counter[10]), .C(clk16MHz), .D(n34[10]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i9 (.Q(counter[9]), .C(clk16MHz), .D(n34[9]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i8 (.Q(counter[8]), .C(clk16MHz), .D(n34[8]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i7 (.Q(counter[7]), .C(clk16MHz), .D(n34[7]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i6 (.Q(counter[6]), .C(clk16MHz), .D(n34[6]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i5 (.Q(counter[5]), .C(clk16MHz), .D(n34[5]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i4 (.Q(counter[4]), .C(clk16MHz), .D(n34[4]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i3 (.Q(counter[3]), .C(clk16MHz), .D(n34[3]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i2 (.Q(counter[2]), .C(clk16MHz), .D(n34[2]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_DFFSR counter_2283__i1 (.Q(counter[1]), .C(clk16MHz), .D(n34[1]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_LUT4 LessThan_25_i10_3_lut (.I0(n436[5]), .I1(n436[6]), .I2(n13_adj_5063), 
            .I3(GND_net), .O(n10_adj_5078));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i30_3_lut (.I0(n12_adj_5072), .I1(n436[17]), .I2(n35_adj_5059), 
            .I3(GND_net), .O(n30_adj_5079));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[6]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[7]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[8]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38988_4_lut (.I0(n13_adj_5063), .I1(n11_adj_5062), .I2(n9_adj_5066), 
            .I3(n54398), .O(n54781));
    defparam i38988_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i38981_4_lut (.I0(n19_adj_5069), .I1(n17_adj_5067), .I2(n15_adj_5064), 
            .I3(n54781), .O(n54774));
    defparam i38981_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39587_4_lut (.I0(n25_adj_5052), .I1(n23_adj_5048), .I2(n21_adj_5070), 
            .I3(n54774), .O(n55380));
    defparam i39587_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39326_4_lut (.I0(n31_adj_5045), .I1(n29_adj_5038), .I2(n27_adj_5065), 
            .I3(n55380), .O(n55119));
    defparam i39326_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[9]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i39683_4_lut (.I0(n37_adj_5035), .I1(n35_adj_5059), .I2(n33_adj_5061), 
            .I3(n55119), .O(n55476));
    defparam i39683_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39577_3_lut (.I0(n6_adj_5084), .I1(n436[10]), .I2(n21_adj_5070), 
            .I3(GND_net), .O(n55370));   // verilog/motorControl.v(56[23:39])
    defparam i39577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i16_3_lut (.I0(n436[9]), .I1(n436[21]), .I2(n43_adj_5034), 
            .I3(GND_net), .O(n16_adj_5085));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_2283_add_4_16 (.CI(n44092), .I0(GND_net), .I1(counter[14]), 
            .CO(n44093));
    SB_LUT4 counter_2283_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(counter[13]), 
            .I3(n44091), .O(n34[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_11 (.CI(n44536), .I0(n17884[8]), .I1(n758), .CO(n44537));
    SB_CARRY add_5096_9 (.CI(n44687), .I0(n12908[6]), .I1(n588), .CO(n44688));
    SB_CARRY add_5235_2 (.CI(GND_net), .I0(n20_adj_5055), .I1(n89_adj_5056), 
            .CO(n44364));
    SB_LUT4 add_5217_7_lut (.I0(GND_net), .I1(n15309[4]), .I2(n451_adj_5086), 
            .I3(n44628), .O(n14588[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_7 (.CI(n44628), .I0(n15309[4]), .I1(n451_adj_5086), 
            .CO(n44629));
    SB_LUT4 add_5487_10_lut (.I0(GND_net), .I1(n19109[7]), .I2(n700), 
            .I3(n44363), .O(n18948[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5487_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i8_3_lut (.I0(n436[4]), .I1(n436[8]), .I2(n17_adj_5067), 
            .I3(GND_net), .O(n8_adj_5087));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5096_8_lut (.I0(GND_net), .I1(n12908[5]), .I2(n515), .I3(n44686), 
            .O(n11938[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5487_9_lut (.I0(GND_net), .I1(n19109[6]), .I2(n627), .I3(n44362), 
            .O(n18948[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5487_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i24_3_lut (.I0(n16_adj_5085), .I1(n436[22]), .I2(n45_adj_5029), 
            .I3(GND_net), .O(n24_adj_5088));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39578_3_lut (.I0(n55370), .I1(n436[11]), .I2(n23_adj_5048), 
            .I3(GND_net), .O(n55371));   // verilog/motorControl.v(56[23:39])
    defparam i39578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38561_4_lut (.I0(n43_adj_5034), .I1(n25_adj_5052), .I2(n23_adj_5048), 
            .I3(n54380), .O(n54353));
    defparam i38561_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5377_10_lut (.I0(GND_net), .I1(n17884[7]), .I2(n685), 
            .I3(n44535), .O(n17493[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_10 (.CI(n44535), .I0(n17884[7]), .I1(n685), .CO(n44536));
    SB_CARRY counter_2283_add_4_15 (.CI(n44091), .I0(GND_net), .I1(counter[13]), 
            .CO(n44092));
    SB_LUT4 mult_17_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_5089));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39356_4_lut (.I0(n24_adj_5088), .I1(n8_adj_5087), .I2(n45_adj_5029), 
            .I3(n54351), .O(n55149));   // verilog/motorControl.v(56[23:39])
    defparam i39356_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39488_3_lut (.I0(n55371), .I1(n436[12]), .I2(n25_adj_5052), 
            .I3(GND_net), .O(n55281));   // verilog/motorControl.v(56[23:39])
    defparam i39488_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5487_9 (.CI(n44362), .I0(n19109[6]), .I1(n627), .CO(n44363));
    SB_LUT4 counter_2283_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(counter[12]), 
            .I3(n44090), .O(n34[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5217_6_lut (.I0(GND_net), .I1(n15309[3]), .I2(n378_adj_5090), 
            .I3(n44627), .O(n14588[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i4_4_lut (.I0(n436[0]), .I1(n436[1]), .I2(n356[1]), 
            .I3(n356[0]), .O(n4_adj_5091));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[10]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY counter_2283_add_4_14 (.CI(n44090), .I0(GND_net), .I1(counter[12]), 
            .CO(n44091));
    SB_LUT4 add_5487_8_lut (.I0(GND_net), .I1(n19109[5]), .I2(n554), .I3(n44361), 
            .O(n18948[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5487_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5377_9_lut (.I0(GND_net), .I1(n17884[6]), .I2(n612), .I3(n44534), 
            .O(n17493[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5487_8 (.CI(n44361), .I0(n19109[5]), .I1(n554), .CO(n44362));
    SB_LUT4 add_5487_7_lut (.I0(GND_net), .I1(n19109[4]), .I2(n481), .I3(n44360), 
            .O(n18948[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5487_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_5_lut (.I0(GND_net), .I1(n257[3]), .I2(n306[3]), .I3(n43297), 
            .O(n356[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5487_7 (.CI(n44360), .I0(n19109[4]), .I1(n481), .CO(n44361));
    SB_LUT4 counter_2283_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(counter[11]), 
            .I3(n44089), .O(n34[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39575_3_lut (.I0(n4_adj_5091), .I1(n436[13]), .I2(n27_adj_5065), 
            .I3(GND_net), .O(n55368));   // verilog/motorControl.v(56[23:39])
    defparam i39575_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_2283_add_4_13 (.CI(n44089), .I0(GND_net), .I1(counter[11]), 
            .CO(n44090));
    SB_CARRY add_5217_6 (.CI(n44627), .I0(n15309[3]), .I1(n378_adj_5090), 
            .CO(n44628));
    SB_LUT4 counter_2283_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(counter[10]), 
            .I3(n44088), .O(n34[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_12 (.CI(n44088), .I0(GND_net), .I1(counter[10]), 
            .CO(n44089));
    SB_LUT4 i39576_3_lut (.I0(n55368), .I1(n436[14]), .I2(n29_adj_5038), 
            .I3(GND_net), .O(n55369));   // verilog/motorControl.v(56[23:39])
    defparam i39576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_2283_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(counter[9]), 
            .I3(n44087), .O(n34[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38575_4_lut (.I0(n33_adj_5061), .I1(n31_adj_5045), .I2(n29_adj_5038), 
            .I3(n54371), .O(n54367));
    defparam i38575_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5377_9 (.CI(n44534), .I0(n17884[6]), .I1(n612), .CO(n44535));
    SB_CARRY counter_2283_add_4_11 (.CI(n44087), .I0(GND_net), .I1(counter[9]), 
            .CO(n44088));
    SB_LUT4 mult_16_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_5093));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2283_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(counter[8]), 
            .I3(n44086), .O(n34[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5487_6_lut (.I0(GND_net), .I1(n19109[3]), .I2(n408), .I3(n44359), 
            .O(n18948[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5487_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_10 (.CI(n44086), .I0(GND_net), .I1(counter[8]), 
            .CO(n44087));
    SB_CARRY add_18_5 (.CI(n43297), .I0(n257[3]), .I1(n306[3]), .CO(n43298));
    SB_CARRY add_5487_6 (.CI(n44359), .I0(n19109[3]), .I1(n408), .CO(n44360));
    SB_LUT4 counter_2283_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n44085), .O(n34[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_9 (.CI(n44085), .I0(GND_net), .I1(counter[7]), 
            .CO(n44086));
    SB_LUT4 add_5487_5_lut (.I0(GND_net), .I1(n19109[2]), .I2(n335_adj_5094), 
            .I3(n44358), .O(n18948[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5487_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5217_5_lut (.I0(GND_net), .I1(n15309[2]), .I2(n305_adj_5095), 
            .I3(n44626), .O(n14588[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5377_8_lut (.I0(GND_net), .I1(n17884[5]), .I2(n539), .I3(n44533), 
            .O(n17493[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_8 (.CI(n44533), .I0(n17884[5]), .I1(n539), .CO(n44534));
    SB_LUT4 add_5377_7_lut (.I0(GND_net), .I1(n17884[4]), .I2(n466), .I3(n44532), 
            .O(n17493[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39709_4_lut (.I0(n30_adj_5079), .I1(n10_adj_5078), .I2(n35_adj_5059), 
            .I3(n54365), .O(n55502));   // verilog/motorControl.v(56[23:39])
    defparam i39709_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5487_5 (.CI(n44358), .I0(n19109[2]), .I1(n335_adj_5094), 
            .CO(n44359));
    SB_LUT4 add_5487_4_lut (.I0(GND_net), .I1(n19109[1]), .I2(n262_adj_5096), 
            .I3(n44357), .O(n18948[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5487_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_7 (.CI(n44532), .I0(n17884[4]), .I1(n466), .CO(n44533));
    SB_LUT4 i39490_3_lut (.I0(n55369), .I1(n436[15]), .I2(n31_adj_5045), 
            .I3(GND_net), .O(n55283));   // verilog/motorControl.v(56[23:39])
    defparam i39490_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5487_4 (.CI(n44357), .I0(n19109[1]), .I1(n262_adj_5096), 
            .CO(n44358));
    SB_LUT4 add_5487_3_lut (.I0(GND_net), .I1(n19109[0]), .I2(n189_adj_5097), 
            .I3(n44356), .O(n18948[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5487_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5487_3 (.CI(n44356), .I0(n19109[0]), .I1(n189_adj_5097), 
            .CO(n44357));
    SB_LUT4 counter_2283_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n44084), .O(n34[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_8 (.CI(n44084), .I0(GND_net), .I1(counter[6]), 
            .CO(n44085));
    SB_LUT4 counter_2283_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n44083), .O(n34[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_7 (.CI(n44083), .I0(GND_net), .I1(counter[5]), 
            .CO(n44084));
    SB_LUT4 counter_2283_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n44082), .O(n34[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_8 (.CI(n44686), .I0(n12908[5]), .I1(n515), .CO(n44687));
    SB_LUT4 add_18_4_lut (.I0(GND_net), .I1(n257[2]), .I2(n306[2]), .I3(n43296), 
            .O(n356[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_6 (.CI(n44082), .I0(GND_net), .I1(counter[4]), 
            .CO(n44083));
    SB_CARRY add_5217_5 (.CI(n44626), .I0(n15309[2]), .I1(n305_adj_5095), 
            .CO(n44627));
    SB_LUT4 add_5377_6_lut (.I0(GND_net), .I1(n17884[3]), .I2(n393), .I3(n44531), 
            .O(n17493[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_4 (.CI(n43296), .I0(n257[2]), .I1(n306[2]), .CO(n43297));
    SB_LUT4 counter_2283_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n44081), .O(n34[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5487_2_lut (.I0(GND_net), .I1(n47_adj_5098), .I2(n116_adj_5099), 
            .I3(GND_net), .O(n18948[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5487_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5487_2 (.CI(GND_net), .I0(n47_adj_5098), .I1(n116_adj_5099), 
            .CO(n44356));
    SB_CARRY add_5377_6 (.CI(n44531), .I0(n17884[3]), .I1(n393), .CO(n44532));
    SB_LUT4 add_18_3_lut (.I0(GND_net), .I1(n257[1]), .I2(n306[1]), .I3(n43295), 
            .O(n356[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5270_18_lut (.I0(GND_net), .I1(n16245[15]), .I2(GND_net), 
            .I3(n44355), .O(n15633[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_5 (.CI(n44081), .I0(GND_net), .I1(counter[3]), 
            .CO(n44082));
    SB_LUT4 add_5270_17_lut (.I0(GND_net), .I1(n16245[14]), .I2(GND_net), 
            .I3(n44354), .O(n15633[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n44080), .O(n34[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_17 (.CI(n44354), .I0(n16245[14]), .I1(GND_net), 
            .CO(n44355));
    SB_LUT4 add_5096_7_lut (.I0(GND_net), .I1(n12908[4]), .I2(n442_adj_5100), 
            .I3(n44685), .O(n11938[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_4 (.CI(n44080), .I0(GND_net), .I1(counter[2]), 
            .CO(n44081));
    SB_LUT4 add_5217_4_lut (.I0(GND_net), .I1(n15309[1]), .I2(n232_adj_5101), 
            .I3(n44625), .O(n14588[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2283_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n44079), .O(n34[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2283_add_4_3 (.CI(n44079), .I0(GND_net), .I1(counter[1]), 
            .CO(n44080));
    SB_LUT4 counter_2283_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n34[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2283_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_3 (.CI(n43295), .I0(n257[1]), .I1(n306[1]), .CO(n43296));
    SB_CARRY counter_2283_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n44079));
    SB_LUT4 add_5377_5_lut (.I0(GND_net), .I1(n17884[2]), .I2(n320), .I3(n44530), 
            .O(n17493[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5270_16_lut (.I0(GND_net), .I1(n16245[13]), .I2(n1114_adj_5103), 
            .I3(n44353), .O(n15633[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_2_lut (.I0(GND_net), .I1(n257[0]), .I2(n306[0]), .I3(GND_net), 
            .O(n356[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_16 (.CI(n44353), .I0(n16245[13]), .I1(n1114_adj_5103), 
            .CO(n44354));
    SB_LUT4 add_5270_15_lut (.I0(GND_net), .I1(n16245[12]), .I2(n1041_adj_5105), 
            .I3(n44352), .O(n15633[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_4 (.CI(n44625), .I0(n15309[1]), .I1(n232_adj_5101), 
            .CO(n44626));
    SB_CARRY add_18_2 (.CI(GND_net), .I0(n257[0]), .I1(n306[0]), .CO(n43295));
    SB_LUT4 add_5217_3_lut (.I0(GND_net), .I1(n15309[0]), .I2(n159_adj_5106), 
            .I3(n44624), .O(n14588[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_3 (.CI(n44624), .I0(n15309[0]), .I1(n159_adj_5106), 
            .CO(n44625));
    SB_CARRY add_5270_15 (.CI(n44352), .I0(n16245[12]), .I1(n1041_adj_5105), 
            .CO(n44353));
    SB_LUT4 add_5270_14_lut (.I0(GND_net), .I1(n16245[11]), .I2(n968), 
            .I3(n44351), .O(n15633[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[11]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[12]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5096_7 (.CI(n44685), .I0(n12908[4]), .I1(n442_adj_5100), 
            .CO(n44686));
    SB_LUT4 i39781_4_lut (.I0(n55283), .I1(n55502), .I2(n35_adj_5059), 
            .I3(n54367), .O(n55574));   // verilog/motorControl.v(56[23:39])
    defparam i39781_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5377_5 (.CI(n44530), .I0(n17884[2]), .I1(n320), .CO(n44531));
    SB_LUT4 i39782_3_lut (.I0(n55574), .I1(n436[18]), .I2(n37_adj_5035), 
            .I3(GND_net), .O(n55575));   // verilog/motorControl.v(56[23:39])
    defparam i39782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39758_3_lut (.I0(n55575), .I1(n436[19]), .I2(n39_adj_5028), 
            .I3(GND_net), .O(n55551));   // verilog/motorControl.v(56[23:39])
    defparam i39758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38563_4_lut (.I0(n43_adj_5034), .I1(n41_adj_5026), .I2(n39_adj_5028), 
            .I3(n55476), .O(n54355));
    defparam i38563_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_9_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n1[23]), .I3(n43294), .O(n130[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n1[22]), .I3(n43293), .O(n130[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_14 (.CI(n44351), .I0(n16245[11]), .I1(n968), .CO(n44352));
    SB_LUT4 add_5377_4_lut (.I0(GND_net), .I1(n17884[1]), .I2(n247), .I3(n44529), 
            .O(n17493[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39615_4_lut (.I0(n55281), .I1(n55149), .I2(n45_adj_5029), 
            .I3(n54353), .O(n55408));   // verilog/motorControl.v(56[23:39])
    defparam i39615_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[13]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5270_13_lut (.I0(GND_net), .I1(n16245[10]), .I2(n895), 
            .I3(n44350), .O(n15633[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39724_3_lut (.I0(n55551), .I1(n436[20]), .I2(n41_adj_5026), 
            .I3(GND_net), .O(n40_adj_5110));   // verilog/motorControl.v(56[23:39])
    defparam i39724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39617_4_lut (.I0(n40_adj_5110), .I1(n55408), .I2(n45_adj_5029), 
            .I3(n54355), .O(n55410));   // verilog/motorControl.v(56[23:39])
    defparam i39617_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_5111));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39618_3_lut (.I0(n55410), .I1(n356[23]), .I2(n436[23]), .I3(GND_net), 
            .O(n55411));   // verilog/motorControl.v(56[23:39])
    defparam i39618_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5270_13 (.CI(n44350), .I0(n16245[10]), .I1(n895), .CO(n44351));
    SB_LUT4 add_5270_12_lut (.I0(GND_net), .I1(n16245[9]), .I2(n822), 
            .I3(n44349), .O(n15633[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_5112));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5096_6_lut (.I0(GND_net), .I1(n12908[3]), .I2(n369_adj_5113), 
            .I3(n44684), .O(n11938[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5217_2_lut (.I0(GND_net), .I1(n17_adj_5114), .I2(n86_adj_5115), 
            .I3(GND_net), .O(n14588[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4994_3_lut (.I0(control_update), .I1(n409), .I2(n55411), 
            .I3(GND_net), .O(n10863));   // verilog/motorControl.v(22[7:21])
    defparam i4994_3_lut.LUT_INIT = 16'ha8a8;
    SB_CARRY add_5270_12 (.CI(n44349), .I0(n16245[9]), .I1(n822), .CO(n44350));
    SB_LUT4 add_5270_11_lut (.I0(GND_net), .I1(n16245[8]), .I2(n749), 
            .I3(n44348), .O(n15633[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_2 (.CI(GND_net), .I0(n17_adj_5114), .I1(n86_adj_5115), 
            .CO(n44624));
    SB_CARRY add_5377_4 (.CI(n44529), .I0(n17884[1]), .I1(n247), .CO(n44530));
    SB_CARRY add_9_24 (.CI(n43293), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n1[22]), .CO(n43294));
    SB_LUT4 add_5377_3_lut (.I0(GND_net), .I1(n17884[0]), .I2(n174), .I3(n44528), 
            .O(n17493[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_11 (.CI(n44348), .I0(n16245[8]), .I1(n749), .CO(n44349));
    SB_LUT4 add_5478_10_lut (.I0(GND_net), .I1(n19029[7]), .I2(n700_adj_5116), 
            .I3(n44623), .O(n18849[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5478_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_3 (.CI(n44528), .I0(n17884[0]), .I1(n174), .CO(n44529));
    SB_LUT4 add_5377_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n17493[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5270_10_lut (.I0(GND_net), .I1(n16245[7]), .I2(n676_adj_5117), 
            .I3(n44347), .O(n15633[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_10 (.CI(n44347), .I0(n16245[7]), .I1(n676_adj_5117), 
            .CO(n44348));
    SB_LUT4 add_5270_9_lut (.I0(GND_net), .I1(n16245[6]), .I2(n603_adj_5118), 
            .I3(n44346), .O(n15633[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n1[21]), .I3(n43292), .O(n130[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5478_9_lut (.I0(GND_net), .I1(n19029[6]), .I2(n627_adj_5119), 
            .I3(n44622), .O(n18849[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5478_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n44528));
    SB_CARRY add_5270_9 (.CI(n44346), .I0(n16245[6]), .I1(n603_adj_5118), 
            .CO(n44347));
    SB_LUT4 add_5270_8_lut (.I0(GND_net), .I1(n16245[5]), .I2(n530_adj_5120), 
            .I3(n44345), .O(n15633[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5403_14_lut (.I0(GND_net), .I1(n18221[11]), .I2(n980_adj_5121), 
            .I3(n44527), .O(n17884[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_23 (.CI(n43292), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n1[21]), .CO(n43293));
    SB_LUT4 add_5403_13_lut (.I0(GND_net), .I1(n18221[10]), .I2(n907_adj_5122), 
            .I3(n44526), .O(n17884[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_8 (.CI(n44345), .I0(n16245[5]), .I1(n530_adj_5120), 
            .CO(n44346));
    SB_LUT4 add_5270_7_lut (.I0(GND_net), .I1(n16245[4]), .I2(n457_adj_5123), 
            .I3(n44344), .O(n15633[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_6 (.CI(n44684), .I0(n12908[3]), .I1(n369_adj_5113), 
            .CO(n44685));
    SB_LUT4 add_9_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n1[20]), .I3(n43291), .O(n130[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_22 (.CI(n43291), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n1[20]), .CO(n43292));
    SB_LUT4 add_9_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n1[19]), .I3(n43290), .O(n130[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_7 (.CI(n44344), .I0(n16245[4]), .I1(n457_adj_5123), 
            .CO(n44345));
    SB_CARRY add_9_21 (.CI(n43290), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n1[19]), .CO(n43291));
    SB_LUT4 mult_16_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_5124));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(deadband[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5125));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5270_6_lut (.I0(GND_net), .I1(n16245[3]), .I2(n384_adj_5126), 
            .I3(n44343), .O(n15633[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(deadband[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5127));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(deadband[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5128));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(deadband[17]), .I1(n356[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5129));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(deadband[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5130));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(deadband[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5131));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_9_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n1[18]), .I3(n43289), .O(n130[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_20 (.CI(n43289), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n1[18]), .CO(n43290));
    SB_LUT4 add_9_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n1[17]), .I3(n43288), .O(n130[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_19 (.CI(n43288), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n1[17]), .CO(n43289));
    SB_LUT4 add_9_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n1[16]), .I3(n43287), .O(n130[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(deadband[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5134));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(deadband[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5135));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[14]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_9_18 (.CI(n43287), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n1[16]), .CO(n43288));
    SB_LUT4 add_9_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n1[15]), .I3(n43286), .O(n130[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_17 (.CI(n43286), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n1[15]), .CO(n43287));
    SB_LUT4 add_9_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n1[14]), .I3(n43285), .O(n130[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_16 (.CI(n43285), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n1[14]), .CO(n43286));
    SB_LUT4 add_9_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n1[13]), .I3(n43284), .O(n130[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_15 (.CI(n43284), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n1[13]), .CO(n43285));
    SB_LUT4 mult_16_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i541_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5478_9 (.CI(n44622), .I0(n19029[6]), .I1(n627_adj_5119), 
            .CO(n44623));
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[15]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[16]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_9_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n1[12]), .I3(n43283), .O(n130[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5403_13 (.CI(n44526), .I0(n18221[10]), .I1(n907_adj_5122), 
            .CO(n44527));
    SB_LUT4 LessThan_19_i25_2_lut (.I0(deadband[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5141));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5270_6 (.CI(n44343), .I0(n16245[3]), .I1(n384_adj_5126), 
            .CO(n44344));
    SB_LUT4 LessThan_19_i45_2_lut (.I0(deadband[22]), .I1(n356[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5142));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_5143));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(deadband[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5144));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5270_5_lut (.I0(GND_net), .I1(n16245[2]), .I2(n311_adj_5145), 
            .I3(n44342), .O(n15633[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5096_5_lut (.I0(GND_net), .I1(n12908[2]), .I2(n296_adj_5146), 
            .I3(n44683), .O(n11938[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5478_8_lut (.I0(GND_net), .I1(n19029[5]), .I2(n554_adj_5147), 
            .I3(n44621), .O(n18849[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5478_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5270_5 (.CI(n44342), .I0(n16245[2]), .I1(n311_adj_5145), 
            .CO(n44343));
    SB_LUT4 add_5270_4_lut (.I0(GND_net), .I1(n16245[1]), .I2(n238_adj_5148), 
            .I3(n44341), .O(n15633[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[17]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5270_4 (.CI(n44341), .I0(n16245[1]), .I1(n238_adj_5148), 
            .CO(n44342));
    SB_LUT4 add_5403_12_lut (.I0(GND_net), .I1(n18221[9]), .I2(n834_adj_5150), 
            .I3(n44525), .O(n17884[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5270_3_lut (.I0(GND_net), .I1(n16245[0]), .I2(n165_adj_5151), 
            .I3(n44340), .O(n15633[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_14 (.CI(n43283), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n1[12]), .CO(n43284));
    SB_LUT4 add_9_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n1[11]), .I3(n43282), .O(n130[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_13 (.CI(n43282), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n1[11]), .CO(n43283));
    SB_CARRY add_5096_5 (.CI(n44683), .I0(n12908[2]), .I1(n296_adj_5146), 
            .CO(n44684));
    SB_CARRY add_5478_8 (.CI(n44621), .I0(n19029[5]), .I1(n554_adj_5147), 
            .CO(n44622));
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[18]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_5153));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n1[10]), .I3(n43281), .O(n130[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(deadband[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5155));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5156));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(deadband[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5157));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5096_4_lut (.I0(GND_net), .I1(n12908[1]), .I2(n223_adj_5158), 
            .I3(n44682), .O(n11938[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5403_12 (.CI(n44525), .I0(n18221[9]), .I1(n834_adj_5150), 
            .CO(n44526));
    SB_CARRY add_5270_3 (.CI(n44340), .I0(n16245[0]), .I1(n165_adj_5151), 
            .CO(n44341));
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[19]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(deadband[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5160));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5270_2_lut (.I0(GND_net), .I1(n23_adj_5161), .I2(n92_adj_5162), 
            .I3(GND_net), .O(n15633[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5270_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_5163));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(deadband[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5164));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_9_12 (.CI(n43281), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n1[10]), .CO(n43282));
    SB_LUT4 add_9_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n1[9]), .I3(n43280), .O(n130[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5403_11_lut (.I0(GND_net), .I1(n18221[8]), .I2(n761_adj_5166), 
            .I3(n44524), .O(n17884[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_4 (.CI(n44682), .I0(n12908[1]), .I1(n223_adj_5158), 
            .CO(n44683));
    SB_LUT4 add_5478_7_lut (.I0(GND_net), .I1(n19029[4]), .I2(n481_adj_5167), 
            .I3(n44620), .O(n18849[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5478_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_11 (.CI(n43280), .I0(\PID_CONTROLLER.integral [9]), .I1(n1[9]), 
            .CO(n43281));
    SB_CARRY add_5270_2 (.CI(GND_net), .I0(n23_adj_5161), .I1(n92_adj_5162), 
            .CO(n44340));
    SB_LUT4 add_9_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n1[8]), .I3(n43279), .O(n130[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_10 (.CI(n43279), .I0(\PID_CONTROLLER.integral [8]), .I1(n1[8]), 
            .CO(n43280));
    SB_LUT4 add_5303_17_lut (.I0(GND_net), .I1(n16789[14]), .I2(GND_net), 
            .I3(n44339), .O(n16245[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(deadband[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5168));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(deadband[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5169));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(deadband[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5170));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(deadband[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5171));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38728_4_lut (.I0(n356[8]), .I1(n356[4]), .I2(n382[8]), .I3(n382[4]), 
            .O(n54521));
    defparam i38728_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i39114_3_lut (.I0(n356[9]), .I1(n54521), .I2(n382[9]), .I3(GND_net), 
            .O(n54907));
    defparam i39114_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_21_i21_rep_164_2_lut (.I0(n356[10]), .I1(n382[10]), 
            .I2(GND_net), .I3(GND_net), .O(n56813));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i21_rep_164_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39112_4_lut (.I0(n356[11]), .I1(n56813), .I2(n382[11]), .I3(n54907), 
            .O(n54905));
    defparam i39112_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i25_rep_159_2_lut (.I0(n356[12]), .I1(n382[12]), 
            .I2(GND_net), .I3(GND_net), .O(n56808));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i25_rep_159_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[20]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5303_16_lut (.I0(GND_net), .I1(n16789[13]), .I2(n1117_adj_5174), 
            .I3(n44338), .O(n16245[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_16 (.CI(n44338), .I0(n16789[13]), .I1(n1117_adj_5174), 
            .CO(n44339));
    SB_LUT4 add_9_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n1[7]), .I3(n43278), .O(n130[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5403_11 (.CI(n44524), .I0(n18221[8]), .I1(n761_adj_5166), 
            .CO(n44525));
    SB_LUT4 add_5096_3_lut (.I0(GND_net), .I1(n12908[0]), .I2(n150_adj_5176), 
            .I3(n44681), .O(n11938[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5403_10_lut (.I0(GND_net), .I1(n18221[7]), .I2(n688_adj_5177), 
            .I3(n44523), .O(n17884[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5303_15_lut (.I0(GND_net), .I1(n16789[12]), .I2(n1044_adj_5178), 
            .I3(n44337), .O(n16245[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_9 (.CI(n43278), .I0(\PID_CONTROLLER.integral [7]), .I1(n1[7]), 
            .CO(n43279));
    SB_CARRY add_5303_15 (.CI(n44337), .I0(n16789[12]), .I1(n1044_adj_5178), 
            .CO(n44338));
    SB_CARRY add_5478_7 (.CI(n44620), .I0(n19029[4]), .I1(n481_adj_5167), 
            .CO(n44621));
    SB_CARRY add_5403_10 (.CI(n44523), .I0(n18221[7]), .I1(n688_adj_5177), 
            .CO(n44524));
    SB_LUT4 add_5403_9_lut (.I0(GND_net), .I1(n18221[6]), .I2(n615_adj_5179), 
            .I3(n44522), .O(n17884[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5303_14_lut (.I0(GND_net), .I1(n16789[11]), .I2(n971_adj_5180), 
            .I3(n44336), .O(n16245[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n1[6]), .I3(n43277), .O(n130[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_14 (.CI(n44336), .I0(n16789[11]), .I1(n971_adj_5180), 
            .CO(n44337));
    SB_LUT4 add_5303_13_lut (.I0(GND_net), .I1(n16789[10]), .I2(n898_adj_5182), 
            .I3(n44335), .O(n16245[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_13 (.CI(n44335), .I0(n16789[10]), .I1(n898_adj_5182), 
            .CO(n44336));
    SB_CARRY add_5403_9 (.CI(n44522), .I0(n18221[6]), .I1(n615_adj_5179), 
            .CO(n44523));
    SB_LUT4 add_5478_6_lut (.I0(GND_net), .I1(n19029[3]), .I2(n408_adj_5183), 
            .I3(n44619), .O(n18849[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5478_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5303_12_lut (.I0(GND_net), .I1(n16789[9]), .I2(n825_adj_5184), 
            .I3(n44334), .O(n16245[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5403_8_lut (.I0(GND_net), .I1(n18221[5]), .I2(n542_adj_5185), 
            .I3(n44521), .O(n17884[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5403_8 (.CI(n44521), .I0(n18221[5]), .I1(n542_adj_5185), 
            .CO(n44522));
    SB_LUT4 i1_3_lut_4_lut_adj_1710 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n19501[0]), 
            .I3(n42958), .O(n19484[1]));   // verilog/motorControl.v(52[18:24])
    defparam i1_3_lut_4_lut_adj_1710.LUT_INIT = 16'h8778;
    SB_LUT4 i28897_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n42958), 
            .I3(n19501[0]), .O(n4_adj_4909));   // verilog/motorControl.v(52[18:24])
    defparam i28897_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_17_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_5186));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38760_4_lut (.I0(n27_adj_5171), .I1(n15_adj_5170), .I2(n13_adj_5169), 
            .I3(n11_adj_5168), .O(n54553));
    defparam i38760_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i38767_4_lut (.I0(n21_adj_5164), .I1(n19_adj_5160), .I2(n17_adj_5157), 
            .I3(n9_adj_5155), .O(n54560));
    defparam i38767_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n356[9]), .I1(n356[21]), .I2(n43_adj_5144), 
            .I3(GND_net), .O(n16_adj_5187));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_5188));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i173_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_8 (.CI(n43277), .I0(\PID_CONTROLLER.integral [6]), .I1(n1[6]), 
            .CO(n43278));
    SB_LUT4 mult_16_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_5189));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[21]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17_adj_5157), 
            .I3(GND_net), .O(n8_adj_5191));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_5187), .I1(n356[22]), .I2(n45_adj_5142), 
            .I3(GND_net), .O(n24_adj_5192));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39154_4_lut (.I0(n13_adj_5169), .I1(n11_adj_5168), .I2(n9_adj_5155), 
            .I3(n54571), .O(n54947));
    defparam i39154_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i28884_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n19484[0]));   // verilog/motorControl.v(52[18:24])
    defparam i28884_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i28886_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n42958));   // verilog/motorControl.v(52[18:24])
    defparam i28886_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[22]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_5194));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_5195));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_5196));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39150_4_lut (.I0(n19_adj_5160), .I1(n17_adj_5157), .I2(n15_adj_5170), 
            .I3(n54947), .O(n54943));
    defparam i39150_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_5303_12 (.CI(n44334), .I0(n16789[9]), .I1(n825_adj_5184), 
            .CO(n44335));
    SB_LUT4 add_9_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n1[5]), .I3(n43276), .O(n130[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39641_4_lut (.I0(n25_adj_5141), .I1(n23_adj_5135), .I2(n21_adj_5164), 
            .I3(n54943), .O(n55434));
    defparam i39641_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39390_4_lut (.I0(n31_adj_5134), .I1(n29_adj_5131), .I2(n27_adj_5171), 
            .I3(n55434), .O(n55183));
    defparam i39390_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39699_4_lut (.I0(n37_adj_5130), .I1(n35_adj_5129), .I2(n33_adj_5128), 
            .I3(n55183), .O(n55492));
    defparam i39699_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_9_7 (.CI(n43276), .I0(\PID_CONTROLLER.integral [5]), .I1(n1[5]), 
            .CO(n43277));
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5418[23]));   // verilog/motorControl.v(53[43:52])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_5198));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5303_11_lut (.I0(GND_net), .I1(n16789[8]), .I2(n752_adj_5199), 
            .I3(n44333), .O(n16245[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_5200));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i271_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5096_3 (.CI(n44681), .I0(n12908[0]), .I1(n150_adj_5176), 
            .CO(n44682));
    SB_CARRY add_5478_6 (.CI(n44619), .I0(n19029[3]), .I1(n408_adj_5183), 
            .CO(n44620));
    SB_LUT4 add_9_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n1[4]), .I3(n43275), .O(n130[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5403_7_lut (.I0(GND_net), .I1(n18221[4]), .I2(n469_adj_5201), 
            .I3(n44520), .O(n17884[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_5202));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38732_4_lut (.I0(n356[6]), .I1(n356[5]), .I2(n382[6]), .I3(n382[5]), 
            .O(n54525));
    defparam i38732_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i39118_3_lut (.I0(n356[7]), .I1(n54525), .I2(n382[7]), .I3(GND_net), 
            .O(n54911));
    defparam i39118_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 mult_16_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_5204));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_5205));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i27_rep_152_2_lut (.I0(n356[13]), .I1(n382[13]), 
            .I2(GND_net), .I3(GND_net), .O(n56801));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i27_rep_152_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39106_4_lut (.I0(n356[14]), .I1(n56801), .I2(n382[14]), .I3(n54911), 
            .O(n54899));
    defparam i39106_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i31_rep_146_2_lut (.I0(n356[15]), .I1(n382[15]), 
            .I2(GND_net), .I3(GND_net), .O(n56795));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i31_rep_146_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i12_3_lut (.I0(n382[7]), .I1(n382[16]), .I2(n356[16]), 
            .I3(GND_net), .O(n12_adj_5208));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38708_4_lut (.I0(n356[16]), .I1(n356[7]), .I2(n382[16]), 
            .I3(n382[7]), .O(n54501));
    defparam i38708_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i35_rep_170_2_lut (.I0(n356[17]), .I1(n382[17]), 
            .I2(GND_net), .I3(GND_net), .O(n56819));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i35_rep_170_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_26_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[0]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5303_11 (.CI(n44333), .I0(n16789[8]), .I1(n752_adj_5199), 
            .CO(n44334));
    SB_LUT4 LessThan_21_i10_3_lut (.I0(n382[5]), .I1(n382[6]), .I2(n356[6]), 
            .I3(GND_net), .O(n10_adj_5210));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i30_3_lut (.I0(n12_adj_5208), .I1(n382[17]), .I2(n356[17]), 
            .I3(GND_net), .O(n30_adj_5211));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_16_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_5212));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38736_4_lut (.I0(n356[3]), .I1(n356[2]), .I2(n382[3]), .I3(n382[2]), 
            .O(n54529));
    defparam i38736_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i9_rep_190_2_lut (.I0(n356[4]), .I1(n382[4]), .I2(GND_net), 
            .I3(GND_net), .O(n56839));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i9_rep_190_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_5213));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5214));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[1]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38734_4_lut (.I0(n356[5]), .I1(n56839), .I2(n382[5]), .I3(n54529), 
            .O(n54527));
    defparam i38734_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_5303_10_lut (.I0(GND_net), .I1(n16789[7]), .I2(n679_adj_5216), 
            .I3(n44332), .O(n16245[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[2]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_21_i13_rep_183_2_lut (.I0(n356[6]), .I1(n382[6]), .I2(GND_net), 
            .I3(GND_net), .O(n56832));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i13_rep_183_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_5218));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5096_2_lut (.I0(GND_net), .I1(n8_adj_5214), .I2(n77_adj_5213), 
            .I3(GND_net), .O(n11938[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5096_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39380_4_lut (.I0(n356[7]), .I1(n56832), .I2(n382[7]), .I3(n54527), 
            .O(n55173));
    defparam i39380_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i17_rep_186_2_lut (.I0(n356[8]), .I1(n382[8]), .I2(GND_net), 
            .I3(GND_net), .O(n56835));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i17_rep_186_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_9_6 (.CI(n43275), .I0(\PID_CONTROLLER.integral [4]), .I1(n1[4]), 
            .CO(n43276));
    SB_CARRY add_5303_10 (.CI(n44332), .I0(n16789[7]), .I1(n679_adj_5216), 
            .CO(n44333));
    SB_LUT4 add_9_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n1[3]), .I3(n43274), .O(n130[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[3]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[4]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_5216));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[5]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39116_4_lut (.I0(n356[9]), .I1(n56835), .I2(n382[9]), .I3(n55173), 
            .O(n54909));
    defparam i39116_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i39525_4_lut (.I0(n356[11]), .I1(n56813), .I2(n382[11]), .I3(n54909), 
            .O(n55318));
    defparam i39525_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_5303_9_lut (.I0(GND_net), .I1(n16789[6]), .I2(n606_adj_5205), 
            .I3(n44331), .O(n16245[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_5222));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i418_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5403_7 (.CI(n44520), .I0(n18221[4]), .I1(n469_adj_5201), 
            .CO(n44521));
    SB_LUT4 mult_16_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_5223));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[6]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5403_6_lut (.I0(GND_net), .I1(n18221[3]), .I2(n396_adj_5204), 
            .I3(n44519), .O(n17884[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38720_4_lut (.I0(n356[13]), .I1(n56808), .I2(n382[13]), .I3(n55318), 
            .O(n54513));
    defparam i38720_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_9_5 (.CI(n43274), .I0(\PID_CONTROLLER.integral [3]), .I1(n1[3]), 
            .CO(n43275));
    SB_LUT4 LessThan_21_i29_rep_150_2_lut (.I0(n356[14]), .I1(n382[14]), 
            .I2(GND_net), .I3(GND_net), .O(n56799));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i29_rep_150_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39374_4_lut (.I0(n356[15]), .I1(n56799), .I2(n382[15]), .I3(n54513), 
            .O(n55167));
    defparam i39374_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_9_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n1[2]), .I3(n43273), .O(n130[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_21_i33_rep_175_2_lut (.I0(n356[16]), .I1(n382[16]), 
            .I2(GND_net), .I3(GND_net), .O(n56824));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i33_rep_175_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39629_4_lut (.I0(n356[17]), .I1(n56824), .I2(n382[17]), .I3(n55167), 
            .O(n55422));
    defparam i39629_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 unary_minus_26_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[7]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_5227));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5478_5_lut (.I0(GND_net), .I1(n19029[2]), .I2(n335_adj_5196), 
            .I3(n44618), .O(n18849[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5478_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_5201));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i316_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5403_6 (.CI(n44519), .I0(n18221[3]), .I1(n396_adj_5204), 
            .CO(n44520));
    SB_LUT4 LessThan_21_i37_rep_141_2_lut (.I0(n356[18]), .I1(n382[18]), 
            .I2(GND_net), .I3(GND_net), .O(n56790));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i37_rep_141_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39731_4_lut (.I0(n356[19]), .I1(n56790), .I2(n382[19]), .I3(n55422), 
            .O(n55524));
    defparam i39731_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i41_rep_138_2_lut (.I0(n356[20]), .I1(n382[20]), 
            .I2(GND_net), .I3(GND_net), .O(n56787));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i41_rep_138_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5303_9 (.CI(n44331), .I0(n16789[6]), .I1(n606_adj_5205), 
            .CO(n44332));
    SB_CARRY add_9_4 (.CI(n43273), .I0(\PID_CONTROLLER.integral [2]), .I1(n1[2]), 
            .CO(n43274));
    SB_LUT4 LessThan_21_i6_3_lut (.I0(n382[2]), .I1(n382[3]), .I2(n356[3]), 
            .I3(GND_net), .O(n6_adj_5229));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39501_3_lut (.I0(n6_adj_5229), .I1(n382[10]), .I2(n356[10]), 
            .I3(GND_net), .O(n55294));   // verilog/motorControl.v(53[33:53])
    defparam i39501_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5478_5 (.CI(n44618), .I0(n19029[2]), .I1(n335_adj_5196), 
            .CO(n44619));
    SB_LUT4 add_5403_5_lut (.I0(GND_net), .I1(n18221[2]), .I2(n323_adj_5093), 
            .I3(n44518), .O(n17884[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5096_2 (.CI(GND_net), .I0(n8_adj_5214), .I1(n77_adj_5213), 
            .CO(n44681));
    SB_LUT4 add_5303_8_lut (.I0(GND_net), .I1(n16789[5]), .I2(n533_adj_5089), 
            .I3(n44330), .O(n16245[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[8]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_21_i16_3_lut (.I0(n382[9]), .I1(n382[21]), .I2(n356[21]), 
            .I3(GND_net), .O(n16_adj_5231));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_5232));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i590_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5303_8 (.CI(n44330), .I0(n16789[5]), .I1(n533_adj_5089), 
            .CO(n44331));
    SB_LUT4 mult_16_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_5233));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_5234));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_5199));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[9]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38694_4_lut (.I0(n356[21]), .I1(n356[9]), .I2(n382[21]), 
            .I3(n382[9]), .O(n54487));
    defparam i38694_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 add_9_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n1[1]), .I3(n43272), .O(n130[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_3 (.CI(n43272), .I0(\PID_CONTROLLER.integral [1]), .I1(n1[1]), 
            .CO(n43273));
    SB_LUT4 add_5139_22_lut (.I0(GND_net), .I1(n13789[19]), .I2(GND_net), 
            .I3(n44680), .O(n12908[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n1[0]), .I3(GND_net), .O(n130[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5478_4_lut (.I0(GND_net), .I1(n19029[1]), .I2(n262), .I3(n44617), 
            .O(n18849[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5478_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5478_4 (.CI(n44617), .I0(n19029[1]), .I1(n262), .CO(n44618));
    SB_CARRY add_9_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), .I1(n1[0]), 
            .CO(n43272));
    SB_LUT4 add_5478_3_lut (.I0(GND_net), .I1(n19029[0]), .I2(n189), .I3(n44616), 
            .O(n18849[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5478_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5403_5 (.CI(n44518), .I0(n18221[2]), .I1(n323_adj_5093), 
            .CO(n44519));
    SB_LUT4 LessThan_21_i8_3_lut (.I0(n382[4]), .I1(n382[8]), .I2(n356[8]), 
            .I3(GND_net), .O(n8_adj_5238));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_16_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_5239));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5303_7_lut (.I0(GND_net), .I1(n16789[4]), .I2(n460_adj_5033), 
            .I3(n44329), .O(n16245[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5403_4_lut (.I0(GND_net), .I1(n18221[1]), .I2(n250_adj_5031), 
            .I3(n44517), .O(n17884[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5403_4 (.CI(n44517), .I0(n18221[1]), .I1(n250_adj_5031), 
            .CO(n44518));
    SB_CARRY add_5303_7 (.CI(n44329), .I0(n16789[4]), .I1(n460_adj_5033), 
            .CO(n44330));
    SB_LUT4 add_5303_6_lut (.I0(GND_net), .I1(n16789[3]), .I2(n387_adj_4992), 
            .I3(n44328), .O(n16245[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_6 (.CI(n44328), .I0(n16789[3]), .I1(n387_adj_4992), 
            .CO(n44329));
    SB_LUT4 LessThan_21_i24_3_lut (.I0(n16_adj_5231), .I1(n382[22]), .I2(n356[22]), 
            .I3(GND_net), .O(n24_adj_5241));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5303_5_lut (.I0(GND_net), .I1(n16789[2]), .I2(n314_adj_4982), 
            .I3(n44327), .O(n16245[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5139_21_lut (.I0(GND_net), .I1(n13789[18]), .I2(GND_net), 
            .I3(n44679), .O(n12908[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_5242));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i230_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5139_21 (.CI(n44679), .I0(n13789[18]), .I1(GND_net), 
            .CO(n44680));
    SB_LUT4 mult_16_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_5243));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5139_20_lut (.I0(GND_net), .I1(n13789[17]), .I2(GND_net), 
            .I3(n44678), .O(n12908[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR result__i0 (.Q(duty[0]), .C(clk16MHz), .E(n28830), .D(n28622), 
            .R(n29234));   // verilog/motorControl.v(43[14] 63[8])
    SB_CARRY add_5303_5 (.CI(n44327), .I0(n16789[2]), .I1(n314_adj_4982), 
            .CO(n44328));
    SB_LUT4 i39502_3_lut (.I0(n55294), .I1(n382[11]), .I2(n356[11]), .I3(GND_net), 
            .O(n55295));   // verilog/motorControl.v(53[33:53])
    defparam i39502_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_16_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_5244));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_5245));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38697_4_lut (.I0(n356[21]), .I1(n56808), .I2(n382[21]), .I3(n54905), 
            .O(n54490));
    defparam i38697_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_17_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_5246));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39352_4_lut (.I0(n24_adj_5241), .I1(n8_adj_5238), .I2(n56785), 
            .I3(n54487), .O(n55145));   // verilog/motorControl.v(53[33:53])
    defparam i39352_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_14_i11_3_lut (.I0(n130[10]), .I1(n182[10]), .I2(n181), 
            .I3(GND_net), .O(n207[10]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i11_3_lut (.I0(n207[10]), .I1(IntegralLimit[10]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [10]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_add_1225_24_lut (.I0(n1[23]), .I1(n11938[21]), .I2(GND_net), 
            .I3(n44723), .O(n11431[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_5247));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i69_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5139_20 (.CI(n44678), .I0(n13789[17]), .I1(GND_net), 
            .CO(n44679));
    SB_LUT4 mult_16_add_1225_23_lut (.I0(GND_net), .I1(n11938[20]), .I2(GND_net), 
            .I3(n44722), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_5248));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39065_3_lut (.I0(n55295), .I1(n382[12]), .I2(n356[12]), .I3(GND_net), 
            .O(n54858));   // verilog/motorControl.v(53[33:53])
    defparam i39065_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n356[7]), .I1(n356[16]), .I2(n33_adj_5128), 
            .I3(GND_net), .O(n12_adj_5249));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(deadband[0]), .I1(n356[1]), .I2(deadband[1]), 
            .I3(n356[0]), .O(n4_adj_5250));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i39505_3_lut (.I0(n4_adj_5250), .I1(n356[13]), .I2(n27_adj_5171), 
            .I3(GND_net), .O(n55298));   // verilog/motorControl.v(53[12:29])
    defparam i39505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39506_3_lut (.I0(n55298), .I1(n356[14]), .I2(n29_adj_5131), 
            .I3(GND_net), .O(n55299));   // verilog/motorControl.v(53[12:29])
    defparam i39506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5303_4_lut (.I0(GND_net), .I1(n16789[1]), .I2(n241_adj_4964), 
            .I3(n44326), .O(n16245[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5303_4 (.CI(n44326), .I0(n16789[1]), .I1(n241_adj_4964), 
            .CO(n44327));
    SB_LUT4 add_5403_3_lut (.I0(GND_net), .I1(n18221[0]), .I2(n177_adj_4962), 
            .I3(n44516), .O(n17884[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5303_3_lut (.I0(GND_net), .I1(n16789[0]), .I2(n168_adj_4960), 
            .I3(n44325), .O(n16245[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n356[5]), .I1(n356[6]), .I2(n13_adj_5169), 
            .I3(GND_net), .O(n10_adj_5251));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_5252));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i22_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter_2283__i0 (.Q(counter[0]), .C(clk16MHz), .D(n34[0]), 
            .R(counter_31__N_3995));   // verilog/motorControl.v(26[16:25])
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_5249), .I1(n356[17]), .I2(n35_adj_5129), 
            .I3(GND_net), .O(n30_adj_5253));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38756_4_lut (.I0(n33_adj_5128), .I1(n31_adj_5134), .I2(n29_adj_5131), 
            .I3(n54553), .O(n54549));
    defparam i38756_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39669_4_lut (.I0(n30_adj_5253), .I1(n10_adj_5251), .I2(n35_adj_5129), 
            .I3(n54547), .O(n55462));   // verilog/motorControl.v(53[12:29])
    defparam i39669_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39057_3_lut (.I0(n55299), .I1(n356[15]), .I2(n31_adj_5134), 
            .I3(GND_net), .O(n54850));   // verilog/motorControl.v(53[12:29])
    defparam i39057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_26_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[10]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_5255));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39753_4_lut (.I0(n54850), .I1(n55462), .I2(n35_adj_5129), 
            .I3(n54549), .O(n55546));   // verilog/motorControl.v(53[12:29])
    defparam i39753_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_5256));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39754_3_lut (.I0(n55546), .I1(n356[18]), .I2(n37_adj_5130), 
            .I3(GND_net), .O(n55547));   // verilog/motorControl.v(53[12:29])
    defparam i39754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_5257));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39507_3_lut (.I0(n6_adj_5258), .I1(n356[10]), .I2(n21_adj_5164), 
            .I3(GND_net), .O(n55300));   // verilog/motorControl.v(53[12:29])
    defparam i39507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39508_3_lut (.I0(n55300), .I1(n356[11]), .I2(n23_adj_5135), 
            .I3(GND_net), .O(n55301));   // verilog/motorControl.v(53[12:29])
    defparam i39508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38740_4_lut (.I0(n43_adj_5144), .I1(n25_adj_5141), .I2(n23_adj_5135), 
            .I3(n54560), .O(n54533));
    defparam i38740_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_5259));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[11]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_5261));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[12]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5416[13]));   // verilog/motorControl.v(57[22:31])
    defparam unary_minus_26_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_5264));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_5185));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_5184));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_5183));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39350_4_lut (.I0(n24_adj_5192), .I1(n8_adj_5191), .I2(n45_adj_5142), 
            .I3(n54531), .O(n55143));   // verilog/motorControl.v(53[12:29])
    defparam i39350_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_17_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_5265));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39055_3_lut (.I0(n55301), .I1(n356[12]), .I2(n25_adj_5141), 
            .I3(GND_net), .O(n54848));   // verilog/motorControl.v(53[12:29])
    defparam i39055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39728_3_lut (.I0(n55547), .I1(n356[19]), .I2(n39_adj_5127), 
            .I3(GND_net), .O(n55521));   // verilog/motorControl.v(53[12:29])
    defparam i39728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_5182));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38742_4_lut (.I0(n43_adj_5144), .I1(n41_adj_5125), .I2(n39_adj_5127), 
            .I3(n55492), .O(n54535));
    defparam i38742_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_5266));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_5180));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39603_4_lut (.I0(n54848), .I1(n55143), .I2(n45_adj_5142), 
            .I3(n54533), .O(n55396));   // verilog/motorControl.v(53[12:29])
    defparam i39603_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39063_3_lut (.I0(n55521), .I1(n356[20]), .I2(n41_adj_5125), 
            .I3(GND_net), .O(n54856));   // verilog/motorControl.v(53[12:29])
    defparam i39063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i4_3_lut (.I0(n54263), .I1(n382[1]), .I2(n356[1]), 
            .I3(GND_net), .O(n4_adj_5268));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39499_3_lut (.I0(n4_adj_5268), .I1(n382[13]), .I2(n356[13]), 
            .I3(GND_net), .O(n55292));   // verilog/motorControl.v(53[33:53])
    defparam i39499_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i39500_3_lut (.I0(n55292), .I1(n382[14]), .I2(n356[14]), .I3(GND_net), 
            .O(n55293));   // verilog/motorControl.v(53[33:53])
    defparam i39500_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_16_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_5179));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_5178));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5303_3 (.CI(n44325), .I0(n16789[0]), .I1(n168_adj_4960), 
            .CO(n44326));
    SB_LUT4 i38710_4_lut (.I0(n356[16]), .I1(n56795), .I2(n382[16]), .I3(n54899), 
            .O(n54503));
    defparam i38710_4_lut.LUT_INIT = 16'h5a7b;
    SB_DFF \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk16MHz), .D(n29289));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 mult_16_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_5177));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39671_4_lut (.I0(n30_adj_5211), .I1(n10_adj_5210), .I2(n56819), 
            .I3(n54501), .O(n55464));   // verilog/motorControl.v(53[33:53])
    defparam i39671_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39067_3_lut (.I0(n55293), .I1(n382[15]), .I2(n356[15]), .I3(GND_net), 
            .O(n54860));   // verilog/motorControl.v(53[33:53])
    defparam i39067_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5478_3 (.CI(n44616), .I0(n19029[0]), .I1(n189), .CO(n44617));
    SB_LUT4 i39755_4_lut (.I0(n54860), .I1(n55464), .I2(n56819), .I3(n54503), 
            .O(n55548));   // verilog/motorControl.v(53[33:53])
    defparam i39755_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_5176));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_5174));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5303_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n16245[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5303_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5403_3 (.CI(n44516), .I0(n18221[0]), .I1(n177_adj_4962), 
            .CO(n44517));
    SB_CARRY add_5303_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n44325));
    SB_LUT4 i39756_3_lut (.I0(n55548), .I1(n382[18]), .I2(n356[18]), .I3(GND_net), 
            .O(n55549));   // verilog/motorControl.v(53[33:53])
    defparam i39756_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY mult_16_add_1225_23 (.CI(n44722), .I0(n11938[20]), .I1(GND_net), 
            .CO(n44723));
    SB_LUT4 i39726_3_lut (.I0(n55549), .I1(n382[19]), .I2(n356[19]), .I3(GND_net), 
            .O(n55519));   // verilog/motorControl.v(53[33:53])
    defparam i39726_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38699_4_lut (.I0(n356[21]), .I1(n56787), .I2(n382[21]), .I3(n55524), 
            .O(n54492));
    defparam i38699_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i45_rep_136_2_lut (.I0(n356[22]), .I1(n382[22]), 
            .I2(GND_net), .I3(GND_net), .O(n56785));   // verilog/motorControl.v(53[33:53])
    defparam LessThan_21_i45_rep_136_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5139_19_lut (.I0(GND_net), .I1(n13789[16]), .I2(GND_net), 
            .I3(n44677), .O(n12908[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5503_9_lut (.I0(GND_net), .I1(n19236[6]), .I2(n630), .I3(n44324), 
            .O(n19109[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5503_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5503_8_lut (.I0(GND_net), .I1(n19236[5]), .I2(n557), .I3(n44323), 
            .O(n19109[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_19 (.CI(n44677), .I0(n13789[16]), .I1(GND_net), 
            .CO(n44678));
    SB_LUT4 add_5403_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n17884[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5403_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5403_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n44516));
    SB_LUT4 add_5139_18_lut (.I0(GND_net), .I1(n13789[15]), .I2(GND_net), 
            .I3(n44676), .O(n12908[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5503_8 (.CI(n44323), .I0(n19236[5]), .I1(n557), .CO(n44324));
    SB_LUT4 i39605_4_lut (.I0(n54858), .I1(n55145), .I2(n56785), .I3(n54490), 
            .O(n55398));   // verilog/motorControl.v(53[33:53])
    defparam i39605_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_5167));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39073_3_lut (.I0(n55519), .I1(n382[20]), .I2(n356[20]), .I3(GND_net), 
            .O(n54866));   // verilog/motorControl.v(53[33:53])
    defparam i39073_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_16_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_5166));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5503_7_lut (.I0(GND_net), .I1(n19236[4]), .I2(n484_adj_4910), 
            .I3(n44322), .O(n19109[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5503_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i8_3_lut (.I0(n130[7]), .I1(n182[7]), .I2(n181), .I3(GND_net), 
            .O(n207[7]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39695_4_lut (.I0(n54866), .I1(n55398), .I2(n56785), .I3(n54492), 
            .O(n55488));   // verilog/motorControl.v(53[33:53])
    defparam i39695_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_15_i8_3_lut (.I0(n207[7]), .I1(IntegralLimit[7]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [7]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39693_4_lut (.I0(n54856), .I1(n55396), .I2(n45_adj_5142), 
            .I3(n54535), .O(n55486));   // verilog/motorControl.v(53[12:29])
    defparam i39693_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(n55488), .I1(control_update), .I2(n356[23]), 
            .I3(n47_adj_5269), .O(n52036));
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'h0c44;
    SB_LUT4 i1_4_lut_adj_1712 (.I0(n52036), .I1(n55486), .I2(deadband[23]), 
            .I3(n356[23]), .O(n29234));
    defparam i1_4_lut_adj_1712.LUT_INIT = 16'h2a02;
    SB_LUT4 add_5478_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n18849[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5478_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5503_7 (.CI(n44322), .I0(n19236[4]), .I1(n484_adj_4910), 
            .CO(n44323));
    SB_LUT4 mult_17_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_5162));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5161));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_22_lut (.I0(GND_net), .I1(n11938[19]), .I2(GND_net), 
            .I3(n44721), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_5158));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i151_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_22 (.CI(n44721), .I0(n11938[19]), .I1(GND_net), 
            .CO(n44722));
    SB_LUT4 mult_17_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_5151));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5459_11_lut (.I0(GND_net), .I1(n18849[8]), .I2(n770_adj_4907), 
            .I3(n43477), .O(n18629[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_5150));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_5148));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_5147));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5459_10_lut (.I0(GND_net), .I1(n18849[7]), .I2(n697), 
            .I3(n43476), .O(n18629[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_5146));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i200_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5459_10 (.CI(n43476), .I0(n18849[7]), .I1(n697), .CO(n43477));
    SB_LUT4 mult_17_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_5145));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5459_9_lut (.I0(GND_net), .I1(n18849[6]), .I2(n624), .I3(n43475), 
            .O(n18629[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_9 (.CI(n43475), .I0(n18849[6]), .I1(n624), .CO(n43476));
    SB_LUT4 mult_16_add_1225_21_lut (.I0(GND_net), .I1(n11938[18]), .I2(GND_net), 
            .I3(n44720), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5459_8_lut (.I0(GND_net), .I1(n18849[5]), .I2(n551), .I3(n43474), 
            .O(n18629[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_18 (.CI(n44676), .I0(n13789[15]), .I1(GND_net), 
            .CO(n44677));
    SB_CARRY add_5478_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n44616));
    SB_LUT4 add_5253_19_lut (.I0(GND_net), .I1(n15956[16]), .I2(GND_net), 
            .I3(n44615), .O(n15309[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5503_6_lut (.I0(GND_net), .I1(n19236[3]), .I2(n411_adj_4892), 
            .I3(n44321), .O(n19109[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5503_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5523_7_lut (.I0(GND_net), .I1(n51035), .I2(n490), .I3(n44515), 
            .O(n19285[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5523_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5503_6 (.CI(n44321), .I0(n19236[3]), .I1(n411_adj_4892), 
            .CO(n44322));
    SB_LUT4 add_5253_18_lut (.I0(GND_net), .I1(n15956[15]), .I2(GND_net), 
            .I3(n44614), .O(n15309[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5523_6_lut (.I0(GND_net), .I1(n19369[3]), .I2(n417_adj_5270), 
            .I3(n44514), .O(n19285[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5523_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5503_5_lut (.I0(GND_net), .I1(n19236[2]), .I2(n338_adj_5271), 
            .I3(n44320), .O(n19109[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5503_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5503_5 (.CI(n44320), .I0(n19236[2]), .I1(n338_adj_5271), 
            .CO(n44321));
    SB_LUT4 add_5503_4_lut (.I0(GND_net), .I1(n19236[1]), .I2(n265_adj_5272), 
            .I3(n44319), .O(n19109[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_8 (.CI(n43474), .I0(n18849[5]), .I1(n551), .CO(n43475));
    SB_LUT4 add_5459_7_lut (.I0(GND_net), .I1(n18849[4]), .I2(n478_adj_5273), 
            .I3(n43473), .O(n18629[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_17_lut (.I0(GND_net), .I1(n13789[14]), .I2(GND_net), 
            .I3(n44675), .O(n12908[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_7 (.CI(n43473), .I0(n18849[4]), .I1(n478_adj_5273), 
            .CO(n43474));
    SB_CARRY add_5503_4 (.CI(n44319), .I0(n19236[1]), .I1(n265_adj_5272), 
            .CO(n44320));
    SB_CARRY mult_16_add_1225_21 (.CI(n44720), .I0(n11938[18]), .I1(GND_net), 
            .CO(n44721));
    SB_LUT4 add_5459_6_lut (.I0(GND_net), .I1(n18849[3]), .I2(n405_adj_5274), 
            .I3(n43472), .O(n18629[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_6 (.CI(n43472), .I0(n18849[3]), .I1(n405_adj_5274), 
            .CO(n43473));
    SB_LUT4 mult_17_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_5126));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_5123));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5459_5_lut (.I0(GND_net), .I1(n18849[2]), .I2(n332_adj_5275), 
            .I3(n43471), .O(n18629[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_5 (.CI(n43471), .I0(n18849[2]), .I1(n332_adj_5275), 
            .CO(n43472));
    SB_LUT4 mult_16_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_5122));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_5121));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_5120));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i357_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5523_6 (.CI(n44514), .I0(n19369[3]), .I1(n417_adj_5270), 
            .CO(n44515));
    SB_LUT4 add_5503_3_lut (.I0(GND_net), .I1(n19236[0]), .I2(n192_adj_5276), 
            .I3(n44318), .O(n19109[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5503_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5523_5_lut (.I0(GND_net), .I1(n19369[2]), .I2(n344_adj_5277), 
            .I3(n44513), .O(n19285[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5523_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5503_3 (.CI(n44318), .I0(n19236[0]), .I1(n192_adj_5276), 
            .CO(n44319));
    SB_LUT4 add_5459_4_lut (.I0(GND_net), .I1(n18849[1]), .I2(n259_adj_5278), 
            .I3(n43470), .O(n18629[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_4 (.CI(n43470), .I0(n18849[1]), .I1(n259_adj_5278), 
            .CO(n43471));
    SB_LUT4 mult_17_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_5119));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_5118));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5459_3_lut (.I0(GND_net), .I1(n18849[0]), .I2(n186_adj_5279), 
            .I3(n43469), .O(n18629[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_3 (.CI(n43469), .I0(n18849[0]), .I1(n186_adj_5279), 
            .CO(n43470));
    SB_LUT4 add_5459_2_lut (.I0(GND_net), .I1(n44_adj_5280), .I2(n113_adj_5281), 
            .I3(GND_net), .O(n18629[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5523_5 (.CI(n44513), .I0(n19369[2]), .I1(n344_adj_5277), 
            .CO(n44514));
    SB_LUT4 mult_17_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_5117));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5253_18 (.CI(n44614), .I0(n15956[15]), .I1(GND_net), 
            .CO(n44615));
    SB_LUT4 add_5503_2_lut (.I0(GND_net), .I1(n50_adj_5282), .I2(n119_adj_5283), 
            .I3(GND_net), .O(n19109[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_2 (.CI(GND_net), .I0(n44_adj_5280), .I1(n113_adj_5281), 
            .CO(n43469));
    SB_LUT4 mult_16_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i15_3_lut (.I0(n130[14]), .I1(n182[14]), .I2(n181), 
            .I3(GND_net), .O(n207[14]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5503_2 (.CI(GND_net), .I0(n50_adj_5282), .I1(n119_adj_5283), 
            .CO(n44318));
    SB_LUT4 add_5523_4_lut (.I0(GND_net), .I1(n19369[1]), .I2(n271_adj_5285), 
            .I3(n44512), .O(n19285[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5523_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5523_4 (.CI(n44512), .I0(n19369[1]), .I1(n271_adj_5285), 
            .CO(n44513));
    SB_LUT4 add_5334_16_lut (.I0(GND_net), .I1(n17269[13]), .I2(n1120_adj_5286), 
            .I3(n44317), .O(n16789[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i15_3_lut (.I0(n207[14]), .I1(IntegralLimit[14]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [14]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_5116));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5334_15_lut (.I0(GND_net), .I1(n17269[12]), .I2(n1047_adj_5287), 
            .I3(n44316), .O(n16789[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_20_lut (.I0(GND_net), .I1(n11938[17]), .I2(GND_net), 
            .I3(n44719), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_17_lut (.I0(GND_net), .I1(n15956[14]), .I2(GND_net), 
            .I3(n44613), .O(n15309[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i504_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5334_15 (.CI(n44316), .I0(n17269[12]), .I1(n1047_adj_5287), 
            .CO(n44317));
    SB_LUT4 add_5523_3_lut (.I0(GND_net), .I1(n19369[0]), .I2(n198_adj_5288), 
            .I3(n44511), .O(n19285[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5523_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_5115));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5114));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5334_14_lut (.I0(GND_net), .I1(n17269[11]), .I2(n974_adj_5289), 
            .I3(n44315), .O(n16789[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_5113));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i249_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5253_17 (.CI(n44613), .I0(n15956[14]), .I1(GND_net), 
            .CO(n44614));
    SB_CARRY add_5523_3 (.CI(n44511), .I0(n19369[0]), .I1(n198_adj_5288), 
            .CO(n44512));
    SB_LUT4 mult_17_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5523_2_lut (.I0(GND_net), .I1(n56_adj_5290), .I2(n125_adj_5291), 
            .I3(GND_net), .O(n19285[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5523_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_17 (.CI(n44675), .I0(n13789[14]), .I1(GND_net), 
            .CO(n44676));
    SB_LUT4 add_5253_16_lut (.I0(GND_net), .I1(n15956[13]), .I2(n1111_adj_5292), 
            .I3(n44612), .O(n15309[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_20 (.CI(n44719), .I0(n11938[17]), .I1(GND_net), 
            .CO(n44720));
    SB_LUT4 add_5139_16_lut (.I0(GND_net), .I1(n13789[13]), .I2(n1102_adj_5293), 
            .I3(n44674), .O(n12908[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_19_lut (.I0(GND_net), .I1(n11938[16]), .I2(GND_net), 
            .I3(n44718), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5334_14 (.CI(n44315), .I0(n17269[11]), .I1(n974_adj_5289), 
            .CO(n44316));
    SB_CARRY add_5253_16 (.CI(n44612), .I0(n15956[13]), .I1(n1111_adj_5292), 
            .CO(n44613));
    SB_CARRY add_5139_16 (.CI(n44674), .I0(n13789[13]), .I1(n1102_adj_5293), 
            .CO(n44675));
    SB_CARRY mult_16_add_1225_19 (.CI(n44718), .I0(n11938[16]), .I1(GND_net), 
            .CO(n44719));
    SB_LUT4 mult_16_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i167_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5523_2 (.CI(GND_net), .I0(n56_adj_5290), .I1(n125_adj_5291), 
            .CO(n44511));
    SB_LUT4 add_5427_13_lut (.I0(GND_net), .I1(n18508[10]), .I2(n910_adj_5294), 
            .I3(n44510), .O(n18221[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_18_lut (.I0(GND_net), .I1(n11938[15]), .I2(GND_net), 
            .I3(n44717), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_15_lut (.I0(GND_net), .I1(n15956[12]), .I2(n1038_adj_5295), 
            .I3(n44611), .O(n15309[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5427_12_lut (.I0(GND_net), .I1(n18508[9]), .I2(n837_adj_5296), 
            .I3(n44509), .O(n18221[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_15 (.CI(n44611), .I0(n15956[12]), .I1(n1038_adj_5295), 
            .CO(n44612));
    SB_LUT4 add_5334_13_lut (.I0(GND_net), .I1(n17269[10]), .I2(n901_adj_5297), 
            .I3(n44314), .O(n16789[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_5106));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5253_14_lut (.I0(GND_net), .I1(n15956[11]), .I2(n965_adj_5298), 
            .I3(n44610), .O(n15309[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_15_lut (.I0(GND_net), .I1(n13789[12]), .I2(n1029_adj_5299), 
            .I3(n44673), .O(n12908[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_15 (.CI(n44673), .I0(n13789[12]), .I1(n1029_adj_5299), 
            .CO(n44674));
    SB_CARRY add_5253_14 (.CI(n44610), .I0(n15956[11]), .I1(n965_adj_5298), 
            .CO(n44611));
    SB_CARRY add_5427_12 (.CI(n44509), .I0(n18508[9]), .I1(n837_adj_5296), 
            .CO(n44510));
    SB_CARRY add_5334_13 (.CI(n44314), .I0(n17269[10]), .I1(n901_adj_5297), 
            .CO(n44315));
    SB_LUT4 add_5427_11_lut (.I0(GND_net), .I1(n18508[8]), .I2(n764_adj_5300), 
            .I3(n44508), .O(n18221[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5334_12_lut (.I0(GND_net), .I1(n17269[9]), .I2(n828_adj_5301), 
            .I3(n44313), .O(n16789[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5334_12 (.CI(n44313), .I0(n17269[9]), .I1(n828_adj_5301), 
            .CO(n44314));
    SB_LUT4 add_5139_14_lut (.I0(GND_net), .I1(n13789[11]), .I2(n956_adj_5302), 
            .I3(n44672), .O(n12908[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5334_11_lut (.I0(GND_net), .I1(n17269[8]), .I2(n755_adj_5303), 
            .I3(n44312), .O(n16789[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5334_11 (.CI(n44312), .I0(n17269[8]), .I1(n755_adj_5303), 
            .CO(n44313));
    SB_LUT4 add_5334_10_lut (.I0(GND_net), .I1(n17269[7]), .I2(n682_adj_5304), 
            .I3(n44311), .O(n16789[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(n29234), .I1(control_update), .I2(GND_net), 
            .I3(GND_net), .O(n28830));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14867_3_lut (.I0(n356[1]), .I1(n436[1]), .I2(n10863), .I3(GND_net), 
            .O(n28938));   // verilog/motorControl.v(43[14] 63[8])
    defparam i14867_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5427_11 (.CI(n44508), .I0(n18508[8]), .I1(n764_adj_5300), 
            .CO(n44509));
    SB_CARRY add_5334_10 (.CI(n44311), .I0(n17269[7]), .I1(n682_adj_5304), 
            .CO(n44312));
    SB_CARRY mult_16_add_1225_18 (.CI(n44717), .I0(n11938[15]), .I1(GND_net), 
            .CO(n44718));
    SB_LUT4 mult_16_add_1225_17_lut (.I0(GND_net), .I1(n11938[14]), .I2(GND_net), 
            .I3(n44716), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_17 (.CI(n44716), .I0(n11938[14]), .I1(GND_net), 
            .CO(n44717));
    SB_CARRY add_5139_14 (.CI(n44672), .I0(n13789[11]), .I1(n956_adj_5302), 
            .CO(n44673));
    SB_LUT4 mult_17_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_5105));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5427_10_lut (.I0(GND_net), .I1(n18508[7]), .I2(n691_adj_5305), 
            .I3(n44507), .O(n18221[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i1_3_lut (.I0(n130[0]), .I1(n182[0]), .I2(n181), .I3(GND_net), 
            .O(n207[0]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i1_3_lut (.I0(n207[0]), .I1(IntegralLimit[0]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [0]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n306[0]));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n257[0]));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_5103));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_5101));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_5100));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_16_lut (.I0(GND_net), .I1(n11938[13]), .I2(n1096_adj_5306), 
            .I3(n44715), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_13_lut (.I0(GND_net), .I1(n13789[10]), .I2(n883_adj_5307), 
            .I3(n44671), .O(n12908[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_13_lut (.I0(GND_net), .I1(n15956[10]), .I2(n892_adj_5308), 
            .I3(n44609), .O(n15309[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5427_10 (.CI(n44507), .I0(n18508[7]), .I1(n691_adj_5305), 
            .CO(n44508));
    SB_LUT4 add_5334_9_lut (.I0(GND_net), .I1(n17269[6]), .I2(n609_adj_5309), 
            .I3(n44310), .O(n16789[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5334_9 (.CI(n44310), .I0(n17269[6]), .I1(n609_adj_5309), 
            .CO(n44311));
    SB_CARRY add_5253_13 (.CI(n44609), .I0(n15956[10]), .I1(n892_adj_5308), 
            .CO(n44610));
    SB_LUT4 add_5427_9_lut (.I0(GND_net), .I1(n18508[6]), .I2(n618_adj_5310), 
            .I3(n44506), .O(n18221[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5334_8_lut (.I0(GND_net), .I1(n17269[5]), .I2(n536_adj_5311), 
            .I3(n44309), .O(n16789[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5334_8 (.CI(n44309), .I0(n17269[5]), .I1(n536_adj_5311), 
            .CO(n44310));
    SB_LUT4 mult_16_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_5099));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5253_12_lut (.I0(GND_net), .I1(n15956[9]), .I2(n819_adj_5312), 
            .I3(n44608), .O(n15309[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_12 (.CI(n44608), .I0(n15956[9]), .I1(n819_adj_5312), 
            .CO(n44609));
    SB_CARRY add_5427_9 (.CI(n44506), .I0(n18508[6]), .I1(n618_adj_5310), 
            .CO(n44507));
    SB_LUT4 add_5334_7_lut (.I0(GND_net), .I1(n17269[4]), .I2(n463_adj_5313), 
            .I3(n44308), .O(n16789[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5427_8_lut (.I0(GND_net), .I1(n18508[5]), .I2(n545_adj_5314), 
            .I3(n44505), .O(n18221[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_5098));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5334_7 (.CI(n44308), .I0(n17269[4]), .I1(n463_adj_5313), 
            .CO(n44309));
    SB_CARRY add_5427_8 (.CI(n44505), .I0(n18508[5]), .I1(n545_adj_5314), 
            .CO(n44506));
    SB_LUT4 add_5334_6_lut (.I0(GND_net), .I1(n17269[3]), .I2(n390_adj_5315), 
            .I3(n44307), .O(n16789[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5334_6 (.CI(n44307), .I0(n17269[3]), .I1(n390_adj_5315), 
            .CO(n44308));
    SB_LUT4 add_5334_5_lut (.I0(GND_net), .I1(n17269[2]), .I2(n317_adj_5316), 
            .I3(n44306), .O(n16789[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5427_7_lut (.I0(GND_net), .I1(n18508[4]), .I2(n472_adj_5317), 
            .I3(n44504), .O(n18221[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5334_5 (.CI(n44306), .I0(n17269[2]), .I1(n317_adj_5316), 
            .CO(n44307));
    SB_LUT4 add_5334_4_lut (.I0(GND_net), .I1(n17269[1]), .I2(n244_adj_5318), 
            .I3(n44305), .O(n16789[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5427_7 (.CI(n44504), .I0(n18508[4]), .I1(n472_adj_5317), 
            .CO(n44505));
    SB_CARRY add_5334_4 (.CI(n44305), .I0(n17269[1]), .I1(n244_adj_5318), 
            .CO(n44306));
    SB_LUT4 add_5334_3_lut (.I0(GND_net), .I1(n17269[0]), .I2(n171_adj_5319), 
            .I3(n44304), .O(n16789[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_13 (.CI(n44671), .I0(n13789[10]), .I1(n883_adj_5307), 
            .CO(n44672));
    SB_LUT4 add_5253_11_lut (.I0(GND_net), .I1(n15956[8]), .I2(n746_adj_5320), 
            .I3(n44607), .O(n15309[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_12_lut (.I0(GND_net), .I1(n13789[9]), .I2(n810_adj_5321), 
            .I3(n44670), .O(n12908[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_12 (.CI(n44670), .I0(n13789[9]), .I1(n810_adj_5321), 
            .CO(n44671));
    SB_CARRY add_5253_11 (.CI(n44607), .I0(n15956[8]), .I1(n746_adj_5320), 
            .CO(n44608));
    SB_LUT4 add_5427_6_lut (.I0(GND_net), .I1(n18508[3]), .I2(n399_adj_5322), 
            .I3(n44503), .O(n18221[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5334_3 (.CI(n44304), .I0(n17269[0]), .I1(n171_adj_5319), 
            .CO(n44305));
    SB_LUT4 add_5334_2_lut (.I0(GND_net), .I1(n29_adj_5323), .I2(n98_adj_5324), 
            .I3(GND_net), .O(n16789[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5334_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5334_2 (.CI(GND_net), .I0(n29_adj_5323), .I1(n98_adj_5324), 
            .CO(n44304));
    SB_CARRY mult_16_add_1225_16 (.CI(n44715), .I0(n11938[13]), .I1(n1096_adj_5306), 
            .CO(n44716));
    SB_CARRY add_5427_6 (.CI(n44503), .I0(n18508[3]), .I1(n399_adj_5322), 
            .CO(n44504));
    SB_LUT4 add_5363_15_lut (.I0(GND_net), .I1(n17689[12]), .I2(n1050_adj_5325), 
            .I3(n44303), .O(n17269[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5427_5_lut (.I0(GND_net), .I1(n18508[2]), .I2(n326_adj_5326), 
            .I3(n44502), .O(n18221[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5363_14_lut (.I0(GND_net), .I1(n17689[11]), .I2(n977_adj_5327), 
            .I3(n44302), .O(n17269[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_14 (.CI(n44302), .I0(n17689[11]), .I1(n977_adj_5327), 
            .CO(n44303));
    SB_CARRY add_5427_5 (.CI(n44502), .I0(n18508[2]), .I1(n326_adj_5326), 
            .CO(n44503));
    SB_LUT4 add_5139_11_lut (.I0(GND_net), .I1(n13789[8]), .I2(n737_adj_5328), 
            .I3(n44669), .O(n12908[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_10_lut (.I0(GND_net), .I1(n15956[7]), .I2(n673_adj_5329), 
            .I3(n44606), .O(n15309[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5363_13_lut (.I0(GND_net), .I1(n17689[10]), .I2(n904_adj_5330), 
            .I3(n44301), .O(n17269[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_13 (.CI(n44301), .I0(n17689[10]), .I1(n904_adj_5330), 
            .CO(n44302));
    SB_LUT4 add_5363_12_lut (.I0(GND_net), .I1(n17689[9]), .I2(n831_adj_5331), 
            .I3(n44300), .O(n17269[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_10 (.CI(n44606), .I0(n15956[7]), .I1(n673_adj_5329), 
            .CO(n44607));
    SB_LUT4 add_5427_4_lut (.I0(GND_net), .I1(n18508[1]), .I2(n253_adj_5332), 
            .I3(n44501), .O(n18221[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5427_4 (.CI(n44501), .I0(n18508[1]), .I1(n253_adj_5332), 
            .CO(n44502));
    SB_LUT4 add_5427_3_lut (.I0(GND_net), .I1(n18508[0]), .I2(n180_adj_5333), 
            .I3(n44500), .O(n18221[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_12 (.CI(n44300), .I0(n17689[9]), .I1(n831_adj_5331), 
            .CO(n44301));
    SB_LUT4 add_5363_11_lut (.I0(GND_net), .I1(n17689[8]), .I2(n758_adj_5334), 
            .I3(n44299), .O(n17269[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_11 (.CI(n44299), .I0(n17689[8]), .I1(n758_adj_5334), 
            .CO(n44300));
    SB_CARRY add_5427_3 (.CI(n44500), .I0(n18508[0]), .I1(n180_adj_5333), 
            .CO(n44501));
    SB_LUT4 add_5363_10_lut (.I0(GND_net), .I1(n17689[7]), .I2(n685_adj_5335), 
            .I3(n44298), .O(n17269[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_15_lut (.I0(GND_net), .I1(n11938[12]), .I2(n1023_adj_5336), 
            .I3(n44714), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_11 (.CI(n44669), .I0(n13789[8]), .I1(n737_adj_5328), 
            .CO(n44670));
    SB_CARRY add_5363_10 (.CI(n44298), .I0(n17689[7]), .I1(n685_adj_5335), 
            .CO(n44299));
    SB_LUT4 add_5253_9_lut (.I0(GND_net), .I1(n15956[6]), .I2(n600_adj_5337), 
            .I3(n44605), .O(n15309[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5427_2_lut (.I0(GND_net), .I1(n38_adj_5338), .I2(n107_adj_5339), 
            .I3(GND_net), .O(n18221[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5363_9_lut (.I0(GND_net), .I1(n17689[6]), .I2(n612_adj_5340), 
            .I3(n44297), .O(n17269[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_9 (.CI(n44297), .I0(n17689[6]), .I1(n612_adj_5340), 
            .CO(n44298));
    SB_CARRY add_5427_2 (.CI(GND_net), .I0(n38_adj_5338), .I1(n107_adj_5339), 
            .CO(n44500));
    SB_LUT4 add_5363_8_lut (.I0(GND_net), .I1(n17689[5]), .I2(n539_adj_5341), 
            .I3(n44296), .O(n17269[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_8 (.CI(n44296), .I0(n17689[5]), .I1(n539_adj_5341), 
            .CO(n44297));
    SB_CARRY mult_16_add_1225_15 (.CI(n44714), .I0(n11938[12]), .I1(n1023_adj_5336), 
            .CO(n44715));
    SB_LUT4 add_5139_10_lut (.I0(GND_net), .I1(n13789[7]), .I2(n664_adj_5342), 
            .I3(n44668), .O(n12908[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_9 (.CI(n44605), .I0(n15956[6]), .I1(n600_adj_5337), 
            .CO(n44606));
    SB_LUT4 add_5449_12_lut (.I0(GND_net), .I1(n18749[9]), .I2(n840_adj_5343), 
            .I3(n44499), .O(n18508[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5363_7_lut (.I0(GND_net), .I1(n17689[4]), .I2(n466_adj_5344), 
            .I3(n44295), .O(n17269[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_7 (.CI(n44295), .I0(n17689[4]), .I1(n466_adj_5344), 
            .CO(n44296));
    SB_LUT4 add_5449_11_lut (.I0(GND_net), .I1(n18749[8]), .I2(n767_adj_5345), 
            .I3(n44498), .O(n18508[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5363_6_lut (.I0(GND_net), .I1(n17689[3]), .I2(n393_adj_5346), 
            .I3(n44294), .O(n17269[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_8_lut (.I0(GND_net), .I1(n15956[5]), .I2(n527_adj_5347), 
            .I3(n44604), .O(n15309[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_8 (.CI(n44604), .I0(n15956[5]), .I1(n527_adj_5347), 
            .CO(n44605));
    SB_CARRY add_5449_11 (.CI(n44498), .I0(n18749[8]), .I1(n767_adj_5345), 
            .CO(n44499));
    SB_CARRY add_5363_6 (.CI(n44294), .I0(n17689[3]), .I1(n393_adj_5346), 
            .CO(n44295));
    SB_LUT4 add_5449_10_lut (.I0(GND_net), .I1(n18749[7]), .I2(n694_adj_5266), 
            .I3(n44497), .O(n18508[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5363_5_lut (.I0(GND_net), .I1(n17689[2]), .I2(n320_adj_5265), 
            .I3(n44293), .O(n17269[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_7_lut (.I0(GND_net), .I1(n15956[4]), .I2(n454_adj_5264), 
            .I3(n44603), .O(n15309[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5449_10 (.CI(n44497), .I0(n18749[7]), .I1(n694_adj_5266), 
            .CO(n44498));
    SB_CARRY add_5363_5 (.CI(n44293), .I0(n17689[2]), .I1(n320_adj_5265), 
            .CO(n44294));
    SB_LUT4 add_5363_4_lut (.I0(GND_net), .I1(n17689[1]), .I2(n247_adj_5259), 
            .I3(n44292), .O(n17269[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_4 (.CI(n44292), .I0(n17689[1]), .I1(n247_adj_5259), 
            .CO(n44293));
    SB_LUT4 add_5363_3_lut (.I0(GND_net), .I1(n17689[0]), .I2(n174_adj_5256), 
            .I3(n44291), .O(n17269[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5449_9_lut (.I0(GND_net), .I1(n18749[6]), .I2(n621_adj_5255), 
            .I3(n44496), .O(n18508[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_3 (.CI(n44291), .I0(n17689[0]), .I1(n174_adj_5256), 
            .CO(n44292));
    SB_LUT4 add_5363_2_lut (.I0(GND_net), .I1(n32_adj_5252), .I2(n101_adj_5247), 
            .I3(GND_net), .O(n17269[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5363_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5363_2 (.CI(GND_net), .I0(n32_adj_5252), .I1(n101_adj_5247), 
            .CO(n44291));
    SB_CARRY add_5253_7 (.CI(n44603), .I0(n15956[4]), .I1(n454_adj_5264), 
            .CO(n44604));
    SB_CARRY add_5449_9 (.CI(n44496), .I0(n18749[6]), .I1(n621_adj_5255), 
            .CO(n44497));
    SB_LUT4 add_5517_8_lut (.I0(GND_net), .I1(n19333[5]), .I2(n560_adj_5246), 
            .I3(n44290), .O(n19236[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5517_7_lut (.I0(GND_net), .I1(n19333[4]), .I2(n487_adj_5245), 
            .I3(n44289), .O(n19236[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5449_8_lut (.I0(GND_net), .I1(n18749[5]), .I2(n548_adj_5244), 
            .I3(n44495), .O(n18508[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5517_7 (.CI(n44289), .I0(n19333[4]), .I1(n487_adj_5245), 
            .CO(n44290));
    SB_LUT4 add_5517_6_lut (.I0(GND_net), .I1(n19333[3]), .I2(n414_adj_5243), 
            .I3(n44288), .O(n19236[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5449_8 (.CI(n44495), .I0(n18749[5]), .I1(n548_adj_5244), 
            .CO(n44496));
    SB_CARRY add_5517_6 (.CI(n44288), .I0(n19333[3]), .I1(n414_adj_5243), 
            .CO(n44289));
    SB_LUT4 add_5517_5_lut (.I0(GND_net), .I1(n19333[2]), .I2(n341_adj_5242), 
            .I3(n44287), .O(n19236[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_10 (.CI(n44668), .I0(n13789[7]), .I1(n664_adj_5342), 
            .CO(n44669));
    SB_LUT4 add_5253_6_lut (.I0(GND_net), .I1(n15956[3]), .I2(n381_adj_5233), 
            .I3(n44602), .O(n15309[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5449_7_lut (.I0(GND_net), .I1(n18749[4]), .I2(n475_adj_5227), 
            .I3(n44494), .O(n18508[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5517_5 (.CI(n44287), .I0(n19333[2]), .I1(n341_adj_5242), 
            .CO(n44288));
    SB_LUT4 add_5517_4_lut (.I0(GND_net), .I1(n19333[1]), .I2(n268_adj_5223), 
            .I3(n44286), .O(n19236[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_9_lut (.I0(GND_net), .I1(n13789[6]), .I2(n591_adj_5222), 
            .I3(n44667), .O(n12908[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_6 (.CI(n44602), .I0(n15956[3]), .I1(n381_adj_5233), 
            .CO(n44603));
    SB_CARRY add_5449_7 (.CI(n44494), .I0(n18749[4]), .I1(n475_adj_5227), 
            .CO(n44495));
    SB_CARRY add_5517_4 (.CI(n44286), .I0(n19333[1]), .I1(n268_adj_5223), 
            .CO(n44287));
    SB_LUT4 add_5449_6_lut (.I0(GND_net), .I1(n18749[3]), .I2(n402_adj_5200), 
            .I3(n44493), .O(n18508[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5517_3_lut (.I0(GND_net), .I1(n19333[0]), .I2(n195_adj_5198), 
            .I3(n44285), .O(n19236[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5517_3 (.CI(n44285), .I0(n19333[0]), .I1(n195_adj_5198), 
            .CO(n44286));
    SB_LUT4 i28838_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [18]), .I3(\Ki[1] ), 
            .O(n19369[0]));   // verilog/motorControl.v(52[27:38])
    defparam i28838_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_5253_5_lut (.I0(GND_net), .I1(n15956[2]), .I2(n308), .I3(n44601), 
            .O(n15309[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5449_6 (.CI(n44493), .I0(n18749[3]), .I1(n402_adj_5200), 
            .CO(n44494));
    SB_LUT4 add_5517_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_4981), 
            .I3(GND_net), .O(n19236[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5517_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_4981), .CO(n44285));
    SB_LUT4 add_5390_14_lut (.I0(GND_net), .I1(n18053[11]), .I2(n980), 
            .I3(n44284), .O(n17689[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5390_13_lut (.I0(GND_net), .I1(n18053[10]), .I2(n907), 
            .I3(n44283), .O(n17689[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5390_13 (.CI(n44283), .I0(n18053[10]), .I1(n907), .CO(n44284));
    SB_LUT4 add_5449_5_lut (.I0(GND_net), .I1(n18749[2]), .I2(n329), .I3(n44492), 
            .O(n18508[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5390_12_lut (.I0(GND_net), .I1(n18053[9]), .I2(n834), 
            .I3(n44282), .O(n17689[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5390_12 (.CI(n44282), .I0(n18053[9]), .I1(n834), .CO(n44283));
    SB_LUT4 add_5390_11_lut (.I0(GND_net), .I1(n18053[8]), .I2(n761), 
            .I3(n44281), .O(n17689[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5390_11 (.CI(n44281), .I0(n18053[8]), .I1(n761), .CO(n44282));
    SB_CARRY add_5449_5 (.CI(n44492), .I0(n18749[2]), .I1(n329), .CO(n44493));
    SB_LUT4 add_5390_10_lut (.I0(GND_net), .I1(n18053[7]), .I2(n688), 
            .I3(n44280), .O(n17689[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28840_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [18]), .I3(\Ki[1] ), 
            .O(n42908));   // verilog/motorControl.v(52[27:38])
    defparam i28840_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_5390_10 (.CI(n44280), .I0(n18053[7]), .I1(n688), .CO(n44281));
    SB_LUT4 add_5449_4_lut (.I0(GND_net), .I1(n18749[1]), .I2(n256), .I3(n44491), 
            .O(n18508[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_5 (.CI(n44601), .I0(n15956[2]), .I1(n308), .CO(n44602));
    SB_LUT4 add_5390_9_lut (.I0(GND_net), .I1(n18053[6]), .I2(n615), .I3(n44279), 
            .O(n17689[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5449_4 (.CI(n44491), .I0(n18749[1]), .I1(n256), .CO(n44492));
    SB_CARRY add_5390_9 (.CI(n44279), .I0(n18053[6]), .I1(n615), .CO(n44280));
    SB_LUT4 add_5390_8_lut (.I0(GND_net), .I1(n18053[5]), .I2(n542), .I3(n44278), 
            .O(n17689[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5390_8 (.CI(n44278), .I0(n18053[5]), .I1(n542), .CO(n44279));
    SB_LUT4 mult_16_add_1225_14_lut (.I0(GND_net), .I1(n11938[11]), .I2(n950), 
            .I3(n44713), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5449_3_lut (.I0(GND_net), .I1(n18749[0]), .I2(n183_adj_4939), 
            .I3(n44490), .O(n18508[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_4_lut (.I0(GND_net), .I1(n15956[1]), .I2(n235), .I3(n44600), 
            .O(n15309[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_9 (.CI(n44667), .I0(n13789[6]), .I1(n591_adj_5222), 
            .CO(n44668));
    SB_LUT4 add_5390_7_lut (.I0(GND_net), .I1(n18053[4]), .I2(n469), .I3(n44277), 
            .O(n17689[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5449_3 (.CI(n44490), .I0(n18749[0]), .I1(n183_adj_4939), 
            .CO(n44491));
    SB_CARRY add_5390_7 (.CI(n44277), .I0(n18053[4]), .I1(n469), .CO(n44278));
    SB_LUT4 add_5390_6_lut (.I0(GND_net), .I1(n18053[3]), .I2(n396), .I3(n44276), 
            .O(n17689[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5449_2_lut (.I0(GND_net), .I1(n41), .I2(n110_adj_4938), 
            .I3(GND_net), .O(n18508[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5449_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_4 (.CI(n44600), .I0(n15956[1]), .I1(n235), .CO(n44601));
    SB_CARRY add_5449_2 (.CI(GND_net), .I0(n41), .I1(n110_adj_4938), .CO(n44490));
    SB_LUT4 mult_17_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3996 [23]), 
            .I1(n11407[21]), .I2(GND_net), .I3(n44489), .O(n10900[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5390_6 (.CI(n44276), .I0(n18053[3]), .I1(n396), .CO(n44277));
    SB_LUT4 add_5390_5_lut (.I0(GND_net), .I1(n18053[2]), .I2(n323), .I3(n44275), 
            .O(n17689[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5390_5 (.CI(n44275), .I0(n18053[2]), .I1(n323), .CO(n44276));
    SB_LUT4 add_5253_3_lut (.I0(GND_net), .I1(n15956[0]), .I2(n162), .I3(n44599), 
            .O(n15309[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5390_4_lut (.I0(GND_net), .I1(n18053[1]), .I2(n250), .I3(n44274), 
            .O(n17689[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_23_lut (.I0(GND_net), .I1(n11407[20]), .I2(GND_net), 
            .I3(n44488), .O(n306[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5390_4 (.CI(n44274), .I0(n18053[1]), .I1(n250), .CO(n44275));
    SB_LUT4 add_5390_3_lut (.I0(GND_net), .I1(n18053[0]), .I2(n177), .I3(n44273), 
            .O(n17689[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_23 (.CI(n44488), .I0(n11407[20]), .I1(GND_net), 
            .CO(n44489));
    SB_CARRY add_5390_3 (.CI(n44273), .I0(n18053[0]), .I1(n177), .CO(n44274));
    SB_LUT4 add_5390_2_lut (.I0(GND_net), .I1(n35_adj_4932), .I2(n104_adj_4931), 
            .I3(GND_net), .O(n17689[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5390_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_22_lut (.I0(GND_net), .I1(n11407[19]), .I2(GND_net), 
            .I3(n44487), .O(n306[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5390_2 (.CI(GND_net), .I0(n35_adj_4932), .I1(n104_adj_4931), 
            .CO(n44273));
    SB_CARRY add_5253_3 (.CI(n44599), .I0(n15956[0]), .I1(n162), .CO(n44600));
    SB_CARRY mult_17_add_1225_22 (.CI(n44487), .I0(n11407[19]), .I1(GND_net), 
            .CO(n44488));
    SB_LUT4 add_5415_13_lut (.I0(GND_net), .I1(n18365[10]), .I2(n910), 
            .I3(n44272), .O(n18053[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5415_12_lut (.I0(GND_net), .I1(n18365[9]), .I2(n837), 
            .I3(n44271), .O(n18053[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5415_12 (.CI(n44271), .I0(n18365[9]), .I1(n837), .CO(n44272));
    SB_LUT4 add_5415_11_lut (.I0(GND_net), .I1(n18365[8]), .I2(n764), 
            .I3(n44270), .O(n18053[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_14 (.CI(n44713), .I0(n11938[11]), .I1(n950), 
            .CO(n44714));
    SB_LUT4 add_5139_8_lut (.I0(GND_net), .I1(n13789[5]), .I2(n518_adj_4922), 
            .I3(n44666), .O(n12908[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5415_11 (.CI(n44270), .I0(n18365[8]), .I1(n764), .CO(n44271));
    SB_LUT4 add_5253_2_lut (.I0(GND_net), .I1(n20), .I2(n89), .I3(GND_net), 
            .O(n15309[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5415_10_lut (.I0(GND_net), .I1(n18365[7]), .I2(n691), 
            .I3(n44269), .O(n18053[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5415_10 (.CI(n44269), .I0(n18365[7]), .I1(n691), .CO(n44270));
    SB_LUT4 mult_16_add_1225_13_lut (.I0(GND_net), .I1(n11938[10]), .I2(n877), 
            .I3(n44712), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_21_lut (.I0(GND_net), .I1(n11407[18]), .I2(GND_net), 
            .I3(n44486), .O(n306[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5415_9_lut (.I0(GND_net), .I1(n18365[6]), .I2(n618), .I3(n44268), 
            .O(n18053[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[23]), 
            .I3(n43424), .O(n436[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[22]), 
            .I3(n43423), .O(n436[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_21 (.CI(n44486), .I0(n11407[18]), .I1(GND_net), 
            .CO(n44487));
    SB_CARRY add_5415_9 (.CI(n44268), .I0(n18365[6]), .I1(n618), .CO(n44269));
    SB_CARRY unary_minus_26_add_3_24 (.CI(n43423), .I0(GND_net), .I1(n1_adj_5416[22]), 
            .CO(n43424));
    SB_LUT4 unary_minus_26_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[21]), 
            .I3(n43422), .O(n436[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_8 (.CI(n44666), .I0(n13789[5]), .I1(n518_adj_4922), 
            .CO(n44667));
    SB_LUT4 add_5139_7_lut (.I0(GND_net), .I1(n13789[4]), .I2(n445_adj_4919), 
            .I3(n44665), .O(n12908[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5415_8_lut (.I0(GND_net), .I1(n18365[5]), .I2(n545), .I3(n44267), 
            .O(n18053[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5415_8 (.CI(n44267), .I0(n18365[5]), .I1(n545), .CO(n44268));
    SB_CARRY unary_minus_26_add_3_23 (.CI(n43422), .I0(GND_net), .I1(n1_adj_5416[21]), 
            .CO(n43423));
    SB_LUT4 unary_minus_26_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[20]), 
            .I3(n43421), .O(n436[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_22 (.CI(n43421), .I0(GND_net), .I1(n1_adj_5416[20]), 
            .CO(n43422));
    SB_CARRY add_5253_2 (.CI(GND_net), .I0(n20), .I1(n89), .CO(n44599));
    SB_LUT4 i28859_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(n4_adj_5348), .I3(n19429[1]), .O(n6_adj_4882));   // verilog/motorControl.v(52[27:38])
    defparam i28859_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_5287_18_lut (.I0(GND_net), .I1(n16533[15]), .I2(GND_net), 
            .I3(n44598), .O(n15956[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_20_lut (.I0(GND_net), .I1(n11407[17]), .I2(GND_net), 
            .I3(n44485), .O(n306[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_20 (.CI(n44485), .I0(n11407[17]), .I1(GND_net), 
            .CO(n44486));
    SB_LUT4 add_5415_7_lut (.I0(GND_net), .I1(n18365[4]), .I2(n472), .I3(n44266), 
            .O(n18053[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5415_7 (.CI(n44266), .I0(n18365[4]), .I1(n472), .CO(n44267));
    SB_LUT4 mult_17_add_1225_19_lut (.I0(GND_net), .I1(n11407[16]), .I2(GND_net), 
            .I3(n44484), .O(n306[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5415_6_lut (.I0(GND_net), .I1(n18365[3]), .I2(n399), .I3(n44265), 
            .O(n18053[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5415_6 (.CI(n44265), .I0(n18365[3]), .I1(n399), .CO(n44266));
    SB_LUT4 add_5415_5_lut (.I0(GND_net), .I1(n18365[2]), .I2(n326), .I3(n44264), 
            .O(n18053[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5287_17_lut (.I0(GND_net), .I1(n16533[14]), .I2(GND_net), 
            .I3(n44597), .O(n15956[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[19]), 
            .I3(n43420), .O(n436[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_21 (.CI(n43420), .I0(GND_net), .I1(n1_adj_5416[19]), 
            .CO(n43421));
    SB_CARRY mult_17_add_1225_19 (.CI(n44484), .I0(n11407[16]), .I1(GND_net), 
            .CO(n44485));
    SB_LUT4 unary_minus_26_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[18]), 
            .I3(n43419), .O(n436[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5415_5 (.CI(n44264), .I0(n18365[2]), .I1(n326), .CO(n44265));
    SB_LUT4 add_5415_4_lut (.I0(GND_net), .I1(n18365[1]), .I2(n253), .I3(n44263), 
            .O(n18053[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_20 (.CI(n43419), .I0(GND_net), .I1(n1_adj_5416[18]), 
            .CO(n43420));
    SB_LUT4 mult_17_add_1225_18_lut (.I0(GND_net), .I1(n11407[15]), .I2(GND_net), 
            .I3(n44483), .O(n306[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_18 (.CI(n44483), .I0(n11407[15]), .I1(GND_net), 
            .CO(n44484));
    SB_CARRY add_5415_4 (.CI(n44263), .I0(n18365[1]), .I1(n253), .CO(n44264));
    SB_LUT4 unary_minus_26_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[17]), 
            .I3(n43418), .O(n436[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5415_3_lut (.I0(GND_net), .I1(n18365[0]), .I2(n180), .I3(n44262), 
            .O(n18053[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_19 (.CI(n43418), .I0(GND_net), .I1(n1_adj_5416[17]), 
            .CO(n43419));
    SB_CARRY add_5415_3 (.CI(n44262), .I0(n18365[0]), .I1(n180), .CO(n44263));
    SB_LUT4 add_5415_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_4911), 
            .I3(GND_net), .O(n18053[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5415_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[16]), 
            .I3(n43417), .O(n436[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_17_lut (.I0(GND_net), .I1(n11407[14]), .I2(GND_net), 
            .I3(n44482), .O(n306[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5287_17 (.CI(n44597), .I0(n16533[14]), .I1(GND_net), 
            .CO(n44598));
    SB_LUT4 add_5287_16_lut (.I0(GND_net), .I1(n16533[13]), .I2(n1114), 
            .I3(n44596), .O(n15956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5415_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_4911), .CO(n44262));
    SB_CARRY mult_17_add_1225_17 (.CI(n44482), .I0(n11407[14]), .I1(GND_net), 
            .CO(n44483));
    SB_LUT4 add_5529_7_lut (.I0(GND_net), .I1(n50780), .I2(n490_adj_4904), 
            .I3(n44261), .O(n19333[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5529_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_18 (.CI(n43417), .I0(GND_net), .I1(n1_adj_5416[16]), 
            .CO(n43418));
    SB_LUT4 mult_17_add_1225_16_lut (.I0(GND_net), .I1(n11407[13]), .I2(n1096), 
            .I3(n44481), .O(n306[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5287_16 (.CI(n44596), .I0(n16533[13]), .I1(n1114), .CO(n44597));
    SB_LUT4 add_5529_6_lut (.I0(GND_net), .I1(n19404[3]), .I2(n417), .I3(n44260), 
            .O(n19333[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5529_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5287_15_lut (.I0(GND_net), .I1(n16533[12]), .I2(n1041), 
            .I3(n44595), .O(n15956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_16 (.CI(n44481), .I0(n11407[13]), .I1(n1096), 
            .CO(n44482));
    SB_LUT4 unary_minus_26_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[15]), 
            .I3(n43416), .O(n436[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5529_6 (.CI(n44260), .I0(n19404[3]), .I1(n417), .CO(n44261));
    SB_CARRY unary_minus_26_add_3_17 (.CI(n43416), .I0(GND_net), .I1(n1_adj_5416[15]), 
            .CO(n43417));
    SB_LUT4 mult_17_add_1225_15_lut (.I0(GND_net), .I1(n11407[12]), .I2(n1023), 
            .I3(n44480), .O(n306[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5529_5_lut (.I0(GND_net), .I1(n19404[2]), .I2(n344), .I3(n44259), 
            .O(n19333[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5529_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[14]), 
            .I3(n43415), .O(n436[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_16 (.CI(n43415), .I0(GND_net), .I1(n1_adj_5416[14]), 
            .CO(n43416));
    SB_CARRY add_5139_7 (.CI(n44665), .I0(n13789[4]), .I1(n445_adj_4919), 
            .CO(n44666));
    SB_CARRY add_5529_5 (.CI(n44259), .I0(n19404[2]), .I1(n344), .CO(n44260));
    SB_LUT4 add_5529_4_lut (.I0(GND_net), .I1(n19404[1]), .I2(n271), .I3(n44258), 
            .O(n19333[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5529_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n43233), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5529_4 (.CI(n44258), .I0(n19404[1]), .I1(n271), .CO(n44259));
    SB_CARRY add_5287_15 (.CI(n44595), .I0(n16533[12]), .I1(n1041), .CO(n44596));
    SB_LUT4 sub_8_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n43232), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_15 (.CI(n44480), .I0(n11407[12]), .I1(n1023), 
            .CO(n44481));
    SB_CARRY sub_8_add_2_24 (.CI(n43232), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n43233));
    SB_LUT4 sub_8_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n43231), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[13]), 
            .I3(n43414), .O(n436[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_23 (.CI(n43231), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n43232));
    SB_CARRY unary_minus_26_add_3_15 (.CI(n43414), .I0(GND_net), .I1(n1_adj_5416[13]), 
            .CO(n43415));
    SB_LUT4 unary_minus_26_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[12]), 
            .I3(n43413), .O(n436[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5529_3_lut (.I0(GND_net), .I1(n19404[0]), .I2(n198_adj_5261), 
            .I3(n44257), .O(n19333[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5529_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5529_3 (.CI(n44257), .I0(n19404[0]), .I1(n198_adj_5261), 
            .CO(n44258));
    SB_CARRY unary_minus_26_add_3_14 (.CI(n43413), .I0(GND_net), .I1(n1_adj_5416[12]), 
            .CO(n43414));
    SB_LUT4 unary_minus_26_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[11]), 
            .I3(n43412), .O(n436[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5529_2_lut (.I0(GND_net), .I1(n56), .I2(n125_adj_5257), 
            .I3(GND_net), .O(n19333[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5529_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n43230), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_13 (.CI(n43412), .I0(GND_net), .I1(n1_adj_5416[11]), 
            .CO(n43413));
    SB_LUT4 unary_minus_26_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[10]), 
            .I3(n43411), .O(n436[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_22 (.CI(n43230), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n43231));
    SB_LUT4 sub_8_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n43229), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_21 (.CI(n43229), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n43230));
    SB_LUT4 sub_8_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n43228), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_14_lut (.I0(GND_net), .I1(n11407[11]), .I2(n950_adj_5248), 
            .I3(n44479), .O(n306[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_20 (.CI(n43228), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n43229));
    SB_CARRY mult_17_add_1225_14 (.CI(n44479), .I0(n11407[11]), .I1(n950_adj_5248), 
            .CO(n44480));
    SB_LUT4 sub_8_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n43227), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5529_2 (.CI(GND_net), .I0(n56), .I1(n125_adj_5257), .CO(n44257));
    SB_CARRY unary_minus_26_add_3_12 (.CI(n43411), .I0(GND_net), .I1(n1_adj_5416[10]), 
            .CO(n43412));
    SB_LUT4 add_5438_12_lut (.I0(GND_net), .I1(n18629[9]), .I2(n840), 
            .I3(n44256), .O(n18365[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5438_11_lut (.I0(GND_net), .I1(n18629[8]), .I2(n767), 
            .I3(n44255), .O(n18365[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_19 (.CI(n43227), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n43228));
    SB_LUT4 add_5139_6_lut (.I0(GND_net), .I1(n13789[3]), .I2(n372_adj_5239), 
            .I3(n44664), .O(n12908[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[9]), 
            .I3(n43410), .O(n436[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5287_14_lut (.I0(GND_net), .I1(n16533[11]), .I2(n968_adj_5234), 
            .I3(n44594), .O(n15956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_11 (.CI(n43410), .I0(GND_net), .I1(n1_adj_5416[9]), 
            .CO(n43411));
    SB_LUT4 mult_17_add_1225_13_lut (.I0(GND_net), .I1(n11407[10]), .I2(n877_adj_5232), 
            .I3(n44478), .O(n306[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5438_11 (.CI(n44255), .I0(n18629[8]), .I1(n767), .CO(n44256));
    SB_LUT4 unary_minus_26_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[8]), 
            .I3(n43409), .O(n436[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n43226), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_18 (.CI(n43226), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n43227));
    SB_LUT4 sub_8_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n43225), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_10 (.CI(n43409), .I0(GND_net), .I1(n1_adj_5416[8]), 
            .CO(n43410));
    SB_CARRY sub_8_add_2_17 (.CI(n43225), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n43226));
    SB_LUT4 unary_minus_26_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[7]), 
            .I3(n43408), .O(n436[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_9 (.CI(n43408), .I0(GND_net), .I1(n1_adj_5416[7]), 
            .CO(n43409));
    SB_LUT4 sub_8_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n43224), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5438_10_lut (.I0(GND_net), .I1(n18629[7]), .I2(n694), 
            .I3(n44254), .O(n18365[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[6]), 
            .I3(n43407), .O(n436[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_8 (.CI(n43407), .I0(GND_net), .I1(n1_adj_5416[6]), 
            .CO(n43408));
    SB_CARRY sub_8_add_2_16 (.CI(n43224), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n43225));
    SB_CARRY add_5438_10 (.CI(n44254), .I0(n18629[7]), .I1(n694), .CO(n44255));
    SB_LUT4 add_5438_9_lut (.I0(GND_net), .I1(n18629[6]), .I2(n621), .I3(n44253), 
            .O(n18365[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5438_9 (.CI(n44253), .I0(n18629[6]), .I1(n621), .CO(n44254));
    SB_LUT4 add_5438_8_lut (.I0(GND_net), .I1(n18629[5]), .I2(n548), .I3(n44252), 
            .O(n18365[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[5]), 
            .I3(n43406), .O(n436[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5438_8 (.CI(n44252), .I0(n18629[5]), .I1(n548), .CO(n44253));
    SB_CARRY mult_17_add_1225_13 (.CI(n44478), .I0(n11407[10]), .I1(n877_adj_5232), 
            .CO(n44479));
    SB_CARRY add_5287_14 (.CI(n44594), .I0(n16533[11]), .I1(n968_adj_5234), 
            .CO(n44595));
    SB_LUT4 add_5438_7_lut (.I0(GND_net), .I1(n18629[4]), .I2(n475), .I3(n44251), 
            .O(n18365[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_7 (.CI(n43406), .I0(GND_net), .I1(n1_adj_5416[5]), 
            .CO(n43407));
    SB_LUT4 unary_minus_26_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[4]), 
            .I3(n43405), .O(n436[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_6 (.CI(n43405), .I0(GND_net), .I1(n1_adj_5416[4]), 
            .CO(n43406));
    SB_LUT4 unary_minus_26_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[3]), 
            .I3(n43404), .O(n436[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n43223), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5438_7 (.CI(n44251), .I0(n18629[4]), .I1(n475), .CO(n44252));
    SB_CARRY unary_minus_26_add_3_5 (.CI(n43404), .I0(GND_net), .I1(n1_adj_5416[3]), 
            .CO(n43405));
    SB_LUT4 mult_17_add_1225_12_lut (.I0(GND_net), .I1(n11407[9]), .I2(n804_adj_5218), 
            .I3(n44477), .O(n306[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[2]), 
            .I3(n43403), .O(n436[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_4 (.CI(n43403), .I0(GND_net), .I1(n1_adj_5416[2]), 
            .CO(n43404));
    SB_CARRY sub_8_add_2_15 (.CI(n43223), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n43224));
    SB_LUT4 unary_minus_26_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[1]), 
            .I3(n43402), .O(n436[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5287_13_lut (.I0(GND_net), .I1(n16533[10]), .I2(n895_adj_5212), 
            .I3(n44593), .O(n15956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_3 (.CI(n43402), .I0(GND_net), .I1(n1_adj_5416[1]), 
            .CO(n43403));
    SB_LUT4 sub_8_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n43222), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_14 (.CI(n43222), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n43223));
    SB_LUT4 unary_minus_26_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5416[0]), 
            .I3(VCC_net), .O(n436[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_12 (.CI(n44477), .I0(n11407[9]), .I1(n804_adj_5218), 
            .CO(n44478));
    SB_LUT4 sub_8_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n43221), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_13 (.CI(n43221), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n43222));
    SB_LUT4 mult_17_add_1225_11_lut (.I0(GND_net), .I1(n11407[8]), .I2(n731_adj_5202), 
            .I3(n44476), .O(n306[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_13 (.CI(n44712), .I0(n11938[10]), .I1(n877), 
            .CO(n44713));
    SB_CARRY unary_minus_26_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5416[0]), 
            .CO(n43402));
    SB_LUT4 sub_8_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n43220), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(n356[23]), .I1(GND_net), .I2(n1_adj_5418[23]), 
            .I3(n43401), .O(n47_adj_5269)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY sub_8_add_2_12 (.CI(n43220), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n43221));
    SB_CARRY add_5139_6 (.CI(n44664), .I0(n13789[3]), .I1(n372_adj_5239), 
            .CO(n44665));
    SB_LUT4 sub_8_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n43219), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5438_6_lut (.I0(GND_net), .I1(n18629[3]), .I2(n402_adj_5195), 
            .I3(n44250), .O(n18365[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5438_6 (.CI(n44250), .I0(n18629[3]), .I1(n402_adj_5195), 
            .CO(n44251));
    SB_CARRY sub_8_add_2_11 (.CI(n43219), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n43220));
    SB_LUT4 add_5438_5_lut (.I0(GND_net), .I1(n18629[2]), .I2(n329_adj_5194), 
            .I3(n44249), .O(n18365[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[22]), 
            .I3(n43400), .O(n382[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n43400), .I0(GND_net), .I1(n1_adj_5418[22]), 
            .CO(n43401));
    SB_CARRY add_5287_13 (.CI(n44593), .I0(n16533[10]), .I1(n895_adj_5212), 
            .CO(n44594));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[21]), 
            .I3(n43399), .O(n382[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5438_5 (.CI(n44249), .I0(n18629[2]), .I1(n329_adj_5194), 
            .CO(n44250));
    SB_LUT4 add_5287_12_lut (.I0(GND_net), .I1(n16533[9]), .I2(n822_adj_5189), 
            .I3(n44592), .O(n15956[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5438_4_lut (.I0(GND_net), .I1(n18629[1]), .I2(n256_adj_5188), 
            .I3(n44248), .O(n18365[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n43399), .I0(GND_net), .I1(n1_adj_5418[21]), 
            .CO(n43400));
    SB_LUT4 sub_8_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n43218), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5438_4 (.CI(n44248), .I0(n18629[1]), .I1(n256_adj_5188), 
            .CO(n44249));
    SB_CARRY mult_17_add_1225_11 (.CI(n44476), .I0(n11407[8]), .I1(n731_adj_5202), 
            .CO(n44477));
    SB_CARRY sub_8_add_2_10 (.CI(n43218), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n43219));
    SB_LUT4 mult_17_add_1225_10_lut (.I0(GND_net), .I1(n11407[7]), .I2(n658_adj_5186), 
            .I3(n44475), .O(n306[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n43217), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[20]), 
            .I3(n43398), .O(n382[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_9 (.CI(n43217), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n43218));
    SB_CARRY unary_minus_20_add_3_22 (.CI(n43398), .I0(GND_net), .I1(n1_adj_5418[20]), 
            .CO(n43399));
    SB_LUT4 sub_8_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n43216), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5438_3_lut (.I0(GND_net), .I1(n18629[0]), .I2(n183_adj_5163), 
            .I3(n44247), .O(n18365[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[19]), 
            .I3(n43397), .O(n382[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5438_3 (.CI(n44247), .I0(n18629[0]), .I1(n183_adj_5163), 
            .CO(n44248));
    SB_CARRY unary_minus_20_add_3_21 (.CI(n43397), .I0(GND_net), .I1(n1_adj_5418[19]), 
            .CO(n43398));
    SB_CARRY mult_17_add_1225_10 (.CI(n44475), .I0(n11407[7]), .I1(n658_adj_5186), 
            .CO(n44476));
    SB_LUT4 add_5438_2_lut (.I0(GND_net), .I1(n41_adj_5156), .I2(n110_adj_5153), 
            .I3(GND_net), .O(n18365[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5438_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[18]), 
            .I3(n43396), .O(n382[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_8 (.CI(n43216), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n43217));
    SB_CARRY unary_minus_20_add_3_20 (.CI(n43396), .I0(GND_net), .I1(n1_adj_5418[18]), 
            .CO(n43397));
    SB_LUT4 sub_8_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n43215), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[17]), 
            .I3(n43395), .O(n382[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_7 (.CI(n43215), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n43216));
    SB_CARRY add_5438_2 (.CI(GND_net), .I0(n41_adj_5156), .I1(n110_adj_5153), 
            .CO(n44247));
    SB_LUT4 add_5139_5_lut (.I0(GND_net), .I1(n13789[2]), .I2(n299_adj_5143), 
            .I3(n44663), .O(n12908[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n43395), .I0(GND_net), .I1(n1_adj_5418[17]), 
            .CO(n43396));
    SB_LUT4 sub_8_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n43214), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[16]), 
            .I3(n43394), .O(n382[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_18 (.CI(n43394), .I0(GND_net), .I1(n1_adj_5418[16]), 
            .CO(n43395));
    SB_LUT4 mult_17_add_1225_9_lut (.I0(GND_net), .I1(n11407[6]), .I2(n585), 
            .I3(n44474), .O(n306[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[15]), 
            .I3(n43393), .O(n382[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_17 (.CI(n43393), .I0(GND_net), .I1(n1_adj_5418[15]), 
            .CO(n43394));
    SB_CARRY mult_17_add_1225_9 (.CI(n44474), .I0(n11407[6]), .I1(n585), 
            .CO(n44475));
    SB_CARRY sub_8_add_2_6 (.CI(n43214), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n43215));
    SB_CARRY add_5287_12 (.CI(n44592), .I0(n16533[9]), .I1(n822_adj_5189), 
            .CO(n44593));
    SB_LUT4 mult_16_add_1225_12_lut (.I0(GND_net), .I1(n11938[9]), .I2(n804), 
            .I3(n44711), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n43213), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_5 (.CI(n44663), .I0(n13789[2]), .I1(n299_adj_5143), 
            .CO(n44664));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[14]), 
            .I3(n43392), .O(n382[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_16 (.CI(n43392), .I0(GND_net), .I1(n1_adj_5418[14]), 
            .CO(n43393));
    SB_LUT4 add_5287_11_lut (.I0(GND_net), .I1(n16533[8]), .I2(n749_adj_5124), 
            .I3(n44591), .O(n15956[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_8_lut (.I0(GND_net), .I1(n11407[5]), .I2(n512_adj_5112), 
            .I3(n44473), .O(n306[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_8 (.CI(n44473), .I0(n11407[5]), .I1(n512_adj_5112), 
            .CO(n44474));
    SB_CARRY sub_8_add_2_5 (.CI(n43213), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n43214));
    SB_LUT4 mult_17_add_1225_7_lut (.I0(GND_net), .I1(n11407[4]), .I2(n439_adj_5111), 
            .I3(n44472), .O(n306[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[13]), 
            .I3(n43391), .O(n382[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n43391), .I0(GND_net), .I1(n1_adj_5418[13]), 
            .CO(n43392));
    SB_CARRY add_5287_11 (.CI(n44591), .I0(n16533[8]), .I1(n749_adj_5124), 
            .CO(n44592));
    SB_LUT4 sub_8_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n43212), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[12]), 
            .I3(n43390), .O(n382[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_4 (.CI(n43212), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n43213));
    SB_CARRY unary_minus_20_add_3_14 (.CI(n43390), .I0(GND_net), .I1(n1_adj_5418[12]), 
            .CO(n43391));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[11]), 
            .I3(n43389), .O(n382[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n43389), .I0(GND_net), .I1(n1_adj_5418[11]), 
            .CO(n43390));
    SB_LUT4 sub_8_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n43211), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_3 (.CI(n43211), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n43212));
    SB_CARRY mult_17_add_1225_7 (.CI(n44472), .I0(n11407[4]), .I1(n439_adj_5111), 
            .CO(n44473));
    SB_LUT4 sub_8_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk16MHz), .D(n29804));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk16MHz), .D(n29803));   // verilog/motorControl.v(43[14] 63[8])
    SB_CARRY sub_8_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n43211));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[10]), 
            .I3(n43388), .O(n382[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n43388), .I0(GND_net), .I1(n1_adj_5418[10]), 
            .CO(n43389));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[9]), 
            .I3(n43387), .O(n382[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n43387), .I0(GND_net), .I1(n1_adj_5418[9]), 
            .CO(n43388));
    SB_DFF \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk16MHz), .D(n29802));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 i1_3_lut_4_lut_adj_1713 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(n4_adj_5348), .I3(n19429[1]), .O(n19369[2]));   // verilog/motorControl.v(52[27:38])
    defparam i1_3_lut_4_lut_adj_1713.LUT_INIT = 16'h8778;
    SB_DFF \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk16MHz), .D(n29801));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk16MHz), .D(n29800));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[8]), 
            .I3(n43386), .O(n382[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n43386), .I0(GND_net), .I1(n1_adj_5418[8]), 
            .CO(n43387));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[7]), 
            .I3(n43385), .O(n382[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n43385), .I0(GND_net), .I1(n1_adj_5418[7]), 
            .CO(n43386));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[6]), 
            .I3(n43384), .O(n382[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n43384), .I0(GND_net), .I1(n1_adj_5418[6]), 
            .CO(n43385));
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[5]), 
            .I3(n43383), .O(n382[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_4_lut (.I0(GND_net), .I1(n13789[1]), .I2(n226_adj_5068), 
            .I3(n44662), .O(n12908[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk16MHz), .D(n29799));   // verilog/motorControl.v(43[14] 63[8])
    SB_CARRY unary_minus_20_add_3_7 (.CI(n43383), .I0(GND_net), .I1(n1_adj_5418[5]), 
            .CO(n43384));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[4]), 
            .I3(n43382), .O(n382[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n43382), .I0(GND_net), .I1(n1_adj_5418[4]), 
            .CO(n43383));
    SB_LUT4 add_5287_10_lut (.I0(GND_net), .I1(n16533[7]), .I2(n676), 
            .I3(n44590), .O(n15956[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[3]), 
            .I3(n43381), .O(n382[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk16MHz), .D(n29798));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk16MHz), .D(n29797));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk16MHz), .D(n29796));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 mult_17_add_1225_6_lut (.I0(GND_net), .I1(n11407[3]), .I2(n366_adj_5054), 
            .I3(n44471), .O(n306[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5287_10 (.CI(n44590), .I0(n16533[7]), .I1(n676), .CO(n44591));
    SB_CARRY mult_16_add_1225_12 (.CI(n44711), .I0(n11938[9]), .I1(n804), 
            .CO(n44712));
    SB_CARRY add_5139_4 (.CI(n44662), .I0(n13789[1]), .I1(n226_adj_5068), 
            .CO(n44663));
    SB_CARRY unary_minus_20_add_3_5 (.CI(n43381), .I0(GND_net), .I1(n1_adj_5418[3]), 
            .CO(n43382));
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[2]), 
            .I3(n43380), .O(n382[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_6 (.CI(n44471), .I0(n11407[3]), .I1(n366_adj_5054), 
            .CO(n44472));
    SB_LUT4 add_5287_9_lut (.I0(GND_net), .I1(n16533[6]), .I2(n603), .I3(n44589), 
            .O(n15956[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_5_lut (.I0(GND_net), .I1(n11407[2]), .I2(n293_adj_5044), 
            .I3(n44470), .O(n306[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_5 (.CI(n44470), .I0(n11407[2]), .I1(n293_adj_5044), 
            .CO(n44471));
    SB_CARRY unary_minus_20_add_3_4 (.CI(n43380), .I0(GND_net), .I1(n1_adj_5418[2]), 
            .CO(n43381));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5418[1]), 
            .I3(n43379), .O(n382[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_4_lut (.I0(GND_net), .I1(n11407[1]), .I2(n220_adj_5040), 
            .I3(n44469), .O(n306[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_4 (.CI(n44469), .I0(n11407[1]), .I1(n220_adj_5040), 
            .CO(n44470));
    SB_LUT4 i38780_2_lut_4_lut (.I0(n130[21]), .I1(n182[21]), .I2(n130[9]), 
            .I3(n182[9]), .O(n54573));
    defparam i38780_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n43379), .I0(GND_net), .I1(n1_adj_5418[1]), 
            .CO(n43380));
    SB_DFF \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk16MHz), .D(n29795));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk16MHz), .D(n29794));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk16MHz), .D(n29793));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(n36533), .I1(GND_net), .I2(n1_adj_5418[0]), 
            .I3(VCC_net), .O(n54263)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5418[0]), 
            .CO(n43379));
    SB_LUT4 i38790_2_lut_4_lut (.I0(n130[16]), .I1(n182[16]), .I2(n130[7]), 
            .I3(n182[7]), .O(n54583));
    defparam i38790_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_13_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[23]), 
            .I3(n43378), .O(n182[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[22]), 
            .I3(n43377), .O(n182[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_24 (.CI(n43377), .I0(GND_net), .I1(n1_adj_5417[22]), 
            .CO(n43378));
    SB_LUT4 unary_minus_13_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[21]), 
            .I3(n43376), .O(n182[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_3_lut (.I0(GND_net), .I1(n11407[0]), .I2(n147_adj_5024), 
            .I3(n44468), .O(n306[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_3 (.CI(n44468), .I0(n11407[0]), .I1(n147_adj_5024), 
            .CO(n44469));
    SB_CARRY unary_minus_13_add_3_23 (.CI(n43376), .I0(GND_net), .I1(n1_adj_5417[21]), 
            .CO(n43377));
    SB_LUT4 unary_minus_13_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[20]), 
            .I3(n43375), .O(n182[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_22 (.CI(n43375), .I0(GND_net), .I1(n1_adj_5417[20]), 
            .CO(n43376));
    SB_DFF \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk16MHz), .D(n29792));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk16MHz), .D(n29791));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk16MHz), .D(n29790));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 unary_minus_13_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[19]), 
            .I3(n43374), .O(n182[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_21 (.CI(n43374), .I0(GND_net), .I1(n1_adj_5417[19]), 
            .CO(n43375));
    SB_LUT4 unary_minus_13_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[18]), 
            .I3(n43373), .O(n182[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_20 (.CI(n43373), .I0(GND_net), .I1(n1_adj_5417[18]), 
            .CO(n43374));
    SB_LUT4 add_5139_3_lut (.I0(GND_net), .I1(n13789[0]), .I2(n153_adj_5020), 
            .I3(n44661), .O(n12908[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[17]), 
            .I3(n43372), .O(n182[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_19 (.CI(n43372), .I0(GND_net), .I1(n1_adj_5417[17]), 
            .CO(n43373));
    SB_LUT4 unary_minus_13_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[16]), 
            .I3(n43371), .O(n182[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_18 (.CI(n43371), .I0(GND_net), .I1(n1_adj_5417[16]), 
            .CO(n43372));
    SB_DFF \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk16MHz), .D(n29789));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk16MHz), .D(n29788));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk16MHz), .D(n29787));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 unary_minus_13_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[15]), 
            .I3(n43370), .O(n182[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_17 (.CI(n43370), .I0(GND_net), .I1(n1_adj_5417[15]), 
            .CO(n43371));
    SB_LUT4 unary_minus_13_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[14]), 
            .I3(n43369), .O(n182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_11_lut (.I0(GND_net), .I1(n11938[8]), .I2(n731), 
            .I3(n44710), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_3 (.CI(n44661), .I0(n13789[0]), .I1(n153_adj_5020), 
            .CO(n44662));
    SB_CARRY add_5287_9 (.CI(n44589), .I0(n16533[6]), .I1(n603), .CO(n44590));
    SB_LUT4 add_5139_2_lut (.I0(GND_net), .I1(n11_adj_5014), .I2(n80_adj_5012), 
            .I3(GND_net), .O(n12908[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5287_8_lut (.I0(GND_net), .I1(n16533[5]), .I2(n530), .I3(n44588), 
            .O(n15956[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_5011), .I2(n74_adj_5009), 
            .I3(GND_net), .O(n306[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_2 (.CI(GND_net), .I0(n5_adj_5011), .I1(n74_adj_5009), 
            .CO(n44468));
    SB_CARRY unary_minus_13_add_3_16 (.CI(n43369), .I0(GND_net), .I1(n1_adj_5417[14]), 
            .CO(n43370));
    SB_LUT4 add_5073_23_lut (.I0(GND_net), .I1(n12425[20]), .I2(GND_net), 
            .I3(n44467), .O(n11407[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk16MHz), .D(n29786));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk16MHz), .D(n29785));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 unary_minus_13_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[13]), 
            .I3(n43368), .O(n182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_15 (.CI(n43368), .I0(GND_net), .I1(n1_adj_5417[13]), 
            .CO(n43369));
    SB_LUT4 unary_minus_13_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[12]), 
            .I3(n43367), .O(n182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_14 (.CI(n43367), .I0(GND_net), .I1(n1_adj_5417[12]), 
            .CO(n43368));
    SB_LUT4 unary_minus_13_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[11]), 
            .I3(n43366), .O(n182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_13 (.CI(n43366), .I0(GND_net), .I1(n1_adj_5417[11]), 
            .CO(n43367));
    SB_LUT4 unary_minus_13_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[10]), 
            .I3(n43365), .O(n182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_12 (.CI(n43365), .I0(GND_net), .I1(n1_adj_5417[10]), 
            .CO(n43366));
    SB_LUT4 unary_minus_13_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[9]), 
            .I3(n43364), .O(n182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_11 (.CI(n43364), .I0(GND_net), .I1(n1_adj_5417[9]), 
            .CO(n43365));
    SB_LUT4 unary_minus_13_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[8]), 
            .I3(n43363), .O(n182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5073_22_lut (.I0(GND_net), .I1(n12425[19]), .I2(GND_net), 
            .I3(n44466), .O(n11407[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_10 (.CI(n43363), .I0(GND_net), .I1(n1_adj_5417[8]), 
            .CO(n43364));
    SB_LUT4 unary_minus_13_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[7]), 
            .I3(n43362), .O(n182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_9 (.CI(n43362), .I0(GND_net), .I1(n1_adj_5417[7]), 
            .CO(n43363));
    SB_DFF \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk16MHz), .D(n29784));   // verilog/motorControl.v(43[14] 63[8])
    SB_CARRY add_5073_22 (.CI(n44466), .I0(n12425[19]), .I1(GND_net), 
            .CO(n44467));
    SB_CARRY add_5287_8 (.CI(n44588), .I0(n16533[5]), .I1(n530), .CO(n44589));
    SB_LUT4 add_5073_21_lut (.I0(GND_net), .I1(n12425[18]), .I2(GND_net), 
            .I3(n44465), .O(n11407[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_21 (.CI(n44465), .I0(n12425[18]), .I1(GND_net), 
            .CO(n44466));
    SB_LUT4 unary_minus_13_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[6]), 
            .I3(n43361), .O(n182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_8 (.CI(n43361), .I0(GND_net), .I1(n1_adj_5417[6]), 
            .CO(n43362));
    SB_LUT4 unary_minus_13_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[5]), 
            .I3(n43360), .O(n182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_2 (.CI(GND_net), .I0(n11_adj_5014), .I1(n80_adj_5012), 
            .CO(n44661));
    SB_LUT4 add_5179_21_lut (.I0(GND_net), .I1(n14588[18]), .I2(GND_net), 
            .I3(n44660), .O(n13789[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5287_7_lut (.I0(GND_net), .I1(n16533[4]), .I2(n457_adj_4987), 
            .I3(n44587), .O(n15956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_7 (.CI(n43360), .I0(GND_net), .I1(n1_adj_5417[5]), 
            .CO(n43361));
    SB_CARRY add_5287_7 (.CI(n44587), .I0(n16533[4]), .I1(n457_adj_4987), 
            .CO(n44588));
    SB_LUT4 add_5073_20_lut (.I0(GND_net), .I1(n12425[17]), .I2(GND_net), 
            .I3(n44464), .O(n11407[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_20 (.CI(n44464), .I0(n12425[17]), .I1(GND_net), 
            .CO(n44465));
    SB_DFF \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk16MHz), .D(n29783));   // verilog/motorControl.v(43[14] 63[8])
    SB_DFF \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk16MHz), .D(n29782));   // verilog/motorControl.v(43[14] 63[8])
    SB_LUT4 i38814_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n130[21]), .I2(IntegralLimit[9]), 
            .I3(n130[9]), .O(n54607));
    defparam i38814_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5287_6_lut (.I0(GND_net), .I1(n16533[3]), .I2(n384), .I3(n44586), 
            .O(n15956[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5073_19_lut (.I0(GND_net), .I1(n12425[16]), .I2(GND_net), 
            .I3(n44463), .O(n11407[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[4]), 
            .I3(n43359), .O(n182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_6 (.CI(n43359), .I0(GND_net), .I1(n1_adj_5417[4]), 
            .CO(n43360));
    SB_LUT4 unary_minus_13_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[3]), 
            .I3(n43358), .O(n182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_5 (.CI(n43358), .I0(GND_net), .I1(n1_adj_5417[3]), 
            .CO(n43359));
    SB_LUT4 unary_minus_13_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[2]), 
            .I3(n43357), .O(n182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_4 (.CI(n43357), .I0(GND_net), .I1(n1_adj_5417[2]), 
            .CO(n43358));
    SB_LUT4 unary_minus_13_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[1]), 
            .I3(n43356), .O(n182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_3 (.CI(n43356), .I0(GND_net), .I1(n1_adj_5417[1]), 
            .CO(n43357));
    SB_LUT4 unary_minus_13_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5417[0]), 
            .I3(VCC_net), .O(n182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5417[0]), 
            .CO(n43356));
    SB_LUT4 i38824_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n130[16]), .I2(IntegralLimit[7]), 
            .I3(n130[7]), .O(n54617));
    defparam i38824_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5073_19 (.CI(n44463), .I0(n12425[16]), .I1(GND_net), 
            .CO(n44464));
    SB_LUT4 add_5073_18_lut (.I0(GND_net), .I1(n12425[15]), .I2(GND_net), 
            .I3(n44462), .O(n11407[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5287_6 (.CI(n44586), .I0(n16533[3]), .I1(n384), .CO(n44587));
    SB_CARRY add_5073_18 (.CI(n44462), .I0(n12425[15]), .I1(GND_net), 
            .CO(n44463));
    SB_LUT4 add_5073_17_lut (.I0(GND_net), .I1(n12425[14]), .I2(GND_net), 
            .I3(n44461), .O(n11407[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_11 (.CI(n44710), .I0(n11938[8]), .I1(n731), 
            .CO(n44711));
    SB_LUT4 add_5179_20_lut (.I0(GND_net), .I1(n14588[17]), .I2(GND_net), 
            .I3(n44659), .O(n13789[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5287_5_lut (.I0(GND_net), .I1(n16533[2]), .I2(n311), .I3(n44585), 
            .O(n15956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_17 (.CI(n44461), .I0(n12425[14]), .I1(GND_net), 
            .CO(n44462));
    SB_LUT4 add_5073_16_lut (.I0(GND_net), .I1(n12425[13]), .I2(n1099_adj_4956), 
            .I3(n44460), .O(n11407[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5287_5 (.CI(n44585), .I0(n16533[2]), .I1(n311), .CO(n44586));
    SB_CARRY add_5073_16 (.CI(n44460), .I0(n12425[13]), .I1(n1099_adj_4956), 
            .CO(n44461));
    SB_LUT4 add_5073_15_lut (.I0(GND_net), .I1(n12425[12]), .I2(n1026_adj_4948), 
            .I3(n44459), .O(n11407[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_20 (.CI(n44659), .I0(n14588[17]), .I1(GND_net), 
            .CO(n44660));
    SB_LUT4 add_5287_4_lut (.I0(GND_net), .I1(n16533[1]), .I2(n238), .I3(n44584), 
            .O(n15956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_15 (.CI(n44459), .I0(n12425[12]), .I1(n1026_adj_4948), 
            .CO(n44460));
    SB_CARRY add_5287_4 (.CI(n44584), .I0(n16533[1]), .I1(n238), .CO(n44585));
    SB_LUT4 add_5073_14_lut (.I0(GND_net), .I1(n12425[11]), .I2(n953_adj_4942), 
            .I3(n44458), .O(n11407[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5287_3_lut (.I0(GND_net), .I1(n16533[0]), .I2(n165), .I3(n44583), 
            .O(n15956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i247_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5073_14 (.CI(n44458), .I0(n12425[11]), .I1(n953_adj_4942), 
            .CO(n44459));
    SB_LUT4 add_5073_13_lut (.I0(GND_net), .I1(n12425[10]), .I2(n880_adj_4940), 
            .I3(n44457), .O(n11407[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5179_19_lut (.I0(GND_net), .I1(n14588[16]), .I2(GND_net), 
            .I3(n44658), .O(n13789[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38812_3_lut_4_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(n130[2]), .O(n54605));   // verilog/motorControl.v(49[21:44])
    defparam i38812_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5073_13 (.CI(n44457), .I0(n12425[10]), .I1(n880_adj_4940), 
            .CO(n44458));
    SB_CARRY add_5287_3 (.CI(n44583), .I0(n16533[0]), .I1(n165), .CO(n44584));
    SB_LUT4 add_5073_12_lut (.I0(GND_net), .I1(n12425[9]), .I2(n807_adj_4927), 
            .I3(n44456), .O(n11407[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5287_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n15956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5287_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i6_3_lut_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(GND_net), .O(n6_adj_5351));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_5073_12 (.CI(n44456), .I0(n12425[9]), .I1(n807_adj_4927), 
            .CO(n44457));
    SB_LUT4 mult_16_add_1225_10_lut (.I0(GND_net), .I1(n11938[7]), .I2(n658), 
            .I3(n44709), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5073_11_lut (.I0(GND_net), .I1(n12425[8]), .I2(n734_adj_4898), 
            .I3(n44455), .O(n11407[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_19 (.CI(n44658), .I0(n14588[16]), .I1(GND_net), 
            .CO(n44659));
    SB_CARRY add_5287_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n44583));
    SB_CARRY add_5073_11 (.CI(n44455), .I0(n12425[8]), .I1(n734_adj_4898), 
            .CO(n44456));
    SB_LUT4 add_5073_10_lut (.I0(GND_net), .I1(n12425[7]), .I2(n661_adj_4878), 
            .I3(n44454), .O(n11407[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5179_18_lut (.I0(GND_net), .I1(n14588[15]), .I2(GND_net), 
            .I3(n44657), .O(n13789[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5179_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38847_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n130[3]), .I2(n130[2]), 
            .I3(IntegralLimit[2]), .O(n54640));   // verilog/motorControl.v(47[12:34])
    defparam i38847_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5495_9_lut (.I0(GND_net), .I1(n19173[6]), .I2(n630_adj_5352), 
            .I3(n44582), .O(n19029[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_10 (.CI(n44454), .I0(n12425[7]), .I1(n661_adj_4878), 
            .CO(n44455));
    SB_LUT4 add_5073_9_lut (.I0(GND_net), .I1(n12425[6]), .I2(n588_adj_5353), 
            .I3(n44453), .O(n11407[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_9 (.CI(n44453), .I0(n12425[6]), .I1(n588_adj_5353), 
            .CO(n44454));
    SB_LUT4 LessThan_10_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n130[3]), 
            .I2(n130[2]), .I3(GND_net), .O(n6_adj_5354));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY mult_16_add_1225_10 (.CI(n44709), .I0(n11938[7]), .I1(n658), 
            .CO(n44710));
    SB_LUT4 add_5073_8_lut (.I0(GND_net), .I1(n12425[5]), .I2(n515_adj_5355), 
            .I3(n44452), .O(n11407[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5495_8_lut (.I0(GND_net), .I1(n19173[5]), .I2(n557_adj_5356), 
            .I3(n44581), .O(n19029[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_8 (.CI(n44452), .I0(n12425[5]), .I1(n515_adj_5355), 
            .CO(n44453));
    SB_LUT4 add_5073_7_lut (.I0(GND_net), .I1(n12425[4]), .I2(n442_adj_5357), 
            .I3(n44451), .O(n11407[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_9_lut (.I0(GND_net), .I1(n11938[6]), .I2(n585_adj_5358), 
            .I3(n44708), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5179_18 (.CI(n44657), .I0(n14588[15]), .I1(GND_net), 
            .CO(n44658));
    SB_CARRY add_5495_8 (.CI(n44581), .I0(n19173[5]), .I1(n557_adj_5356), 
            .CO(n44582));
    SB_CARRY add_5073_7 (.CI(n44451), .I0(n12425[4]), .I1(n442_adj_5357), 
            .CO(n44452));
    SB_LUT4 add_5073_6_lut (.I0(GND_net), .I1(n12425[3]), .I2(n369_adj_5359), 
            .I3(n44450), .O(n11407[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_6 (.CI(n44450), .I0(n12425[3]), .I1(n369_adj_5359), 
            .CO(n44451));
    SB_CARRY mult_16_add_1225_9 (.CI(n44708), .I0(n11938[6]), .I1(n585_adj_5358), 
            .CO(n44709));
    SB_LUT4 add_5073_5_lut (.I0(GND_net), .I1(n12425[2]), .I2(n296), .I3(n44449), 
            .O(n11407[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_5347));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_5346));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_5345));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_5344));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_5343));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_5342));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28981_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_5360), 
            .I3(n19453[1]), .O(n6));   // verilog/motorControl.v(52[18:24])
    defparam i28981_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_1714 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n19453[1]), 
            .I3(n4_adj_5360), .O(n19404[2]));   // verilog/motorControl.v(52[18:24])
    defparam i1_3_lut_4_lut_adj_1714.LUT_INIT = 16'h8778;
    SB_LUT4 mult_17_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i17_3_lut (.I0(n130[16]), .I1(n182[16]), .I2(n181), 
            .I3(GND_net), .O(n207[16]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i17_3_lut (.I0(n207[16]), .I1(IntegralLimit[16]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [16]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_5341));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_5340));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_5339));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_5338));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_5337));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_5336));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_5335));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_5097));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_5096));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_5095));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_5094));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_5334));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_5333));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_5332));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_5331));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_5330));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_5329));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_5328));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_5327));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_5326));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_5325));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i10_3_lut (.I0(n130[9]), .I1(n182[9]), .I2(n181), .I3(GND_net), 
            .O(n207[9]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i10_3_lut (.I0(n207[9]), .I1(IntegralLimit[9]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [9]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_5324));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5323));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_5322));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_5321));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_5320));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_5319));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_5318));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_5317));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_5316));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_5315));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1715 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n19453[0]), 
            .I3(n43040), .O(n19404[1]));   // verilog/motorControl.v(52[18:24])
    defparam i1_3_lut_4_lut_adj_1715.LUT_INIT = 16'h8778;
    SB_LUT4 i28973_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n43040), 
            .I3(n19453[0]), .O(n4_adj_5360));   // verilog/motorControl.v(52[18:24])
    defparam i28973_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_16_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_5314));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_5313));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_5312));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_5311));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_5310));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28960_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n19404[0]));   // verilog/motorControl.v(52[18:24])
    defparam i28960_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i28962_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n43040));   // verilog/motorControl.v(52[18:24])
    defparam i28962_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38778_3_lut_4_lut (.I0(deadband[3]), .I1(n356[3]), .I2(n356[2]), 
            .I3(deadband[2]), .O(n54571));   // verilog/motorControl.v(53[12:29])
    defparam i38778_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n356[3]), 
            .I2(n356[2]), .I3(GND_net), .O(n6_adj_5258));   // verilog/motorControl.v(53[12:29])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_17_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_5309));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_5308));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38754_2_lut_4_lut (.I0(deadband[16]), .I1(n356[16]), .I2(deadband[7]), 
            .I3(n356[7]), .O(n54547));
    defparam i38754_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i38605_3_lut_4_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(n356[2]), .O(n54398));   // verilog/motorControl.v(56[23:39])
    defparam i38605_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_25_i6_3_lut_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(GND_net), .O(n6_adj_5084));   // verilog/motorControl.v(56[23:39])
    defparam LessThan_25_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_16_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_5307));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_5306));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_5305));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38691_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n356[3]), .I2(n356[2]), 
            .I3(PWMLimit[2]), .O(n54484));   // verilog/motorControl.v(54[14:29])
    defparam i38691_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_23_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n356[3]), 
            .I2(n356[2]), .I3(GND_net), .O(n6_adj_5006));   // verilog/motorControl.v(54[14:29])
    defparam LessThan_23_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i14551_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28621), 
            .I3(PWMLimit[0]), .O(n28622));
    defparam i14551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14868_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28938), 
            .I3(PWMLimit[1]), .O(n28939));
    defparam i14868_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14758_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28828), 
            .I3(PWMLimit[23]), .O(n28829));
    defparam i14758_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_14_i3_3_lut (.I0(n130[2]), .I1(n182[2]), .I2(n181), .I3(GND_net), 
            .O(n207[2]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i3_3_lut (.I0(n207[2]), .I1(IntegralLimit[2]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [2]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14763_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28833), 
            .I3(PWMLimit[22]), .O(n28834));
    defparam i14763_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_17_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14768_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28838), 
            .I3(PWMLimit[21]), .O(n28839));
    defparam i14768_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14773_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28843), 
            .I3(PWMLimit[20]), .O(n28844));
    defparam i14773_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14778_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28848), 
            .I3(PWMLimit[19]), .O(n28849));
    defparam i14778_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14783_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28853), 
            .I3(PWMLimit[18]), .O(n28854));
    defparam i14783_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14788_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28858), 
            .I3(PWMLimit[17]), .O(n28859));
    defparam i14788_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_4_lut_adj_1716 (.I0(n62), .I1(n131), .I2(n201_adj_5362), 
            .I3(n42908), .O(n19369[1]));   // verilog/motorControl.v(52[27:38])
    defparam i1_3_lut_4_lut_adj_1716.LUT_INIT = 16'h6996;
    SB_LUT4 i14793_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28863), 
            .I3(PWMLimit[16]), .O(n28864));
    defparam i14793_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14798_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28868), 
            .I3(PWMLimit[15]), .O(n28869));
    defparam i14798_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14803_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28873), 
            .I3(PWMLimit[14]), .O(n28874));
    defparam i14803_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 LessThan_10_i9_2_lut (.I0(IntegralLimit[4]), .I1(n130[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5363));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i11_2_lut (.I0(IntegralLimit[5]), .I1(n130[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5364));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i13_2_lut (.I0(IntegralLimit[6]), .I1(n130[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5365));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28935_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[19]), .I2(n4_adj_5366), 
            .I3(n19484[1]), .O(n6_adj_4908));   // verilog/motorControl.v(52[18:24])
    defparam i28935_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_16_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_5090));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i15_2_lut (.I0(IntegralLimit[7]), .I1(n130[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5367));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i21_2_lut (.I0(IntegralLimit[10]), .I1(n130[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5368));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i9_2_lut (.I0(n130[4]), .I1(n182[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5369));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14808_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28878), 
            .I3(PWMLimit[13]), .O(n28879));
    defparam i14808_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 LessThan_12_i11_2_lut (.I0(n130[5]), .I1(n182[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5370));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i13_2_lut (.I0(n130[6]), .I1(n182[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5371));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14813_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28883), 
            .I3(PWMLimit[12]), .O(n28884));
    defparam i14813_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 LessThan_12_i15_2_lut (.I0(n130[7]), .I1(n182[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5372));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i21_2_lut (.I0(n130[10]), .I1(n182[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5373));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14818_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28888), 
            .I3(PWMLimit[11]), .O(n28889));
    defparam i14818_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_4_lut_adj_1717 (.I0(\Kp[3] ), .I1(n1[19]), .I2(n19484[1]), 
            .I3(n4_adj_5366), .O(n19453[2]));   // verilog/motorControl.v(52[18:24])
    defparam i1_3_lut_4_lut_adj_1717.LUT_INIT = 16'h8778;
    SB_LUT4 i14823_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28893), 
            .I3(PWMLimit[10]), .O(n28894));
    defparam i14823_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut_4_lut_adj_1718 (.I0(n62_adj_4891), .I1(n131_adj_4890), 
            .I2(n204_adj_4880), .I3(n19484[0]), .O(n19453[1]));   // verilog/motorControl.v(52[18:24])
    defparam i1_3_lut_4_lut_adj_1718.LUT_INIT = 16'h8778;
    SB_LUT4 mult_17_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_5304));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14828_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28898), 
            .I3(PWMLimit[9]), .O(n28899));
    defparam i14828_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14833_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28903), 
            .I3(PWMLimit[8]), .O(n28904));
    defparam i14833_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14838_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28908), 
            .I3(PWMLimit[7]), .O(n28909));
    defparam i14838_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14843_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28913), 
            .I3(PWMLimit[6]), .O(n28914));
    defparam i14843_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_17_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_5303));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38738_2_lut_4_lut (.I0(deadband[21]), .I1(n356[21]), .I2(deadband[9]), 
            .I3(n356[9]), .O(n54531));
    defparam i38738_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i14848_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28918), 
            .I3(PWMLimit[5]), .O(n28919));
    defparam i14848_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14853_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28923), 
            .I3(PWMLimit[4]), .O(n28924));
    defparam i14853_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i28927_3_lut_4_lut (.I0(n62_adj_4891), .I1(n131_adj_4890), .I2(n204_adj_4880), 
            .I3(n19484[0]), .O(n4_adj_5366));   // verilog/motorControl.v(52[18:24])
    defparam i28927_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i14858_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28928), 
            .I3(PWMLimit[3]), .O(n28929));
    defparam i14858_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_17_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i16_3_lut (.I0(n130[15]), .I1(n182[15]), .I2(n181), 
            .I3(GND_net), .O(n207[15]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_5302));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i16_3_lut (.I0(n207[15]), .I1(IntegralLimit[15]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [15]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14863_3_lut_4_lut (.I0(control_update), .I1(n409), .I2(n28933), 
            .I3(PWMLimit[2]), .O(n28934));
    defparam i14863_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mult_16_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_5301));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_5300));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i39_2_lut (.I0(IntegralLimit[19]), .I1(n130[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5374));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i41_2_lut (.I0(IntegralLimit[20]), .I1(n130[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5375));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i37_2_lut (.I0(IntegralLimit[18]), .I1(n130[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5376));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i35_2_lut (.I0(IntegralLimit[17]), .I1(n130[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5377));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i31_2_lut (.I0(IntegralLimit[15]), .I1(n130[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5378));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i33_2_lut (.I0(IntegralLimit[16]), .I1(n130[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5379));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i27_2_lut (.I0(IntegralLimit[13]), .I1(n130[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5380));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i29_2_lut (.I0(IntegralLimit[14]), .I1(n130[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5381));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i45_2_lut (.I0(IntegralLimit[22]), .I1(n130[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5382));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i25_2_lut (.I0(IntegralLimit[12]), .I1(n130[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5383));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_5299));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i23_2_lut (.I0(IntegralLimit[11]), .I1(n130[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5384));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i17_2_lut (.I0(IntegralLimit[8]), .I1(n130[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5385));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i19_2_lut (.I0(IntegralLimit[9]), .I1(n130[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5386));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i43_2_lut (.I0(IntegralLimit[21]), .I1(n130[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5387));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_5298));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38837_4_lut (.I0(n21_adj_5368), .I1(n19_adj_5386), .I2(n17_adj_5385), 
            .I3(n9_adj_5363), .O(n54630));
    defparam i38837_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i38830_4_lut (.I0(n27_adj_5380), .I1(n15_adj_5367), .I2(n13_adj_5365), 
            .I3(n11_adj_5364), .O(n54623));
    defparam i38830_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_10_i12_3_lut (.I0(n130[7]), .I1(n130[16]), .I2(n33_adj_5379), 
            .I3(GND_net), .O(n12_adj_5388));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i10_3_lut (.I0(n130[5]), .I1(n130[6]), .I2(n13_adj_5365), 
            .I3(GND_net), .O(n10_adj_5389));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i30_3_lut (.I0(n12_adj_5388), .I1(n130[17]), .I2(n35_adj_5377), 
            .I3(GND_net), .O(n30_adj_5390));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39234_4_lut (.I0(n13_adj_5365), .I1(n11_adj_5364), .I2(n9_adj_5363), 
            .I3(n54640), .O(n55027));
    defparam i39234_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39230_4_lut (.I0(n19_adj_5386), .I1(n17_adj_5385), .I2(n15_adj_5367), 
            .I3(n55027), .O(n55023));
    defparam i39230_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_17_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_5359));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39653_4_lut (.I0(n25_adj_5383), .I1(n23_adj_5384), .I2(n21_adj_5368), 
            .I3(n55023), .O(n55446));
    defparam i39653_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39424_4_lut (.I0(n31_adj_5378), .I1(n29_adj_5381), .I2(n27_adj_5380), 
            .I3(n55446), .O(n55217));
    defparam i39424_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39703_4_lut (.I0(n37_adj_5376), .I1(n35_adj_5377), .I2(n33_adj_5379), 
            .I3(n55217), .O(n55496));
    defparam i39703_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_10_i16_3_lut (.I0(n130[9]), .I1(n130[21]), .I2(n43_adj_5387), 
            .I3(GND_net), .O(n16_adj_5391));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39523_3_lut (.I0(n6_adj_5354), .I1(n130[10]), .I2(n21_adj_5368), 
            .I3(GND_net), .O(n55316));   // verilog/motorControl.v(47[12:34])
    defparam i39523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39524_3_lut (.I0(n55316), .I1(n130[11]), .I2(n23_adj_5384), 
            .I3(GND_net), .O(n55317));   // verilog/motorControl.v(47[12:34])
    defparam i39524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_5297));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i8_3_lut (.I0(n130[4]), .I1(n130[8]), .I2(n17_adj_5385), 
            .I3(GND_net), .O(n8_adj_5392));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i24_3_lut (.I0(n16_adj_5391), .I1(n130[22]), .I2(n45_adj_5382), 
            .I3(GND_net), .O(n24_adj_5393));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38816_4_lut (.I0(n43_adj_5387), .I1(n25_adj_5383), .I2(n23_adj_5384), 
            .I3(n54630), .O(n54609));
    defparam i38816_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39346_4_lut (.I0(n24_adj_5393), .I1(n8_adj_5392), .I2(n45_adj_5382), 
            .I3(n54607), .O(n55139));   // verilog/motorControl.v(47[12:34])
    defparam i39346_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39035_3_lut (.I0(n55317), .I1(n130[12]), .I2(n25_adj_5383), 
            .I3(GND_net), .O(n54828));   // verilog/motorControl.v(47[12:34])
    defparam i39035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i4_4_lut (.I0(n130[0]), .I1(n130[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_5394));   // verilog/motorControl.v(47[12:34])
    defparam LessThan_10_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i39521_3_lut (.I0(n4_adj_5394), .I1(n130[13]), .I2(n27_adj_5380), 
            .I3(GND_net), .O(n55314));   // verilog/motorControl.v(47[12:34])
    defparam i39521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39522_3_lut (.I0(n55314), .I1(n130[14]), .I2(n29_adj_5381), 
            .I3(GND_net), .O(n55315));   // verilog/motorControl.v(47[12:34])
    defparam i39522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38826_4_lut (.I0(n33_adj_5379), .I1(n31_adj_5378), .I2(n29_adj_5381), 
            .I3(n54623), .O(n54619));
    defparam i38826_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39665_4_lut (.I0(n30_adj_5390), .I1(n10_adj_5389), .I2(n35_adj_5377), 
            .I3(n54617), .O(n55458));   // verilog/motorControl.v(47[12:34])
    defparam i39665_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39037_3_lut (.I0(n55315), .I1(n130[15]), .I2(n31_adj_5378), 
            .I3(GND_net), .O(n54830));   // verilog/motorControl.v(47[12:34])
    defparam i39037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39749_4_lut (.I0(n54830), .I1(n55458), .I2(n35_adj_5377), 
            .I3(n54619), .O(n55542));   // verilog/motorControl.v(47[12:34])
    defparam i39749_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39750_3_lut (.I0(n55542), .I1(n130[18]), .I2(n37_adj_5376), 
            .I3(GND_net), .O(n55543));   // verilog/motorControl.v(47[12:34])
    defparam i39750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39734_3_lut (.I0(n55543), .I1(n130[19]), .I2(n39_adj_5374), 
            .I3(GND_net), .O(n55527));   // verilog/motorControl.v(47[12:34])
    defparam i39734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38818_4_lut (.I0(n43_adj_5387), .I1(n41_adj_5375), .I2(n39_adj_5374), 
            .I3(n55496), .O(n54611));
    defparam i38818_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39599_4_lut (.I0(n54828), .I1(n55139), .I2(n45_adj_5382), 
            .I3(n54609), .O(n55392));   // verilog/motorControl.v(47[12:34])
    defparam i39599_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_5296));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_5358));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39043_3_lut (.I0(n55527), .I1(n130[20]), .I2(n41_adj_5375), 
            .I3(GND_net), .O(n54836));   // verilog/motorControl.v(47[12:34])
    defparam i39043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39689_4_lut (.I0(n54836), .I1(n55392), .I2(n45_adj_5382), 
            .I3(n54611), .O(n55482));   // verilog/motorControl.v(47[12:34])
    defparam i39689_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39690_3_lut (.I0(n55482), .I1(IntegralLimit[23]), .I2(n130[23]), 
            .I3(GND_net), .O(n155));   // verilog/motorControl.v(47[12:34])
    defparam i39690_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_12_i41_2_lut (.I0(n130[20]), .I1(n182[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5395));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i37_2_lut (.I0(n130[18]), .I1(n182[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5396));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i39_2_lut (.I0(n130[19]), .I1(n182[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5397));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_5357));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i35_2_lut (.I0(n130[17]), .I1(n182[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5398));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i19_2_lut (.I0(n130[9]), .I1(n182[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5399));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i31_2_lut (.I0(n130[15]), .I1(n182[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5400));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i33_2_lut (.I0(n130[16]), .I1(n182[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5401));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_5295));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i29_2_lut (.I0(n130[14]), .I1(n182[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5402));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i27_2_lut (.I0(n130[13]), .I1(n182[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5403));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i23_2_lut (.I0(n130[11]), .I1(n182[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5404));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i25_2_lut (.I0(n130[12]), .I1(n182[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5405));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i43_2_lut (.I0(n130[21]), .I1(n182[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5406));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i45_2_lut (.I0(n130[22]), .I1(n182[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5407));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_5294));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i17_2_lut (.I0(n130[8]), .I1(n182[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5408));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38802_4_lut (.I0(n21_adj_5373), .I1(n19_adj_5399), .I2(n17_adj_5408), 
            .I3(n9_adj_5369), .O(n54595));
    defparam i38802_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28945_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [22]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [21]), .I3(\Ki[1] ), 
            .O(n19493[0]));   // verilog/motorControl.v(52[27:38])
    defparam i28945_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i38796_4_lut (.I0(n27_adj_5403), .I1(n15_adj_5372), .I2(n13_adj_5371), 
            .I3(n11_adj_5370), .O(n54589));
    defparam i38796_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_12_i12_3_lut (.I0(n182[7]), .I1(n182[16]), .I2(n33_adj_5401), 
            .I3(GND_net), .O(n12_adj_5409));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i10_3_lut (.I0(n182[5]), .I1(n182[6]), .I2(n13_adj_5371), 
            .I3(GND_net), .O(n10_adj_5410));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i30_3_lut (.I0(n12_adj_5409), .I1(n182[17]), .I2(n35_adj_5398), 
            .I3(GND_net), .O(n30_adj_5411));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39198_4_lut (.I0(n13_adj_5371), .I1(n11_adj_5370), .I2(n9_adj_5369), 
            .I3(n54605), .O(n54991));
    defparam i39198_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39194_4_lut (.I0(n19_adj_5399), .I1(n17_adj_5408), .I2(n15_adj_5372), 
            .I3(n54991), .O(n54987));
    defparam i39194_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39647_4_lut (.I0(n25_adj_5405), .I1(n23_adj_5404), .I2(n21_adj_5373), 
            .I3(n54987), .O(n55440));
    defparam i39647_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39408_4_lut (.I0(n31_adj_5400), .I1(n29_adj_5402), .I2(n27_adj_5403), 
            .I3(n55440), .O(n55201));
    defparam i39408_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39701_4_lut (.I0(n37_adj_5396), .I1(n35_adj_5398), .I2(n33_adj_5401), 
            .I3(n55201), .O(n55494));
    defparam i39701_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_12_i16_3_lut (.I0(n182[9]), .I1(n182[21]), .I2(n43_adj_5406), 
            .I3(GND_net), .O(n16_adj_5412));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_5293));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39515_3_lut (.I0(n6_adj_5351), .I1(n182[10]), .I2(n21_adj_5373), 
            .I3(GND_net), .O(n55308));   // verilog/motorControl.v(49[21:44])
    defparam i39515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39516_3_lut (.I0(n55308), .I1(n182[11]), .I2(n23_adj_5404), 
            .I3(GND_net), .O(n55309));   // verilog/motorControl.v(49[21:44])
    defparam i39516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_5292));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_5291));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i8_3_lut (.I0(n182[4]), .I1(n182[8]), .I2(n17_adj_5408), 
            .I3(GND_net), .O(n8_adj_5413));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i24_3_lut (.I0(n16_adj_5412), .I1(n182[22]), .I2(n45_adj_5407), 
            .I3(GND_net), .O(n24_adj_5414));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38782_4_lut (.I0(n43_adj_5406), .I1(n25_adj_5405), .I2(n23_adj_5404), 
            .I3(n54595), .O(n54575));
    defparam i38782_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39348_4_lut (.I0(n24_adj_5414), .I1(n8_adj_5413), .I2(n45_adj_5407), 
            .I3(n54573), .O(n55141));   // verilog/motorControl.v(49[21:44])
    defparam i39348_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39045_3_lut (.I0(n55309), .I1(n182[12]), .I2(n25_adj_5405), 
            .I3(GND_net), .O(n54838));   // verilog/motorControl.v(49[21:44])
    defparam i39045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i4_4_lut (.I0(n130[0]), .I1(n182[1]), .I2(n130[1]), 
            .I3(n182[0]), .O(n4_adj_5415));   // verilog/motorControl.v(49[21:44])
    defparam LessThan_12_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_17_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_5290));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39513_3_lut (.I0(n4_adj_5415), .I1(n182[13]), .I2(n27_adj_5403), 
            .I3(GND_net), .O(n55306));   // verilog/motorControl.v(49[21:44])
    defparam i39513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39514_3_lut (.I0(n55306), .I1(n182[14]), .I2(n29_adj_5402), 
            .I3(GND_net), .O(n55307));   // verilog/motorControl.v(49[21:44])
    defparam i39514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38792_4_lut (.I0(n33_adj_5401), .I1(n31_adj_5400), .I2(n29_adj_5402), 
            .I3(n54589), .O(n54585));
    defparam i38792_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_5356));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39667_4_lut (.I0(n30_adj_5411), .I1(n10_adj_5410), .I2(n35_adj_5398), 
            .I3(n54583), .O(n55460));   // verilog/motorControl.v(49[21:44])
    defparam i39667_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_17_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_5289));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_5355));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_5288));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39047_3_lut (.I0(n55307), .I1(n182[15]), .I2(n31_adj_5400), 
            .I3(GND_net), .O(n54840));   // verilog/motorControl.v(49[21:44])
    defparam i39047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_5086));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39751_4_lut (.I0(n54840), .I1(n55460), .I2(n35_adj_5398), 
            .I3(n54585), .O(n55544));   // verilog/motorControl.v(49[21:44])
    defparam i39751_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39752_3_lut (.I0(n55544), .I1(n182[18]), .I2(n37_adj_5396), 
            .I3(GND_net), .O(n55545));   // verilog/motorControl.v(49[21:44])
    defparam i39752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28947_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [22]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [21]), .I3(\Ki[1] ), 
            .O(n43024));   // verilog/motorControl.v(52[27:38])
    defparam i28947_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i39730_3_lut (.I0(n55545), .I1(n182[19]), .I2(n39_adj_5397), 
            .I3(GND_net), .O(n55523));   // verilog/motorControl.v(49[21:44])
    defparam i39730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38784_4_lut (.I0(n43_adj_5406), .I1(n41_adj_5395), .I2(n39_adj_5397), 
            .I3(n55494), .O(n54577));
    defparam i38784_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39601_4_lut (.I0(n54838), .I1(n55141), .I2(n45_adj_5407), 
            .I3(n54575), .O(n55394));   // verilog/motorControl.v(49[21:44])
    defparam i39601_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39053_3_lut (.I0(n55523), .I1(n182[20]), .I2(n41_adj_5395), 
            .I3(GND_net), .O(n54846));   // verilog/motorControl.v(49[21:44])
    defparam i39053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39691_4_lut (.I0(n54846), .I1(n55394), .I2(n45_adj_5407), 
            .I3(n54577), .O(n55484));   // verilog/motorControl.v(49[21:44])
    defparam i39691_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39692_3_lut (.I0(n55484), .I1(n130[23]), .I2(n182[23]), .I3(GND_net), 
            .O(n181));   // verilog/motorControl.v(49[21:44])
    defparam i39692_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_14_i2_3_lut (.I0(n130[1]), .I1(n182[1]), .I2(n181), .I3(GND_net), 
            .O(n207[1]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i2_3_lut (.I0(n207[1]), .I1(IntegralLimit[1]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [1]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_5287));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28851_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n42908), .I3(n201_adj_5362), 
            .O(n4_adj_5348));   // verilog/motorControl.v(52[27:38])
    defparam i28851_3_lut_4_lut.LUT_INIT = 16'hf660;
    SB_LUT4 i28762_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [20]), .I3(\Ki[1] ), 
            .O(n19469[0]));   // verilog/motorControl.v(52[27:38])
    defparam i28762_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i28764_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3996 [20]), .I3(\Ki[1] ), 
            .O(n42826));   // verilog/motorControl.v(52[27:38])
    defparam i28764_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_5286));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_5285));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_5283));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38559_2_lut_4_lut (.I0(n356[21]), .I1(n436[21]), .I2(n356[9]), 
            .I3(n436[9]), .O(n54351));
    defparam i38559_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_5282));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38573_2_lut_4_lut (.I0(n356[16]), .I1(n436[16]), .I2(n356[7]), 
            .I3(n436[7]), .O(n54365));
    defparam i38573_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i38607_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(PWMLimit[9]), 
            .I3(n356[9]), .O(n54400));
    defparam i38607_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_5281));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_5280));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28821_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(n4_adj_4966), .I3(n19469[1]), .O(n6_adj_4884));   // verilog/motorControl.v(52[27:38])
    defparam i28821_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_16_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i7_3_lut (.I0(n130[6]), .I1(n182[6]), .I2(n181), .I3(GND_net), 
            .O(n207[6]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i7_3_lut (.I0(n207[6]), .I1(IntegralLimit[6]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [6]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_5279));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_5278));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_5056));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5055));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_5051));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_5277));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_5047));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_5276));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_5046));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1719 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [19]), 
            .I2(n4_adj_4966), .I3(n19469[1]), .O(n19429[2]));   // verilog/motorControl.v(52[27:38])
    defparam i1_3_lut_4_lut_adj_1719.LUT_INIT = 16'h8778;
    SB_LUT4 mult_17_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_5275));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38633_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(PWMLimit[7]), 
            .I3(n356[7]), .O(n54426));
    defparam i38633_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_5039));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_5274));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_5018));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_5273));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_5272));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_5271));   // verilog/motorControl.v(52[18:24])
    defparam mult_16_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_5270));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n19429[2]), .I1(n6_adj_4882), .I2(\Ki[4] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3996 [18]), .O(n19369[3]));   // verilog/motorControl.v(52[27:38])
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'h9666;
    SB_LUT4 mult_17_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_5353));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i18_3_lut (.I0(n130[17]), .I1(n182[17]), .I2(n181), 
            .I3(GND_net), .O(n207[17]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_14_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28914_2_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(\Kp[1] ), 
            .I3(n1[19]), .O(n19453[0]));   // verilog/motorControl.v(52[18:24])
    defparam i28914_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mux_15_i18_3_lut (.I0(n207[17]), .I1(IntegralLimit[17]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3996 [17]));   // verilog/motorControl.v(49[18] 51[12])
    defparam mux_15_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_5002));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_5352));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i136_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n201_adj_5362));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3996 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_5001));   // verilog/motorControl.v(52[27:38])
    defparam mult_17_i36_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (clk16MHz, \state[3] , n6, GND_net, read, \state[0] , 
            enable_slow_N_4393, n6271, \state[1] , n48226, VCC_net, 
            n36101, n49533, n49611, n48264, n29303, rw, n48368, 
            data_ready, n7354, \state[2] , \state_7__N_4290[0] , n4, 
            n4_adj_19, n35819, scl_enable, n26, \state_7__N_4306[3] , 
            n7936, sda_enable, n29357, \saved_addr[0] , \state[0]_adj_20 , 
            n29269, data, n29268, n29267, n29266, n29265, n29264, 
            n29263, n10, n10_adj_21, n8, n29727, n54311, n27267, 
            n27262, scl, sda_out) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    output \state[3] ;
    output n6;
    input GND_net;
    input read;
    output \state[0] ;
    output enable_slow_N_4393;
    output [0:0]n6271;
    output \state[1] ;
    input n48226;
    input VCC_net;
    output n36101;
    input n49533;
    output n49611;
    input n48264;
    input n29303;
    output rw;
    input n48368;
    output data_ready;
    output n7354;
    output \state[2] ;
    output \state_7__N_4290[0] ;
    output n4;
    output n4_adj_19;
    output n35819;
    output scl_enable;
    output n26;
    input \state_7__N_4306[3] ;
    input n7936;
    output sda_enable;
    input n29357;
    output \saved_addr[0] ;
    output \state[0]_adj_20 ;
    input n29269;
    output [7:0]data;
    input n29268;
    input n29267;
    input n29266;
    input n29265;
    input n29264;
    input n29263;
    output n10;
    output n10_adj_21;
    input n8;
    input n29727;
    output n54311;
    output n27267;
    output n27262;
    output scl;
    output sda_out;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [15:0]delay_counter_15__N_4192;
    
    wire n28826;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    
    wire n29219, n27130, n28, n26_c, n27, n25, enable;
    wire [15:0]n4876;
    
    wire n43355, n43354, n43353, n43352, n43351, n43350, n43349, 
        n43348, n43347, n43346, n43345, n43344, n43343, n43342, 
        n43341;
    
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[1]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[2]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[3]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[4]), .S(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[5]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[6]), .S(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[7]), .S(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[8]), .S(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[9]), .S(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i2_2_lut (.I0(\state[3] ), .I1(n27130), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26_c));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26_c), .I3(n28), .O(n27130));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1487_Mux_0_i1_4_lut (.I0(read), .I1(n27130), .I2(\state[0] ), 
            .I3(enable_slow_N_4393), .O(n6271[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_1487_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n28826), .D(delay_counter_15__N_4192[10]), .S(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n28826), .D(delay_counter_15__N_4192[11]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFSR enable_39 (.Q(enable), .C(clk16MHz), .D(n6271[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n28826), .D(delay_counter_15__N_4192[12]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n28826), .D(delay_counter_15__N_4192[13]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n28826), .D(delay_counter_15__N_4192[14]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n28826), .D(delay_counter_15__N_4192[15]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFE state__i1 (.Q(\state[1] ), .C(clk16MHz), .E(VCC_net), .D(n48226));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i15156_2_lut (.I0(n28826), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29219));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15156_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n28826));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i22041_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_4393), 
            .I3(GND_net), .O(n36101));   // verilog/eeprom.v(51[5:9])
    defparam i22041_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i33876_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n49533), 
            .I3(enable_slow_N_4393), .O(n49611));   // verilog/eeprom.v(51[5:9])
    defparam i33876_4_lut_4_lut.LUT_INIT = 16'hfcf8;
    SB_LUT4 i39795_2_lut (.I0(n27130), .I1(enable_slow_N_4393), .I2(GND_net), 
            .I3(GND_net), .O(n4876[4]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i39795_2_lut.LUT_INIT = 16'h2222;
    SB_DFF state__i0 (.Q(\state[0] ), .C(clk16MHz), .D(n48264));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n28826), 
            .D(delay_counter_15__N_4192[0]), .R(n29219));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF rw_43 (.Q(rw), .C(clk16MHz), .D(n29303));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(clk16MHz), .D(n48368));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_1035_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n4876[4]), 
            .I3(n43355), .O(delay_counter_15__N_4192[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1035_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n4876[4]), 
            .I3(n43354), .O(delay_counter_15__N_4192[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_16 (.CI(n43354), .I0(delay_counter[14]), .I1(n4876[4]), 
            .CO(n43355));
    SB_LUT4 add_1035_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n4876[4]), 
            .I3(n43353), .O(delay_counter_15__N_4192[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_15 (.CI(n43353), .I0(delay_counter[13]), .I1(n4876[4]), 
            .CO(n43354));
    SB_LUT4 add_1035_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n4876[4]), 
            .I3(n43352), .O(delay_counter_15__N_4192[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_14 (.CI(n43352), .I0(delay_counter[12]), .I1(n4876[4]), 
            .CO(n43353));
    SB_LUT4 add_1035_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n4876[4]), 
            .I3(n43351), .O(delay_counter_15__N_4192[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_13 (.CI(n43351), .I0(delay_counter[11]), .I1(n4876[4]), 
            .CO(n43352));
    SB_LUT4 add_1035_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n4876[4]), 
            .I3(n43350), .O(delay_counter_15__N_4192[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_12 (.CI(n43350), .I0(delay_counter[10]), .I1(n4876[4]), 
            .CO(n43351));
    SB_LUT4 add_1035_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n4876[4]), 
            .I3(n43349), .O(delay_counter_15__N_4192[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_11 (.CI(n43349), .I0(delay_counter[9]), .I1(n4876[4]), 
            .CO(n43350));
    SB_LUT4 add_1035_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n4876[4]), 
            .I3(n43348), .O(delay_counter_15__N_4192[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_10 (.CI(n43348), .I0(delay_counter[8]), .I1(n4876[4]), 
            .CO(n43349));
    SB_LUT4 add_1035_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n4876[4]), 
            .I3(n43347), .O(delay_counter_15__N_4192[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_9 (.CI(n43347), .I0(delay_counter[7]), .I1(n4876[4]), 
            .CO(n43348));
    SB_LUT4 add_1035_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n4876[4]), 
            .I3(n43346), .O(delay_counter_15__N_4192[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_8 (.CI(n43346), .I0(delay_counter[6]), .I1(n4876[4]), 
            .CO(n43347));
    SB_LUT4 add_1035_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n4876[4]), 
            .I3(n43345), .O(delay_counter_15__N_4192[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_7 (.CI(n43345), .I0(delay_counter[5]), .I1(n4876[4]), 
            .CO(n43346));
    SB_LUT4 add_1035_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n4876[4]), 
            .I3(n43344), .O(delay_counter_15__N_4192[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_6 (.CI(n43344), .I0(delay_counter[4]), .I1(n4876[4]), 
            .CO(n43345));
    SB_LUT4 add_1035_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n4876[4]), 
            .I3(n43343), .O(delay_counter_15__N_4192[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_5 (.CI(n43343), .I0(delay_counter[3]), .I1(n4876[4]), 
            .CO(n43344));
    SB_LUT4 add_1035_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n4876[4]), 
            .I3(n43342), .O(delay_counter_15__N_4192[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_4 (.CI(n43342), .I0(delay_counter[2]), .I1(n4876[4]), 
            .CO(n43343));
    SB_LUT4 add_1035_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n4876[4]), 
            .I3(n43341), .O(delay_counter_15__N_4192[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_3 (.CI(n43341), .I0(delay_counter[1]), .I1(n4876[4]), 
            .CO(n43342));
    SB_LUT4 add_1035_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n4876[4]), 
            .I3(GND_net), .O(delay_counter_15__N_4192[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1035_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1035_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n4876[4]), 
            .CO(n43341));
    i2c_controller i2c (.n7354(n7354), .\state[2] (\state[2] ), .\state_7__N_4290[0] (\state_7__N_4290[0] ), 
            .enable_slow_N_4393(enable_slow_N_4393), .GND_net(GND_net), 
            .\state[3] (\state[3] ), .n4(n4), .n4_adj_17(n4_adj_19), .n35819(n35819), 
            .clk16MHz(clk16MHz), .scl_enable(scl_enable), .n26(n26), .\state_7__N_4306[3] (\state_7__N_4306[3] ), 
            .n7936(n7936), .sda_enable(sda_enable), .n29357(n29357), .\saved_addr[0] (\saved_addr[0] ), 
            .VCC_net(VCC_net), .\state[0] (\state[0]_adj_20 ), .n29269(n29269), 
            .data({data}), .n29268(n29268), .n29267(n29267), .n29266(n29266), 
            .n29265(n29265), .n29264(n29264), .n29263(n29263), .n10(n10), 
            .enable(enable), .n10_adj_18(n10_adj_21), .n8(n8), .n29727(n29727), 
            .n54311(n54311), .n27267(n27267), .n27262(n27262), .scl(scl), 
            .sda_out(sda_out)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (n7354, \state[2] , \state_7__N_4290[0] , enable_slow_N_4393, 
            GND_net, \state[3] , n4, n4_adj_17, n35819, clk16MHz, 
            scl_enable, n26, \state_7__N_4306[3] , n7936, sda_enable, 
            n29357, \saved_addr[0] , VCC_net, \state[0] , n29269, 
            data, n29268, n29267, n29266, n29265, n29264, n29263, 
            n10, enable, n10_adj_18, n8, n29727, n54311, n27267, 
            n27262, scl, sda_out) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output n7354;
    output \state[2] ;
    output \state_7__N_4290[0] ;
    output enable_slow_N_4393;
    input GND_net;
    output \state[3] ;
    output n4;
    output n4_adj_17;
    output n35819;
    input clk16MHz;
    output scl_enable;
    output n26;
    input \state_7__N_4306[3] ;
    input n7936;
    output sda_enable;
    input n29357;
    output \saved_addr[0] ;
    input VCC_net;
    output \state[0] ;
    input n29269;
    output [7:0]data;
    input n29268;
    input n29267;
    input n29266;
    input n29265;
    input n29264;
    input n29263;
    output n10;
    input enable;
    output n10_adj_18;
    input n8;
    input n29727;
    output n54311;
    output n27267;
    output n27262;
    output scl;
    output sda_out;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n5;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n36572, n35999, n36031, enable_slow_N_4392, n48426, n50642;
    wire [7:0]n119;
    
    wire n28748;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n29132;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n10_c, n29081, i2c_clk_N_4379, scl_enable_N_4380, n15, n49539, 
        n7347, n37, n28691;
    wire [5:0]n29;
    
    wire n19511, n7849, n29075, n43507, n43506, n43505, n43504, 
        n43503, n43502, n43501;
    wire [0:0]n7051;
    
    wire n29072, sda_out_adj_4864, n54255, n54227, n7050, n7, n10_adj_4865, 
        n54319, n11, n12, n34_adj_4868, n33_adj_4869, n9, state_7__N_4289, 
        n11_adj_4870, n36403, n11_adj_4871, n44208, n44207, n44206, 
        n44205, n44204, n11_adj_4872, n4_adj_4873;
    
    SB_DFFESS state_i0_i1 (.Q(state[1]), .C(i2c_clk), .E(n7354), .D(n5), 
            .S(n36572));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n7354), .D(n35999), 
            .S(n36031));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i39826_2_lut (.I0(\state_7__N_4290[0] ), .I1(enable_slow_N_4393), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4392));   // verilog/i2c_controller.v(62[6:32])
    defparam i39826_2_lut.LUT_INIT = 16'h7777;
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n7354), .D(n48426), 
            .S(n50642));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n28748), .D(n119[1]), 
            .S(n29132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n28748), .D(n119[2]), 
            .S(n29132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n28748), .D(n119[3]), 
            .R(n29132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n28748), .D(n119[4]), 
            .R(n29132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n28748), .D(n119[5]), 
            .R(n29132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n28748), .D(n119[6]), 
            .R(n29132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n28748), .D(n119[7]), 
            .R(n29132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 equal_385_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_385_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_383_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_17));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_383_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n29081));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i21759_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35819));
    defparam i21759_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n29081), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4379));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4379));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4380));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 i1_2_lut_adj_1693 (.I0(\state[2] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n26));
    defparam i1_2_lut_adj_1693.LUT_INIT = 16'heeee;
    SB_LUT4 i33809_2_lut (.I0(\state_7__N_4306[3] ), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n49539));
    defparam i33809_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(n7347), .I1(n49539), .I2(n7936), .I3(n37), 
            .O(n28748));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_DFFE enable_slow_120 (.Q(\state_7__N_4290[0] ), .C(clk16MHz), .E(n28691), 
            .D(enable_slow_N_4392));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFSR counter2_2294_2295__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n29081));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n7849), 
            .D(n19511), .S(n29075));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFSR counter2_2294_2295__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n29081));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2294_2295__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n29081));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2294_2295__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n29081));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2294_2295__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n29081));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29357));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n43507), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n43506), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n43506), .I0(counter[6]), .I1(VCC_net), 
            .CO(n43507));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n43505), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n43505), .I0(counter[5]), .I1(VCC_net), 
            .CO(n43506));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n43504), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n43504), .I0(counter[4]), .I1(VCC_net), 
            .CO(n43505));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n43503), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n43503), .I0(counter[3]), .I1(VCC_net), 
            .CO(n43504));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n43502), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n43502), .I0(counter[2]), .I1(VCC_net), 
            .CO(n43503));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n43501), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n43501), .I0(counter[1]), .I1(VCC_net), 
            .CO(n43502));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n43501));
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4864), .C(i2c_clk), .E(n29072), 
            .D(n7051[0]));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n28748), .D(n119[0]), 
            .S(n29132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i38616_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n54255));   // verilog/i2c_controller.v(198[28:35])
    defparam i38616_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i38583_4_lut (.I0(n54255), .I1(state[1]), .I2(counter[0]), 
            .I3(counter[2]), .O(n54227));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i38583_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 mux_1682_i1_4_lut (.I0(n54227), .I1(\state[0] ), .I2(n7050), 
            .I3(\state[2] ), .O(n7051[0]));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam mux_1682_i1_4_lut.LUT_INIT = 16'h303a;
    SB_DFFSR counter2_2294_2295__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n29081));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29269));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29268));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29267));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29266));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29265));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29264));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29263));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_adj_1694 (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_1694.LUT_INIT = 16'h4444;
    SB_LUT4 i38626_4_lut (.I0(n10_adj_4865), .I1(n10), .I2(\state_7__N_4306[3] ), 
            .I3(enable), .O(n54319));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i38626_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut (.I0(state[1]), .I1(n7), .I2(n54319), .I3(\state[0] ), 
            .O(n48426));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i40426_2_lut (.I0(\state_7__N_4306[3] ), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n35999));
    defparam i40426_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_18));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10_adj_18), 
            .O(n7347));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[1]), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34_adj_4868));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33_adj_4869));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_LUT4 equal_309_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4865));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_309_i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i39806_4_lut (.I0(state_7__N_4289), .I1(n7347), .I2(n11_adj_4870), 
            .I3(n36403), .O(n7354));
    defparam i39806_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n11_adj_4871), .I1(n11), .I2(\state_7__N_4306[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'h5755;
    SB_LUT4 equal_2273_i19_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4393));   // verilog/i2c_controller.v(77[47:62])
    defparam equal_2273_i19_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n29727));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 counter2_2294_2295_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n44208), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2294_2295_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n44207), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2294_2295_add_4_6 (.CI(n44207), .I0(GND_net), .I1(counter2[4]), 
            .CO(n44208));
    SB_LUT4 counter2_2294_2295_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n44206), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2294_2295_add_4_5 (.CI(n44206), .I0(GND_net), .I1(counter2[3]), 
            .CO(n44207));
    SB_LUT4 counter2_2294_2295_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n44205), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2294_2295_add_4_4 (.CI(n44205), .I0(GND_net), .I1(counter2[2]), 
            .CO(n44206));
    SB_LUT4 counter2_2294_2295_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n44204), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2294_2295_add_4_3 (.CI(n44204), .I0(GND_net), .I1(counter2[1]), 
            .CO(n44205));
    SB_LUT4 counter2_2294_2295_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2294_2295_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2294_2295_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n44204));
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4871));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 equal_309_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_309_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i38685_3_lut_4_lut (.I0(n11_adj_4870), .I1(n11_adj_4872), .I2(enable_slow_N_4393), 
            .I3(\state_7__N_4290[0] ), .O(n54311));
    defparam i38685_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 i40433_3_lut_4_lut (.I0(n11_adj_4870), .I1(n11_adj_4872), .I2(n15), 
            .I3(n7354), .O(n36572));
    defparam i40433_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i22395_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_4289));
    defparam i22395_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11_adj_4872));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10), .I2(counter[0]), .I3(GND_net), 
            .O(n27267));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1696 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n27262));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_1696.LUT_INIT = 16'hfefe;
    SB_LUT4 i40431_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11_adj_4872), 
            .I3(n7354), .O(n36031));   // verilog/i2c_controller.v(151[5:14])
    defparam i40431_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4870));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i22342_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n36403));
    defparam i22342_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i40429_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(state[1]), 
            .I3(n7354), .O(n50642));
    defparam i40429_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[0] ), .I1(\state[3] ), .I2(state[1]), 
            .I3(\state[2] ), .O(n29072));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0316;
    SB_LUT4 i21755_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i21755_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2711_2_lut (.I0(sda_out_adj_4864), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2711_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22421_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[2] ), 
            .I3(n15), .O(scl_enable_N_4380));   // verilog/i2c_controller.v(77[47:62])
    defparam i22421_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_4_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[3] ), 
            .I3(\state[2] ), .O(n7050));   // verilog/i2c_controller.v(77[47:62])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h001a;
    SB_LUT4 i1_2_lut_adj_1697 (.I0(\state[2] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4873));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i1_2_lut_adj_1697.LUT_INIT = 16'h4444;
    SB_LUT4 i33779_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n49539), .O(n29132));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i33779_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_4_lut_adj_1698 (.I0(\state[3] ), .I1(\state[2] ), .I2(state[1]), 
            .I3(\state[0] ), .O(n37));
    defparam i1_4_lut_4_lut_adj_1698.LUT_INIT = 16'h1154;
    SB_LUT4 i1_3_lut (.I0(state[1]), .I1(n33_adj_4869), .I2(n37), .I3(GND_net), 
            .O(n29075));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i39840_4_lut (.I0(n7050), .I1(n34_adj_4868), .I2(n4_adj_4873), 
            .I3(n37), .O(n7849));
    defparam i39840_4_lut.LUT_INIT = 16'haf8c;
    SB_LUT4 i40423_2_lut (.I0(\state[0] ), .I1(n7050), .I2(GND_net), .I3(GND_net), 
            .O(n19511));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i40423_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_3_lut_adj_1699 (.I0(enable), .I1(\state_7__N_4290[0] ), 
            .I2(enable_slow_N_4393), .I3(GND_net), .O(n28691));
    defparam i1_2_lut_3_lut_adj_1699.LUT_INIT = 16'heaea;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n29426, deadband, clk16MHz, n29425, n29424, n29423, 
            n29422, GND_net, \data_in_frame[16] , rx_data, \data_in_frame[5] , 
            n29421, \data_in_frame[14] , \data_in_frame[12] , \data_in_frame[15] , 
            \data_out_frame[6] , \data_out_frame[7] , \data_in_frame[10] , 
            \data_out_frame[4] , \data_out_frame[5] , n4452, \FRAME_MATCHER.i_31__N_2845 , 
            n22902, \data_in_frame[3] , n29419, \data_in_frame[2] , 
            \data_in_frame[1] , \data_in_frame[21] , \data_out_frame[8] , 
            \data_out_frame[9] , \data_out_frame[10] , \data_out_frame[11] , 
            \data_out_frame[14] , \data_out_frame[15] , \data_out_frame[12] , 
            \data_out_frame[13] , \data_out_frame[16] , \data_out_frame[17] , 
            \data_out_frame[18] , \data_out_frame[19] , \data_out_frame[22] , 
            \data_out_frame[23] , \data_out_frame[20] , \data_out_frame[21] , 
            n29418, \data_in_frame[6] , n29417, \data_in_frame[4] , 
            \data_in_frame[9] , \data_in_frame[13] , \data_in[1] , \data_in[2] , 
            \data_in[3] , \data_in[0] , \data_in[1][1] , \data_in[2][5] , 
            \data_in[1][6] , \data_in[1][3] , \data_in[2][0] , \data_in[1][2] , 
            \data_in[2][6] , \data_in[2][3] , \data_in[3][3] , \data_in[3][5] , 
            \data_in[3][6] , \data_in[2][1] , rx_data_ready, n63, n3303, 
            n4599, n48672, n4, n48616, \data_in_frame[8] , n29416, 
            n29415, \Kp[2] , setpoint, ID, \data_in_frame[11] , n29411, 
            \Kp[3] , tx_active, \data_in_frame[20] , n29410, \Kp[4] , 
            \data_in_frame[23] , \FRAME_MATCHER.state[0] , n29409, \Kp[5] , 
            n29408, \Kp[6] , n29407, \Kp[7] , n29406, \Kp[8] , n29405, 
            \Kp[9] , n29404, \Kp[10] , n29403, \Kp[11] , n29402, 
            \Kp[12] , n29401, \Kp[13] , n29400, \Kp[14] , n29396, 
            \Kp[15] , n29395, \Ki[1] , n29394, \Ki[2] , n29391, 
            \Ki[3] , n29390, \Ki[4] , n29389, \Ki[5] , n29388, \Ki[6] , 
            n29387, \Ki[7] , n29386, \Ki[8] , n29385, \Ki[9] , n29384, 
            \Ki[10] , n29378, \Ki[11] , n29377, \Ki[12] , n29376, 
            \Ki[13] , n29375, \Ki[14] , \data_out_frame[25] , \data_out_frame[24] , 
            n29374, \Ki[15] , n29373, n29372, n29371, n29370, n29369, 
            n29368, n29366, n29365, n29364, n29363, n29362, n29361, 
            n29360, n29358, n29355, n29354, n29353, n29352, n29351, 
            n29349, n29347, n29346, n29345, n29343, n29341, n29340, 
            n29339, n29338, n29337, n29336, n29335, n29334, n29333, 
            n29332, n29331, n29330, n29329, n29328, n29327, n29326, 
            n29325, n29323, n29322, n50602, n122, \FRAME_MATCHER.i_31__N_2843 , 
            n5, n57092, n29321, n29957, n29956, n29955, n29954, 
            n29953, n29952, n29951, n29950, n29949, n29948, n29947, 
            n29946, n29945, n29944, n29943, n29942, n29941, n29940, 
            n29939, n29938, n29937, n29936, n29935, n29934, n29933, 
            n29932, n29931, n29930, n29929, n29928, n29927, n29926, 
            n29925, n29924, n29923, n29922, n29921, n29920, n29919, 
            n29918, n29917, n29916, n29915, n29914, n29913, n29912, 
            n29911, n29910, n29909, n29908, n29907, n29906, n29905, 
            n29904, n29903, n29902, n29901, n29900, n29899, n29898, 
            n29897, n29896, n29895, n29894, n29893, n29892, n29891, 
            n29890, n29889, n29888, n29887, n29886, n29885, n29884, 
            n29883, n29882, DE_c, LED_c, n29319, n29318, n29316, 
            n29315, n29314, n29313, n29312, n29311, n29310, n29307, 
            n29306, n29305, n29304, n29300, n29299, n29298, n29297, 
            n29296, n29881, n29880, n29879, n29878, n29877, n29876, 
            n29875, n29874, n29873, n29872, n29871, n29870, n29869, 
            n29868, n29867, n29859, n29858, n29857, n29856, n29855, 
            n29854, n29853, n29852, n29851, control_mode, n29295, 
            n29850, n29849, n29848, n29847, n29846, n29845, n29294, 
            n29844, current_limit, n29293, n29843, n29842, n29841, 
            n29840, n29292, n29291, n29290, n29288, n29287, n29286, 
            n48016, n29284, PWMLimit, n29283, n29282, n29280, neopxl_color, 
            n29279, n29278, \Ki[0] , n29277, \Kp[0] , n29276, IntegralLimit, 
            n29275, n29274, n29273, n29839, n29838, n29837, n29836, 
            n29835, n29834, n63_adj_6, n29833, n29832, n9, n29831, 
            n29830, n29829, n29828, n29260, n29259, n29827, n29826, 
            n29825, n29824, n29823, n29822, n29821, n29820, n29256, 
            n29819, n29818, n29817, n29816, n29815, n29814, n29813, 
            n29812, n29811, n29810, n29809, n29808, n29807, n56702, 
            n29762, n29761, n29760, n29759, n29758, n29757, n29756, 
            n29755, n29754, n29753, n29752, n29751, n29726, n29725, 
            n29724, n29723, n29722, n29721, n29720, n29719, n29718, 
            n29717, n29716, n29707, n29706, n29705, n29704, n29703, 
            n29702, n29701, n29687, n29686, n29685, n29666, n29665, 
            n29664, n29663, n29662, n29661, n29660, n29659, n29658, 
            n29657, n29656, n29655, n29654, n29653, n29652, n29651, 
            n29650, n29649, n29648, n29646, n29645, n29644, n29643, 
            n29483, n29482, n29481, n29480, n29479, n29478, n29477, 
            n29476, n29468, n29467, n29466, n29465, n29464, n29463, 
            n29462, n29461, n29460, n29459, n29458, n29457, n29456, 
            n29455, n29454, n29453, n29452, n29451, n29450, n29449, 
            n29448, n29447, n29446, n29445, \Kp[1] , n29442, n29441, 
            n29440, n29439, n29438, n29437, n29434, n29433, n29432, 
            n29431, n29430, n29429, n29428, n5_adj_7, n50620, n24373, 
            n48646, n48638, \state[0] , \state[2] , \state[3] , n7936, 
            n28758, n29184, \r_Bit_Index[0] , r_SM_Main, \r_SM_Main_2__N_3848[1] , 
            VCC_net, tx_o, n29324, n29732, n56700, n4_adj_8, tx_enable, 
            n19731, n28762, n29186, n29420, r_SM_Main_adj_16, r_Rx_Data, 
            \r_SM_Main_2__N_3777[2] , n35837, RX_N_10, n4_adj_12, n4_adj_13, 
            n29735, \r_Bit_Index[0]_adj_14 , n48270, n29261, n4_adj_15, 
            n29769, n29767, n29766, n48565, n29749, n29748, n29740, 
            n27227, n27232) /* synthesis syn_module_defined=1 */ ;
    input n29426;
    output [23:0]deadband;
    input clk16MHz;
    input n29425;
    input n29424;
    input n29423;
    input n29422;
    input GND_net;
    output [7:0]\data_in_frame[16] ;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[5] ;
    input n29421;
    output [7:0]\data_in_frame[14] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[15] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    output n4452;
    output \FRAME_MATCHER.i_31__N_2845 ;
    output n22902;
    output [7:0]\data_in_frame[3] ;
    input n29419;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[21] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[22] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[21] ;
    input n29418;
    output [7:0]\data_in_frame[6] ;
    input n29417;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[0] ;
    output \data_in[1][1] ;
    output \data_in[2][5] ;
    output \data_in[1][6] ;
    output \data_in[1][3] ;
    output \data_in[2][0] ;
    output \data_in[1][2] ;
    output \data_in[2][6] ;
    output \data_in[2][3] ;
    output \data_in[3][3] ;
    output \data_in[3][5] ;
    output \data_in[3][6] ;
    output \data_in[2][1] ;
    output rx_data_ready;
    output n63;
    output n3303;
    output n4599;
    output n48672;
    output n4;
    output n48616;
    output [7:0]\data_in_frame[8] ;
    input n29416;
    input n29415;
    output \Kp[2] ;
    output [23:0]setpoint;
    input [7:0]ID;
    output [7:0]\data_in_frame[11] ;
    input n29411;
    output \Kp[3] ;
    output tx_active;
    output [7:0]\data_in_frame[20] ;
    input n29410;
    output \Kp[4] ;
    output [7:0]\data_in_frame[23] ;
    output \FRAME_MATCHER.state[0] ;
    input n29409;
    output \Kp[5] ;
    input n29408;
    output \Kp[6] ;
    input n29407;
    output \Kp[7] ;
    input n29406;
    output \Kp[8] ;
    input n29405;
    output \Kp[9] ;
    input n29404;
    output \Kp[10] ;
    input n29403;
    output \Kp[11] ;
    input n29402;
    output \Kp[12] ;
    input n29401;
    output \Kp[13] ;
    input n29400;
    output \Kp[14] ;
    input n29396;
    output \Kp[15] ;
    input n29395;
    output \Ki[1] ;
    input n29394;
    output \Ki[2] ;
    input n29391;
    output \Ki[3] ;
    input n29390;
    output \Ki[4] ;
    input n29389;
    output \Ki[5] ;
    input n29388;
    output \Ki[6] ;
    input n29387;
    output \Ki[7] ;
    input n29386;
    output \Ki[8] ;
    input n29385;
    output \Ki[9] ;
    input n29384;
    output \Ki[10] ;
    input n29378;
    output \Ki[11] ;
    input n29377;
    output \Ki[12] ;
    input n29376;
    output \Ki[13] ;
    input n29375;
    output \Ki[14] ;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[24] ;
    input n29374;
    output \Ki[15] ;
    input n29373;
    input n29372;
    input n29371;
    input n29370;
    input n29369;
    input n29368;
    input n29366;
    input n29365;
    input n29364;
    input n29363;
    input n29362;
    input n29361;
    input n29360;
    input n29358;
    input n29355;
    input n29354;
    input n29353;
    input n29352;
    input n29351;
    input n29349;
    input n29347;
    input n29346;
    input n29345;
    input n29343;
    input n29341;
    input n29340;
    input n29339;
    input n29338;
    input n29337;
    input n29336;
    input n29335;
    input n29334;
    input n29333;
    input n29332;
    input n29331;
    input n29330;
    input n29329;
    input n29328;
    input n29327;
    input n29326;
    input n29325;
    input n29323;
    input n29322;
    output n50602;
    output n122;
    output \FRAME_MATCHER.i_31__N_2843 ;
    output n5;
    output n57092;
    input n29321;
    input n29957;
    input n29956;
    input n29955;
    input n29954;
    input n29953;
    input n29952;
    input n29951;
    input n29950;
    input n29949;
    input n29948;
    input n29947;
    input n29946;
    input n29945;
    input n29944;
    input n29943;
    input n29942;
    input n29941;
    input n29940;
    input n29939;
    input n29938;
    input n29937;
    input n29936;
    input n29935;
    input n29934;
    input n29933;
    input n29932;
    input n29931;
    input n29930;
    input n29929;
    input n29928;
    input n29927;
    input n29926;
    input n29925;
    input n29924;
    input n29923;
    input n29922;
    input n29921;
    input n29920;
    input n29919;
    input n29918;
    input n29917;
    input n29916;
    input n29915;
    input n29914;
    input n29913;
    input n29912;
    input n29911;
    input n29910;
    input n29909;
    input n29908;
    input n29907;
    input n29906;
    input n29905;
    input n29904;
    input n29903;
    input n29902;
    input n29901;
    input n29900;
    input n29899;
    input n29898;
    input n29897;
    input n29896;
    input n29895;
    input n29894;
    input n29893;
    input n29892;
    input n29891;
    input n29890;
    input n29889;
    input n29888;
    input n29887;
    input n29886;
    input n29885;
    input n29884;
    input n29883;
    input n29882;
    output DE_c;
    output LED_c;
    input n29319;
    input n29318;
    input n29316;
    input n29315;
    input n29314;
    input n29313;
    input n29312;
    input n29311;
    input n29310;
    input n29307;
    input n29306;
    input n29305;
    input n29304;
    input n29300;
    input n29299;
    input n29298;
    input n29297;
    input n29296;
    input n29881;
    input n29880;
    input n29879;
    input n29878;
    input n29877;
    input n29876;
    input n29875;
    input n29874;
    input n29873;
    input n29872;
    input n29871;
    input n29870;
    input n29869;
    input n29868;
    input n29867;
    input n29859;
    input n29858;
    input n29857;
    input n29856;
    input n29855;
    input n29854;
    input n29853;
    input n29852;
    input n29851;
    output [7:0]control_mode;
    input n29295;
    input n29850;
    input n29849;
    input n29848;
    input n29847;
    input n29846;
    input n29845;
    input n29294;
    input n29844;
    output [15:0]current_limit;
    input n29293;
    input n29843;
    input n29842;
    input n29841;
    input n29840;
    input n29292;
    input n29291;
    input n29290;
    input n29288;
    input n29287;
    input n29286;
    input n48016;
    input n29284;
    output [23:0]PWMLimit;
    input n29283;
    input n29282;
    input n29280;
    output [23:0]neopxl_color;
    input n29279;
    input n29278;
    output \Ki[0] ;
    input n29277;
    output \Kp[0] ;
    input n29276;
    output [23:0]IntegralLimit;
    input n29275;
    input n29274;
    input n29273;
    input n29839;
    input n29838;
    input n29837;
    input n29836;
    input n29835;
    input n29834;
    output n63_adj_6;
    input n29833;
    input n29832;
    input n9;
    input n29831;
    input n29830;
    input n29829;
    input n29828;
    input n29260;
    input n29259;
    input n29827;
    input n29826;
    input n29825;
    input n29824;
    input n29823;
    input n29822;
    input n29821;
    input n29820;
    input n29256;
    input n29819;
    input n29818;
    input n29817;
    input n29816;
    input n29815;
    input n29814;
    input n29813;
    input n29812;
    input n29811;
    input n29810;
    input n29809;
    input n29808;
    input n29807;
    input n56702;
    input n29762;
    input n29761;
    input n29760;
    input n29759;
    input n29758;
    input n29757;
    input n29756;
    input n29755;
    input n29754;
    input n29753;
    input n29752;
    input n29751;
    input n29726;
    input n29725;
    input n29724;
    input n29723;
    input n29722;
    input n29721;
    input n29720;
    input n29719;
    input n29718;
    input n29717;
    input n29716;
    input n29707;
    input n29706;
    input n29705;
    input n29704;
    input n29703;
    input n29702;
    input n29701;
    input n29687;
    input n29686;
    input n29685;
    input n29666;
    input n29665;
    input n29664;
    input n29663;
    input n29662;
    input n29661;
    input n29660;
    input n29659;
    input n29658;
    input n29657;
    input n29656;
    input n29655;
    input n29654;
    input n29653;
    input n29652;
    input n29651;
    input n29650;
    input n29649;
    input n29648;
    input n29646;
    input n29645;
    input n29644;
    input n29643;
    input n29483;
    input n29482;
    input n29481;
    input n29480;
    input n29479;
    input n29478;
    input n29477;
    input n29476;
    input n29468;
    input n29467;
    input n29466;
    input n29465;
    input n29464;
    input n29463;
    input n29462;
    input n29461;
    input n29460;
    input n29459;
    input n29458;
    input n29457;
    input n29456;
    input n29455;
    input n29454;
    input n29453;
    input n29452;
    input n29451;
    input n29450;
    input n29449;
    input n29448;
    input n29447;
    input n29446;
    input n29445;
    output \Kp[1] ;
    input n29442;
    input n29441;
    input n29440;
    input n29439;
    input n29438;
    input n29437;
    input n29434;
    input n29433;
    input n29432;
    input n29431;
    input n29430;
    input n29429;
    input n29428;
    output n5_adj_7;
    output n50620;
    output n24373;
    output n48646;
    output n48638;
    input \state[0] ;
    input \state[2] ;
    input \state[3] ;
    output n7936;
    output n28758;
    output n29184;
    output \r_Bit_Index[0] ;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3848[1] ;
    input VCC_net;
    output tx_o;
    input n29324;
    input n29732;
    input n56700;
    output n4_adj_8;
    output tx_enable;
    output n19731;
    output n28762;
    output n29186;
    input n29420;
    output [2:0]r_SM_Main_adj_16;
    output r_Rx_Data;
    output \r_SM_Main_2__N_3777[2] ;
    output n35837;
    input RX_N_10;
    output n4_adj_12;
    output n4_adj_13;
    input n29735;
    output \r_Bit_Index[0]_adj_14 ;
    input n48270;
    input n29261;
    output n4_adj_15;
    input n29769;
    input n29767;
    input n29766;
    input n48565;
    input n29749;
    input n29748;
    input n29740;
    output n27227;
    output n27232;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n56584, n56533, n7;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(103[12:33])
    wire [7:0]tx_data;   // verilog/coms.v(106[13:20])
    
    wire n56437, n54306, n56578;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(116[11:12])
    
    wire n4623, n3, n28010, n4_c, n8, n48649, n29603, n2, n3_adj_4624, 
        n45442, n6, n49029, n8_adj_4625;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(97[12:25])
    
    wire n29636, n49308, n29637;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(97[12:25])
    
    wire n52138, n29638, n53050, n52140, n53048, n29639, n27961, 
        n49403, n49284, n49400, n52148, n56563, n54307, n27208, 
        n4_adj_4626, n2_adj_4627;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(113[11:16])
    
    wire n48182, n49397, n49321, n52152, n48983, n28107, Kp_23__N_1398, 
        n52158;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(97[12:25])
    
    wire n7672, n7674, n7675, n3_adj_4628, n7676, n45492, n45488, 
        n49299, n52164, n7677, n7678, n7679, n7680;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(97[12:25])
    
    wire n7681, n7682, n7683, n56647, n54301, n7684, n7685, n7686, 
        n48749, n46462, n45524, n52170, n29640, n7687, n7688, 
        n7689, n7690, n46365, n48986, n7691, n7692, n7693, n7694, 
        n7695, n7696, n29641, n7_adj_4629, n50318, n48942, n29642, 
        n29281, n52988, n52989, n52893, n52892, n10, n52973, n52974, 
        n52884, n52883, n56299, n54305, n45424, n49358, n48781, 
        n52184, n51079, n35747, n48658, n10_adj_4630, n8_adj_4631, 
        n29588, n49165, n45137, n49406, n48184, Kp_23__N_1602, n48936, 
        n27621, n48758;
    wire [0:0]n6223;
    wire [2:0]r_SM_Main_2__N_3851;
    
    wire n7824, n3_adj_4632;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(97[12:25])
    
    wire n52508, n27556, n52514, n28328, n26308, n48811, n27946, 
        n3_adj_4633, n3_adj_4634, n49170, n3_adj_4635, n3_adj_4636, 
        n3_adj_4637, n3_adj_4638, n3_adj_4639, n49052, n48799, n10_adj_4640, 
        n25573, n3_adj_4641, n3_adj_4642, n3_adj_4643, n29589, n52801, 
        n3_adj_4644, n27328, n15, n27114;
    wire [7:0]\data_in[1]_c ;   // verilog/coms.v(96[12:19])
    
    wire n10_adj_4645;
    wire [7:0]\data_in[2]_c ;   // verilog/coms.v(96[12:19])
    
    wire n3_adj_4646, n16, n29590, n17, n29591;
    wire [7:0]\data_in[3]_c ;   // verilog/coms.v(96[12:19])
    
    wire n5_c, n29592, n46475, n50466, n10_adj_4647;
    wire [7:0]\data_in[0]_c ;   // verilog/coms.v(96[12:19])
    
    wire n14, n27291, n18, \FRAME_MATCHER.rx_data_ready_prev , n161, 
        n20, n15_adj_4648, n63_c, n27661, n49004, n49393, n49420, 
        n20_adj_4649, n19, n52807, n16_adj_4651, n17_adj_4652, n49363, 
        n63_adj_4653, n27244, n5_adj_4654, n771, n36594, n6_adj_4655, 
        tx_transmit_N_3748, n3_adj_4656, n3_adj_4657, n11, n144, n21, 
        n3_adj_4658, n3_adj_4659, n16_adj_4660, n3_adj_4661, n3_adj_4662, 
        n3_adj_4663, n3_adj_4664, n15_adj_4665, n27325, n27132, n48820, 
        n49387, n49176, n17_adj_4666, n44, n42, n43, n41, n48881, 
        n40, n39, n50, n45, n48722, \FRAME_MATCHER.i_31__N_2839 , 
        n29593, n56377, n7_adj_4668, n27465, n29594, n29595, n27583, 
        n28384, n4_adj_4669, n27549, n27685, n48847, n48878, n46432, 
        n28078, n6_adj_4670, n46531, n48893, n48718, n49149, n6_adj_4671, 
        n48887, n27916, Kp_23__N_1130, n48958, Kp_23__N_1174, n48805, 
        n49198, n45988, n45537, n49415, n27564, n52620, n27570, 
        n28047, n14_adj_4672, n27506, n10_adj_4673, n50634, n46502, 
        n45470, n28075, n20_adj_4674, n28032, n19_adj_4675, n45422, 
        n27639, n27601, n27649, n21_adj_4676, n6_adj_4677, n52102, 
        n7_adj_4678, n27913, n31, n52104, n31_adj_4679, n23547, 
        n52106, n52961, n48641, n24561, n28627, n7673, n52962, 
        n52911, n52910, n49999, n29580, n29581, n12, n52114, n10_adj_4680, 
        n48919, n49204, n52118, n52116, n49069, n52124, n27445, 
        n49087, Kp_23__N_1206, n29582, n52594, n52596, n49384, n48768, 
        n52602, n52608, n45436, n48925, n52614, n2_adj_4681, n49257, 
        n52952, n52953, n11_adj_4682, n2_adj_4683, n52944, n52943, 
        n29583, n52891, n2_adj_4684, n52889, n2_adj_4685, n2_adj_4686, 
        n29414;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(97[12:25])
    
    wire n29413, n2_adj_4687, n29584, n2_adj_4688, n9_c, n2_adj_4689, 
        n27631, n49084, n52946, n52947, n49012, n45384, n50425, 
        n2_adj_4690, n35749, n52983, n52982, n48736, n46448, n48960, 
        n10_adj_4691, n2_adj_4692, n50208, n48974;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(98[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(98[12:26])
    
    wire n56572, n52916, n2_adj_4693, n49333, n50850, n2_adj_4694, 
        n2_adj_4695, n50005, n8_adj_4696, n52917, n2_adj_4697, n52998, 
        n52252, n2_adj_4698, n52997, n46240, n48679, n118, n45510, 
        n46389, n46481, n6_adj_4699, n2_adj_4700, n53042, n36499, 
        n53043, n29585, n105, n27239, n2_adj_4701, n56717, n11_adj_4702, 
        n2_adj_4703, n46429, n52522, n52902, n48560, n176, n41981, 
        n52901, n28717, n49010, n46415, n52672, n46577, n29586, 
        n52666, n56614, n56617, n29587, n49105, n52226, n52228, 
        n52863, n49127, n49318, n52234, n52864, n52862, n49248, 
        n52240, n52202, n29523, n52204, n56431, n52208, n46393, 
        n49272, n52214, n52904, n52905, n53016, n2_adj_4704, n53015, 
        n52928, n52929, n52935, n48681, n49426, n52220, n50753, 
        n29572, n46407, n52244, n46363, n52934, n52949, n52950, 
        n52959, n52958, n52955, n7_adj_4705, n52956, n52923, n52922, 
        n29573, n29574, n29575, n29576, n49305, n14_adj_4706, n29577, 
        n56389, n56608, n56497, n7_adj_4707, n29578, n1;
    wire [31:0]\FRAME_MATCHER.state_31__N_2943 ;
    
    wire n13, n29579, n48644, n49096, n13_adj_4708, n52254;
    wire [7:0]n9046;
    
    wire n28649, n29210, Kp_23__N_1587, n6_adj_4709, n49351, n49173, 
        n8_adj_4710, n29564, n49151, n48728, n52644, n27969, n49423, 
        n48742, n29565, n51116, n49296, n50394, n29566, n27608, 
        Kp_23__N_1536, Kp_23__N_1539, n2_adj_4711, n56575, n45514, 
        n48992, n50581, n52258, n46426, n49266, n2_adj_4712, n3_adj_4713, 
        n2_adj_4714, n3_adj_4715, n29567, n27822, n28335, n8_adj_4716, 
        n29568, n52260, n52262, n50588, n50811, n29367, n52360, 
        Kp_23__N_1098, n46436, n29569, n50405, n28051, n49230, n29359, 
        n29356, n56566, n49007, n52436, n52328, n52334, n29570, 
        n52450, n52268, n27590, n29571, n28477, n52442, n52454, 
        Kp_23__N_1324, n49207, n49045, n52272, n49336, n50889, n45486, 
        n52274, n8_adj_4717, n29556, n28295, n52580, n49245, n52584, 
        n52919, n52920, n29557, n35692, n29348, n35686, n35689, 
        n28105, n48817, n52590, n56569, n56560, n48773, n53004, 
        n53003, n50782, n50686, n50306, n50411, n50065, n29558, 
        n52895, n52896, n29559, n50541, n50073, n50544, n50966, 
        n49279, n48945, n27615, n12_adj_4718, n52913, n52914, n56530, 
        n52908, n52907, n50662, n53046, n53045, n50903, n46444, 
        n29560, n6_adj_4719, n27669, n50534, n29561, n52426, n27119, 
        n56641, n50504, n51075, n2_adj_4720, n3_adj_4721, n2_adj_4722, 
        n3_adj_4723, n45569, n49093, n48971, n52472, n52478, n48916, 
        n48922, n49157, n52484, n49260, n52490, n46409, n48704, 
        n29562, n29563, n2_adj_4725, n3_adj_4726, n2_adj_4727, n3_adj_4728, 
        n2_adj_4729, n3_adj_4730, n52881, n52528, n52882, n52880, 
        n52552, n10_adj_4731, n48905, n12_adj_4732, n49192, n52544, 
        n48866, Kp_23__N_1203, n28387, n48710, n49201, n10_adj_4733, 
        n27922, Kp_23__N_1416, n48731, n49154, n48896, n45132, n52080, 
        n45522, n45571, n49167, n52700, n28353, n46500, n52300, 
        n52314, n49354, n52320, n48967, n52306, n52326, n46367, 
        n52898, n52899, n56494, n52344, n49189, n28468, n52965, 
        n52964, n8_adj_4734, n29548, n4_adj_4735, n52458, n49263, 
        n29549, n28129, n29550, n27515, n27552, n6_adj_4736, n6_adj_4737, 
        n46507, n43271, n43270, n43269, n29551, n27278, n171, 
        n124, n29552, n29040, n49607, n56488, n56491, n56482, 
        n56485, n56476, n56479, n56470, n56473, n29553, n29554, 
        n29555, n52678, n48796, n56434, n43268, n56428, n29866, 
        n56422, n29865, n56425, n29864, n29863, n56416, n29862, 
        n56419, n29861, n29860, n56398, n56401, n3_adj_4738, n52284, 
        n52288, n48933, n43267, n56602, n43266, n48674, n48086, 
        n48084, n56386, n56374;
    wire [31:0]n92;
    
    wire n5_adj_4739, n44910, n1_adj_4741, n56701, n48110, n48102, 
        n48082, n43265, n48080, n48078, n43264, n3746, n43263, 
        n43262, n43261, n43260, n43259, n43258, n4_adj_4742, n7_adj_4744, 
        n48114, n48076, n46498, n46440, n12_adj_4745, n48012, n49074, 
        n5_adj_4746, n48014, n46052, n48995, n45453, n50908, n12_adj_4747, 
        n46477, n49278, n48074, n48096, n49114, n6_adj_4748, n43257, 
        n49275, n49375, n49217, n22, n48094, n51165, n49293, n45480, 
        n20_adj_4749, n15_adj_4750, n49269, n50160, n24, n48072, 
        n48092, n2_adj_4751, n43256, n48090, n2_adj_4752, n43255, 
        n2_adj_4753, n43254, n2_adj_4754, n43253, n43252, n48088, 
        n43251, n48018, n27448, n49020, n50561, n12_adj_4755, n51086, 
        n49118, n50784, n46456, n51199, n43250, n50467, n50101, 
        n49064, n49287, n49075, n56590, n7_adj_4756, n48665, n29508, 
        n29509, n29510, n29511, n2520, n49195, n29512, n48048, 
        n29513, n29514, n48050, n48180, n48052, n48178, n48054, 
        n48176, n48056, n48174, n48058, n48172, n48060, n48170, 
        n48062, n48168, n48064, n48166, n48066, n48164, n48068, 
        n48162, n48070, n48160, n48158, n48156, n48150, n48142, 
        n48134, n48132, n48130, n48128, n48126, n48124, n48122, 
        n48120, n48118, n48116, n48010, n48980, n29515, n43249, 
        n27421, n49026, n10_adj_4757, n43248, n43247, n43246, n27905, 
        n48964, n43245, n43244, n43243, n43242, n29500, n43241, 
        n43240, n29501, n43239, n43238, n49061, n43237, n29502, 
        n29503, n29504, n4_adj_4758, n46452, n49342, n46387, n7_adj_4759, 
        n43236, n29505, n29506, n29507, n43235, n43234, n49214, 
        n8_adj_4760, n4_adj_4761, n28257, n48823, n48861, n49130, 
        n29492, n50938, n48952, n28410, n29493, n46504, n48707, 
        n29494, n29495, n45389, n48701, n49330, n6_adj_4762, n49042, 
        n50783, n28094, n14_adj_4763, n46454, n49139, n13_adj_4764, 
        n29496, n56326, n8_adj_4765, n56329, n56320, n45478, n48955, 
        n12_adj_4766, n29497, n26, n56323, n29498, n29499, n41963, 
        n27894, n19_adj_4767, Kp_23__N_1079, n52716, n48850, n45604, 
        n24_adj_4768, n29484, n28, n29485, n16_adj_4769, n29486, 
        n29487, n29488, n29489, n29490, n50646, n27153, n29491, 
        n48755, n6_adj_4770, n56656, n48989, n26792, n49019, n10_adj_4771, 
        n45590, n26789, n56659, n49039, n6_adj_4772, n28318, n27985, 
        n7_adj_4773, n29635, n29634, n29633, n29632, n29631, n29630, 
        n29629, n29628, n29627, n29626, n29625, n29624, n29623, 
        n29622, n29621, n29620, n29619, n29618, n29617, n29616, 
        n29615, n29614, n29613, n29612, n29611, n29610, n29609, 
        n29608, n29607, n29606, n29605, n29604, n29602, n29601, 
        n29600, n29599, n29598, n29597, n29596, n48802, n49180, 
        n49372, n16_adj_4774, n29547, n29546, n29545, n29544, n29543, 
        n29542, n29541, n29540, n29539, n29538, n29537, n29536, 
        n29535, n29534, n29533, n29532, n29531, n29530, n29529, 
        n29528, n29527, n29526, n46395, n49315, n50720, n49090, 
        n17_adj_4775, n29525, n29524, n29522, n29521, n29520, n29519, 
        n46513, n1247, n10_adj_4776, n46138, n49034, n29518, n29517, 
        n29516, n29475, n29474, n29473, n29472, n29471, n29470, 
        n29469, n10_adj_4777, n49220, n45438, n10_adj_4778, n28275, 
        n56650, n56653, n28401, n25317, n10_adj_4779, n48687, n49186, 
        n14_adj_4780, n27347, n28289, n27848, n49000, n10_adj_4781, 
        n50826, n6_adj_4782, n48858, n48690, n10_adj_4783, n28140, 
        n45376, n48853, n27863, n49226, n45584, n49302, n49327, 
        n6_adj_4784, n48834, n8_adj_4785, n27580, n9_adj_4786, n49077, 
        n49082, n49339, n49162, n46403, n48684, n49312, n48746, 
        n10_adj_4787, n48713, n48939, n12_adj_4788, n28394, n49210, 
        n1191, n48725, n1168, n49145, n49239, n10_adj_4789, n17_adj_4790, 
        n10_adj_4791, n49345, n48890, n14_adj_4792, n48884, n10_adj_4793, 
        n10_adj_4794, n48739, n4_adj_4795, n48912, n46610, n27343, 
        n28_adj_4796, n1182, n48841, n26_adj_4797, n28398, n27, 
        n25, n51207, n48930, n49233, n49378, n16_adj_4798, n49251, 
        n49108, n17_adj_4799, n49079, n51208, n10_adj_4800, n49324, 
        n6_adj_4801, n49111, n25447, n49048, n10_adj_4802, n46361, 
        n6_adj_4803, n28_adj_4804, n26_adj_4805, n48977, n27_adj_4806, 
        n25_adj_4807, n54303, n56596, n26997, n52875, n46520, n13_adj_4808, 
        n28381, n52876, n14_adj_4809, n15_adj_4810, n49121, n52874, 
        n49429, n6_adj_4811, n46391, n49348, n49183, n49366, n48789, 
        n49023, n28143, n7_adj_4812, n10_adj_4813, n49142, n48645, 
        n27576, n10_adj_4814, n49369, n46599, n48844, n1519, n1516, 
        n27356, n27711, n165, n48902, n49242, n27891, n40_adj_4815, 
        n38, n39_adj_4816, n37, n42_adj_4817, n46, n41_adj_4818, 
        n12_adj_4819, n13_adj_4820, n46355, n14_adj_4821, n48872, 
        n6_adj_4822, n10_adj_4823, n50291, n18_adj_4824, n19_adj_4825, 
        n49254, n10_adj_4826, n14_adj_4827, n56644, n50278, n49136, 
        n49412, n6_adj_4829, n49056, n10_adj_4830, n6_adj_4831, n14_adj_4832, 
        n49133, n15_adj_4833, n48838, n6_adj_4834, n49223, n10_adj_4835, 
        n53035, n53033, n7_adj_4836, n52870, n52868, n7_adj_4837, 
        n53026, n53024, n7_adj_4838, n14_adj_4839, n56638, n1668, 
        n14_adj_4840, n8_adj_4841, n7_adj_4842, n6_adj_4843, n56293, 
        n14_adj_4844, n54289, n54302, n52869, n54300, n56626, n53025, 
        n48899, n57, n23, n26_adj_4845, n29, n22_adj_4846, n32, 
        n27_adj_4847, n56296, n6_adj_4848, n16_adj_4849, n56290, n17_adj_4850, 
        n50821, n12_adj_4851, n10_adj_4852, n14_adj_4853, n56620;
    
    SB_LUT4 n56584_bdd_4_lut (.I0(n56584), .I1(n56533), .I2(n7), .I3(byte_transmit_counter[4]), 
            .O(tx_data[2]));
    defparam n56584_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_40739 (.I0(byte_transmit_counter[3]), 
            .I1(n56437), .I2(n54306), .I3(byte_transmit_counter[4]), .O(n56578));
    defparam byte_transmit_counter_3__bdd_4_lut_40739.LUT_INIT = 16'he4aa;
    SB_DFF deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n29426));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n29425));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n29424));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n29423));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n29422));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 select_713_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_713_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[16] [5]), .I1(n28010), .I2(GND_net), 
            .I3(GND_net), .O(n4_c));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15527_3_lut_4_lut (.I0(n8), .I1(n48649), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n29603));
    defparam i15527_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n29421));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk16MHz), 
            .D(n2), .S(n3_adj_4624));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut (.I0(\data_in_frame[14] [3]), .I1(n45442), .I2(n6), 
            .I3(\data_in_frame[12] [2]), .O(n49029));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i15560_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48649), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n29636));
    defparam i15560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_956 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49308));
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h6666;
    SB_LUT4 i15561_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48649), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n29637));
    defparam i15561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_957 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[17] [0]), 
            .I2(\data_in_frame[16] [6]), .I3(\data_in_frame[15] [7]), .O(n52138));
    defparam i1_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 i15562_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48649), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n29638));
    defparam i15562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37258_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n53050));
    defparam i37258_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i1_4_lut_adj_958 (.I0(n52138), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[10] [6]), .I3(\data_in_frame[17] [3]), .O(n52140));
    defparam i1_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_LUT4 i37256_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53048));
    defparam i37256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15563_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48649), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n29639));
    defparam i15563_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_959 (.I0(n27961), .I1(n49403), .I2(n49284), .I3(n49400), 
            .O(n52148));
    defparam i1_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i38632_2_lut (.I0(n56563), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54307));
    defparam i38632_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [29]), .O(n48182));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i1_4_lut_adj_960 (.I0(n52148), .I1(n49397), .I2(n49321), .I3(n52140), 
            .O(n52152));
    defparam i1_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2845 ), .I2(n22902), 
            .I3(GND_net), .O(n2_adj_4627));   // verilog/coms.v(260[6] 262[9])
    defparam i2_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_4_lut_adj_961 (.I0(n48983), .I1(n28107), .I2(Kp_23__N_1398), 
            .I3(n52152), .O(n52158));
    defparam i1_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2112_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n7672), .I3(GND_net), .O(n7674));
    defparam mux_2112_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n7672), .I3(GND_net), .O(n7675));
    defparam mux_2112_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_713_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4628));
    defparam select_713_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_2112_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n7672), .I3(GND_net), .O(n7676));
    defparam mux_2112_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_962 (.I0(n45492), .I1(n45488), .I2(n49299), .I3(n52158), 
            .O(n52164));
    defparam i1_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2112_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n7672), .I3(GND_net), .O(n7677));
    defparam mux_2112_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n7672), .I3(GND_net), .O(n7678));
    defparam mux_2112_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n7672), .I3(GND_net), .O(n7679));
    defparam mux_2112_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n29419));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 mux_2112_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n7672), .I3(GND_net), .O(n7680));
    defparam mux_2112_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n7672), .I3(GND_net), .O(n7681));
    defparam mux_2112_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n7672), .I3(GND_net), .O(n7682));
    defparam mux_2112_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n7672), .I3(GND_net), .O(n7683));
    defparam mux_2112_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38750_2_lut (.I0(n56647), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54301));
    defparam i38750_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_2112_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n7672), .I3(GND_net), .O(n7684));
    defparam mux_2112_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n7672), .I3(GND_net), .O(n7685));
    defparam mux_2112_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n7672), .I3(GND_net), .O(n7686));
    defparam mux_2112_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_963 (.I0(n48749), .I1(n46462), .I2(n45524), .I3(n52164), 
            .O(n52170));
    defparam i1_4_lut_adj_963.LUT_INIT = 16'h9669;
    SB_LUT4 i15564_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48649), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n29640));
    defparam i15564_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_2112_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n7672), .I3(GND_net), .O(n7687));
    defparam mux_2112_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n7672), .I3(GND_net), .O(n7688));
    defparam mux_2112_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n7672), .I3(GND_net), .O(n7689));
    defparam mux_2112_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n7672), .I3(GND_net), .O(n7690));
    defparam mux_2112_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_964 (.I0(\data_in_frame[21] [1]), .I1(n46365), 
            .I2(GND_net), .I3(GND_net), .O(n48986));
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2112_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n7672), .I3(GND_net), .O(n7691));
    defparam mux_2112_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n7672), .I3(GND_net), .O(n7692));
    defparam mux_2112_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n7672), .I3(GND_net), .O(n7693));
    defparam mux_2112_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n7672), .I3(GND_net), .O(n7694));
    defparam mux_2112_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n7672), .I3(GND_net), .O(n7695));
    defparam mux_2112_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2112_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n7672), .I3(GND_net), .O(n7696));
    defparam mux_2112_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15565_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48649), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n29641));
    defparam i15565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut (.I0(n7_adj_4629), .I1(\data_in_frame[18] [6]), .I2(\data_in_frame[21] [0]), 
            .I3(n50318), .O(n48942));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i15566_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48649), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n29642));
    defparam i15566_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15205_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48649), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n29281));
    defparam i15205_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37196_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52988));
    defparam i37196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37197_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52989));
    defparam i37197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37101_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52893));
    defparam i37101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37100_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52892));
    defparam i37100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_340_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10));   // verilog/coms.v(155[7:23])
    defparam equal_340_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i37181_3_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52973));
    defparam i37181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37182_3_lut (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52974));
    defparam i37182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37092_3_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52884));
    defparam i37092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37091_3_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[21] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52883));
    defparam i37091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38749_2_lut (.I0(n56299), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54305));
    defparam i38749_2_lut.LUT_INIT = 16'h2222;
    SB_DFF deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n29418));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_965 (.I0(n45424), .I1(n49358), .I2(n48781), .I3(n52184), 
            .O(n51079));
    defparam i1_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_966 (.I0(n35747), .I1(n10), .I2(GND_net), .I3(GND_net), 
            .O(n48658));
    defparam i1_2_lut_adj_966.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_348_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4630));   // verilog/coms.v(155[7:23])
    defparam equal_348_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15512_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48649), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n29588));
    defparam i15512_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n29417));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_967 (.I0(\data_in_frame[18] [5]), .I1(n49165), 
            .I2(n51079), .I3(n45137), .O(n49406));
    defparam i1_4_lut_adj_967.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_968 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [30]), .O(n48184));
    defparam i1_2_lut_4_lut_adj_968.LUT_INIT = 16'hf800;
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[16] [2]), .I1(Kp_23__N_1602), .I2(n48936), 
            .I3(n27621), .O(n48983));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_969 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n48758));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_DFFSR tx_transmit_4011 (.Q(r_SM_Main_2__N_3851[0]), .C(clk16MHz), 
            .D(n6223[0]), .R(n7824));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 select_713_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4632));
    defparam select_713_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n52508));
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_971 (.I0(n27556), .I1(\data_in_frame[2] [7]), .I2(n52508), 
            .I3(\data_in_frame[4] [6]), .O(n52514));
    defparam i1_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_972 (.I0(n28328), .I1(n26308), .I2(n48811), .I3(n52514), 
            .O(n27946));
    defparam i1_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 select_713_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4633));
    defparam select_713_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4634));
    defparam select_713_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_973 (.I0(\data_in_frame[14] [0]), .I1(n27946), 
            .I2(n49170), .I3(\data_in_frame[9] [4]), .O(n48936));
    defparam i3_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_974 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[16] [1]), 
            .I2(\data_in_frame[16] [0]), .I3(GND_net), .O(n49321));   // verilog/coms.v(86[17:63])
    defparam i2_3_lut_adj_974.LUT_INIT = 16'h9696;
    SB_LUT4 select_713_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4635));
    defparam select_713_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4636));
    defparam select_713_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4637));
    defparam select_713_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4638));
    defparam select_713_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4639));
    defparam select_713_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_975 (.I0(n49052), .I1(n48799), .I2(\data_in_frame[13] [5]), 
            .I3(n49321), .O(n10_adj_4640));   // verilog/coms.v(86[17:63])
    defparam i4_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_976 (.I0(n35747), .I1(n10_adj_4630), .I2(GND_net), 
            .I3(GND_net), .O(n48649));
    defparam i1_2_lut_adj_976.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_3_lut (.I0(n48936), .I1(n10_adj_4640), .I2(\data_in_frame[13] [7]), 
            .I3(GND_net), .O(n25573));   // verilog/coms.v(86[17:63])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_713_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4641));
    defparam select_713_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4642));
    defparam select_713_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4643));
    defparam select_713_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15513_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48649), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n29589));
    defparam i15513_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37059_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [2]), .I2(\data_in[3] [0]), 
            .I3(GND_net), .O(n52801));
    defparam i37059_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_713_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4644));
    defparam select_713_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut (.I0(\data_in[1] [5]), .I1(\data_in[1] [4]), .I2(n27328), 
            .I3(\data_in[0] [3]), .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(\data_in[2] [4]), .I2(n52801), .I3(\data_in[0] [6]), 
            .O(n27114));
    defparam i8_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut_adj_977 (.I0(\data_in[1]_c [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1][1] ), .I3(\data_in[0] [4]), .O(n10_adj_4645));
    defparam i4_4_lut_adj_977.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_978 (.I0(\data_in[3] [4]), .I1(n10_adj_4645), .I2(\data_in[2]_c [7]), 
            .I3(GND_net), .O(n27328));
    defparam i5_3_lut_adj_978.LUT_INIT = 16'hdfdf;
    SB_LUT4 select_713_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4646));
    defparam select_713_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_979 (.I0(\data_in[2][5] ), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16));
    defparam i6_4_lut_adj_979.LUT_INIT = 16'hfffe;
    SB_LUT4 i15514_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48649), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n29590));
    defparam i15514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut (.I0(\data_in[1][6] ), .I1(\data_in[1][3] ), .I2(\data_in[2][0] ), 
            .I3(\data_in[1][2] ), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i15515_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48649), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n29591));
    defparam i15515_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_in[2][6] ), .I2(n16), .I3(\data_in[3]_c [7]), 
            .O(n5_c));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i15516_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48649), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n29592));
    defparam i15516_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_980 (.I0(n48983), .I1(n46475), .I2(\data_in_frame[16] [3]), 
            .I3(GND_net), .O(n50466));
    defparam i2_3_lut_adj_980.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut (.I0(\data_in[2][3] ), .I1(\data_in[3]_c [1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4647));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_981 (.I0(\data_in[0] [2]), .I1(\data_in[3][3] ), 
            .I2(\data_in[3][5] ), .I3(\data_in[0]_c [7]), .O(n14));
    defparam i6_4_lut_adj_981.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_982 (.I0(\data_in[3][6] ), .I1(n14), .I2(n10_adj_4647), 
            .I3(\data_in[2][1] ), .O(n27291));
    defparam i7_4_lut_adj_982.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_983 (.I0(\data_in[2] [4]), .I1(n27291), .I2(\data_in[1] [5]), 
            .I3(n5_c), .O(n18));
    defparam i7_4_lut_adj_983.LUT_INIT = 16'hfffd;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(154[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i9_4_lut_adj_984 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n27328), .O(n20));
    defparam i9_4_lut_adj_984.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4648));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n15_adj_4648), .I1(n20), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_c));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i3_4_lut_adj_985 (.I0(n27661), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[17] [0]), .I3(n49004), .O(n49393));
    defparam i3_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_986 (.I0(n49029), .I1(n49393), .I2(GND_net), 
            .I3(GND_net), .O(n49420));
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_987 (.I0(\data_in[2][6] ), .I1(\data_in[2][0] ), 
            .I2(n27291), .I3(\data_in[0] [5]), .O(n20_adj_4649));
    defparam i8_4_lut_adj_987.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_988 (.I0(n27114), .I1(\data_in[3]_c [7]), .I2(\data_in[1][6] ), 
            .I3(\data_in[2][5] ), .O(n19));
    defparam i7_4_lut_adj_988.LUT_INIT = 16'hfeff;
    SB_LUT4 i37065_4_lut (.I0(\data_in[0] [1]), .I1(\data_in[3] [2]), .I2(\data_in[1][2] ), 
            .I3(\data_in[1][3] ), .O(n52807));
    defparam i37065_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n52807), .I1(n19), .I2(n20_adj_4649), .I3(GND_net), 
            .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i6_4_lut_adj_989 (.I0(n5_c), .I1(\data_in[0]_c [7]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3][6] ), .O(n16_adj_4651));
    defparam i6_4_lut_adj_989.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_990 (.I0(n27114), .I1(\data_in[3][3] ), .I2(\data_in[2][3] ), 
            .I3(\data_in[2][1] ), .O(n17_adj_4652));
    defparam i7_4_lut_adj_990.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_adj_991 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49363));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_992 (.I0(n17_adj_4652), .I1(\data_in[3][5] ), .I2(n16_adj_4651), 
            .I3(\data_in[3]_c [1]), .O(n63_adj_4653));
    defparam i9_4_lut_adj_992.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_993 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27244));   // verilog/coms.v(255[5:25])
    defparam i1_2_lut_adj_993.LUT_INIT = 16'hbbbb;
    SB_LUT4 i21891_4_lut (.I0(n5_adj_4654), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(158[9:60])
    defparam i21891_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i40484_2_lut (.I0(n36594), .I1(n6_adj_4655), .I2(GND_net), 
            .I3(GND_net), .O(tx_transmit_N_3748));
    defparam i40484_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 select_713_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4656));
    defparam select_713_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4657));
    defparam select_713_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27_3_lut (.I0(n11), .I1(n144), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n21));
    defparam i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_713_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4658));
    defparam select_713_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4659));
    defparam select_713_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_994 (.I0(\data_in_frame[21] [2]), .I1(n49363), 
            .I2(\data_in_frame[18] [7]), .I3(n49420), .O(n16_adj_4660));
    defparam i6_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 select_713_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4661));
    defparam select_713_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4662));
    defparam select_713_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4663));
    defparam select_713_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4664));
    defparam select_713_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_2_lut (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4665));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_995 (.I0(\FRAME_MATCHER.i [4]), .I1(n27325), .I2(GND_net), 
            .I3(GND_net), .O(n27132));   // verilog/coms.v(155[7:23])
    defparam i1_2_lut_adj_995.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_996 (.I0(n48820), .I1(n49387), .I2(\data_in_frame[19] [2]), 
            .I3(n49176), .O(n17_adj_4666));
    defparam i7_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_LUT4 i21892_4_lut (.I0(n8_adj_4625), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27132), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(228[9:54])
    defparam i21892_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(\data_in_frame[21] [3]), .I1(n17_adj_4666), .I2(n15_adj_4665), 
            .I3(n16_adj_4660), .O(n48881));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40), .O(n27325));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21893_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27325), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(260[9:58])
    defparam i21893_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_997 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n48722));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_998 (.I0(n4599), .I1(n4_adj_4626), .I2(GND_net), 
            .I3(GND_net), .O(n48672));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_999 (.I0(\FRAME_MATCHER.i_31__N_2839 ), .I1(n771), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/coms.v(158[6] 160[9])
    defparam i1_2_lut_adj_999.LUT_INIT = 16'h2222;
    SB_LUT4 i15517_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48649), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n29593));
    defparam i15517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n56578_bdd_4_lut (.I0(n56578), .I1(n56377), .I2(n7_adj_4668), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n56578_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1000 (.I0(\FRAME_MATCHER.i_31__N_2845 ), .I1(n4452), 
            .I2(GND_net), .I3(GND_net), .O(n48616));
    defparam i1_2_lut_adj_1000.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1001 (.I0(n63_adj_4653), .I1(n63), .I2(n63_c), 
            .I3(GND_net), .O(n22902));   // verilog/coms.v(158[6] 160[9])
    defparam i2_3_lut_adj_1001.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1002 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27465));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'h6666;
    SB_LUT4 i15518_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48649), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n29594));
    defparam i15518_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15519_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48649), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n29595));
    defparam i15519_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut (.I0(n27583), .I1(n28384), .I2(\data_in_frame[8] [2]), 
            .I3(GND_net), .O(n4_adj_4669));   // verilog/coms.v(77[16:43])
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1003 (.I0(n27549), .I1(n27685), .I2(n48847), 
            .I3(\data_in_frame[5] [5]), .O(n48878));
    defparam i1_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1004 (.I0(n46432), .I1(n27465), .I2(n28078), 
            .I3(n6_adj_4670), .O(n46531));
    defparam i4_4_lut_adj_1004.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1005 (.I0(n48893), .I1(n48718), .I2(\data_in_frame[6] [0]), 
            .I3(GND_net), .O(n49149));   // verilog/coms.v(86[17:28])
    defparam i1_3_lut_adj_1005.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1006 (.I0(n6_adj_4671), .I1(n48887), .I2(\data_in_frame[6] [6]), 
            .I3(GND_net), .O(n27916));   // verilog/coms.v(75[16:43])
    defparam i1_3_lut_adj_1006.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1007 (.I0(Kp_23__N_1130), .I1(n49149), .I2(n48878), 
            .I3(\data_in_frame[7] [7]), .O(n48958));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1007.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_1__4__I_0_2_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1174));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_1__4__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1008 (.I0(n48805), .I1(n49198), .I2(Kp_23__N_1174), 
            .I3(\data_in_frame[3] [5]), .O(n45988));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(\data_in_frame[4] [5]), .I1(n45537), 
            .I2(GND_net), .I3(GND_net), .O(n48718));
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1010 (.I0(\data_in_frame[6] [7]), .I1(n49415), 
            .I2(\data_in_frame[6] [6]), .I3(GND_net), .O(n48893));   // verilog/coms.v(86[17:28])
    defparam i1_3_lut_adj_1010.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1011 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n48847));
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1012 (.I0(\data_in_frame[6] [5]), .I1(n27564), 
            .I2(\data_in_frame[6] [1]), .I3(\data_in_frame[6] [2]), .O(n49415));
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52620));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1014 (.I0(n48893), .I1(n27570), .I2(n48718), 
            .I3(n28047), .O(n14_adj_4672));
    defparam i6_4_lut_adj_1014.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(n28047), .I1(n27506), .I2(n52620), 
            .I3(\data_in_frame[4] [6]), .O(n48887));   // verilog/coms.v(75[16:43])
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1016 (.I0(\data_in_frame[8] [1]), .I1(n14_adj_4672), 
            .I2(n10_adj_4673), .I3(\data_in_frame[1] [3]), .O(n50634));
    defparam i7_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1017 (.I0(n45988), .I1(\data_in_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46502));
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1018 (.I0(n45470), .I1(n28075), .I2(n50634), 
            .I3(n28078), .O(n20_adj_4674));
    defparam i8_4_lut_adj_1018.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_1019 (.I0(n48958), .I1(n28032), .I2(n27916), 
            .I3(n46502), .O(n19_adj_4675));
    defparam i7_4_lut_adj_1019.LUT_INIT = 16'hfdff;
    SB_LUT4 i9_4_lut_adj_1020 (.I0(n45422), .I1(n27639), .I2(n27601), 
            .I3(n27649), .O(n21_adj_4676));
    defparam i9_4_lut_adj_1020.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_4_lut_adj_1021 (.I0(n27946), .I1(n21_adj_4676), .I2(n19_adj_4675), 
            .I3(n20_adj_4674), .O(n6_adj_4677));
    defparam i1_4_lut_adj_1021.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1022 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[5] [1]), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[5] [6]), .O(n52102));
    defparam i1_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1023 (.I0(n7_adj_4678), .I1(n4_adj_4669), .I2(n27913), 
            .I3(n6_adj_4677), .O(n31));
    defparam i4_4_lut_adj_1023.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1024 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[0] [4]), .O(n52104));
    defparam i1_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i4697_3_lut (.I0(n31_adj_4679), .I1(n31), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n23547));
    defparam i4697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1025 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[5] [7]), .O(n52106));
    defparam i1_4_lut_adj_1025.LUT_INIT = 16'h6996;
    SB_LUT4 i37169_3_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[17] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52961));
    defparam i37169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39814_4_lut (.I0(n48641), .I1(n23547), .I2(n24561), .I3(\FRAME_MATCHER.state [2]), 
            .O(n28627));
    defparam i39814_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 mux_2112_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n7672), .I3(GND_net), .O(n7673));
    defparam mux_2112_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37170_3_lut (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[19] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52962));
    defparam i37170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37119_3_lut (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[23] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52911));
    defparam i37119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37118_3_lut (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[21] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52910));
    defparam i37118_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(rx_data_ready));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n29416));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n29415));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15504_3_lut_4_lut (.I0(n10_adj_4630), .I1(n49999), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n29580));
    defparam i15504_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n28627), .D(n7673));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15505_3_lut_4_lut (.I0(n10_adj_4630), .I1(n49999), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n29581));
    defparam i15505_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_1026 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12));   // verilog/coms.v(239[12:32])
    defparam i4_4_lut_adj_1026.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_3_lut_adj_1027 (.I0(n52104), .I1(n48847), .I2(n52102), 
            .I3(GND_net), .O(n52114));
    defparam i1_3_lut_adj_1027.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1028 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4680));   // verilog/coms.v(239[12:32])
    defparam i2_4_lut_adj_1028.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1029 (.I0(n48919), .I1(n49204), .I2(n48722), 
            .I3(n52106), .O(n52118));
    defparam i1_4_lut_adj_1029.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1030 (.I0(n52116), .I1(n49069), .I2(n52118), 
            .I3(n52114), .O(n52124));
    defparam i1_4_lut_adj_1030.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(n27445), .I1(n49087), .I2(Kp_23__N_1206), 
            .I3(n52124), .O(n45537));
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_LUT4 i15506_3_lut_4_lut (.I0(n10_adj_4630), .I1(n49999), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n29582));
    defparam i15506_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n52594));
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1033 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[7] [1]), .I3(GND_net), .O(n52596));
    defparam i1_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n49384), .I1(n52596), .I2(n48768), 
            .I3(n52594), .O(n52602));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(n45537), .I1(n48887), .I2(n49415), 
            .I3(n52602), .O(n52608));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1036 (.I0(n46531), .I1(n45436), .I2(n48925), 
            .I3(n52608), .O(n52614));
    defparam i1_4_lut_adj_1036.LUT_INIT = 16'h9669;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n2_adj_4681), .S(n3_adj_4664));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1037 (.I0(\data_in_frame[14] [2]), .I1(n52614), 
            .I2(n49257), .I3(n45442), .O(n46475));
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'h9669;
    SB_LUT4 i37160_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52952));
    defparam i37160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37161_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52953));
    defparam i37161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1038 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_4682));   // verilog/coms.v(239[12:32])
    defparam i3_4_lut_adj_1038.LUT_INIT = 16'h7bde;
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n2_adj_4683), .S(n3_adj_4661));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37152_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52944));
    defparam i37152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37151_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52943));
    defparam i37151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15507_3_lut_4_lut (.I0(n10_adj_4630), .I1(n49999), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n29583));
    defparam i15507_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i37099_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n52891));
    defparam i37099_4_lut.LUT_INIT = 16'hec2c;
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n2_adj_4684), .S(n3_adj_4658));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37097_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52889));
    defparam i37097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(\data_in_frame[16] [4]), .I1(n46475), 
            .I2(GND_net), .I3(GND_net), .O(n49176));
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'h9999;
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n2_adj_4685), .S(n3_adj_4657));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n2_adj_4686), .S(n3_adj_4656));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n29414));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n29413));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk16MHz), 
            .D(n2_adj_4687), .S(n3_adj_4646));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n29411));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1602));   // verilog/coms.v(86[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15508_3_lut_4_lut (.I0(n10_adj_4630), .I1(n49999), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n29584));
    defparam i15508_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n2_adj_4688), .S(n3_adj_4644));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1040 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_c));   // verilog/coms.v(239[12:32])
    defparam i1_4_lut_adj_1040.LUT_INIT = 16'h7bde;
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n2_adj_4689), .S(n3_adj_4643));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1041 (.I0(n27631), .I1(\data_in_frame[15] [1]), 
            .I2(n49084), .I3(GND_net), .O(n49299));
    defparam i1_3_lut_adj_1041.LUT_INIT = 16'h6969;
    SB_LUT4 i37154_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52946));
    defparam i37154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37155_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52947));
    defparam i37155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1042 (.I0(n9_c), .I1(n11_adj_4682), .I2(n10_adj_4680), 
            .I3(n12), .O(n24561));   // verilog/coms.v(239[12:32])
    defparam i7_4_lut_adj_1042.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(n49012), .I1(n45384), .I2(n50425), 
            .I3(n49299), .O(n46462));
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'h9669;
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n2_adj_4690), .S(n3_adj_4642));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_3_lut_adj_1044 (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n6_adj_4655));
    defparam i2_3_lut_adj_1044.LUT_INIT = 16'hfefe;
    SB_LUT4 i21689_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3851[0]), .I2(GND_net), 
            .I3(GND_net), .O(n35749));
    defparam i21689_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i37191_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52983));
    defparam i37191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37190_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52982));
    defparam i37190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1045 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[10] [5]), .I3(\data_in_frame[12] [7]), .O(n48736));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1045.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1046 (.I0(\data_in_frame[20] [3]), .I1(n46448), 
            .I2(\data_in_frame[22] [5]), .I3(n48960), .O(n10_adj_4691));
    defparam i4_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n2_adj_4692), .S(n3_adj_4641));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i5_3_lut_adj_1047 (.I0(\data_in_frame[20] [4]), .I1(n10_adj_4691), 
            .I2(\data_in_frame[18] [1]), .I3(GND_net), .O(n50208));
    defparam i5_3_lut_adj_1047.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n48974));
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_40764 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n56572));
    defparam byte_transmit_counter_0__bdd_4_lut_40764.LUT_INIT = 16'he4aa;
    SB_LUT4 i37124_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52916));
    defparam i37124_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n2_adj_4693), .S(n3_adj_4639));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_4_lut_adj_1049 (.I0(\data_in_frame[20] [4]), .I1(n49333), 
            .I2(\data_in_frame[20] [5]), .I3(\data_in_frame[22] [6]), .O(n50850));
    defparam i2_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n2_adj_4694), .S(n3_adj_4638));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n2_adj_4695), .S(n3_adj_4637));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1050 (.I0(n50005), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[20] [2]), .I3(\data_in_frame[20] [3]), .O(n8_adj_4696));
    defparam i3_4_lut_adj_1050.LUT_INIT = 16'h9669;
    SB_LUT4 i37125_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52917));
    defparam i37125_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n29410));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n2_adj_4697), .S(n3_adj_4636));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37206_3_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52998));
    defparam i37206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1051 (.I0(n50850), .I1(\data_in_frame[23] [4]), 
            .I2(n50208), .I3(n48881), .O(n52252));   // verilog/coms.v(269[9:85])
    defparam i1_4_lut_adj_1051.LUT_INIT = 16'hf7fd;
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n2_adj_4698), .S(n3_adj_4635));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37205_3_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[21] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52997));
    defparam i37205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(n46240), .I1(n48679), .I2(GND_net), 
            .I3(GND_net), .O(n118));
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1053 (.I0(n45510), .I1(\data_in_frame[19] [5]), 
            .I2(n46389), .I3(n46481), .O(n6_adj_4699));   // verilog/coms.v(86[17:28])
    defparam i1_4_lut_adj_1053.LUT_INIT = 16'h9669;
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n2_adj_4700), .S(n3_adj_4634));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37250_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53042));
    defparam i37250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22436_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n36499));
    defparam i22436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1054 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n36499), .I3(byte_transmit_counter[2]), .O(n36594));
    defparam i2_4_lut_adj_1054.LUT_INIT = 16'h8880;
    SB_LUT4 i37251_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53043));
    defparam i37251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15509_3_lut_4_lut (.I0(n10_adj_4630), .I1(n49999), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n29585));
    defparam i15509_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_1055 (.I0(\FRAME_MATCHER.state[0] ), .I1(n35749), 
            .I2(n6_adj_4655), .I3(n105), .O(n27239));
    defparam i3_4_lut_adj_1055.LUT_INIT = 16'hfdff;
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n2_adj_4701), .S(n3_adj_4633));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n29409));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_rep_68_2_lut (.I0(\data_in_frame[21] [5]), .I1(\data_in_frame[21] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n56717));   // verilog/coms.v(86[17:28])
    defparam i1_rep_68_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1056 (.I0(n144), .I1(n11_adj_4702), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n7824));
    defparam i1_3_lut_adj_1056.LUT_INIT = 16'hecec;
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n2_adj_4703), .S(n3_adj_4632));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1057 (.I0(n28075), .I1(n46429), .I2(n28078), 
            .I3(n52522), .O(n45488));   // verilog/coms.v(72[16:27])
    defparam i1_4_lut_adj_1057.LUT_INIT = 16'h9669;
    SB_LUT4 i37110_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52902));
    defparam i37110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(n144), .I1(n48560), .I2(GND_net), .I3(GND_net), 
            .O(n176));   // verilog/coms.v(113[11:16])
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'heeee;
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n29408));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n29407));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n29406));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n29405));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n29404));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i38_4_lut (.I0(n27239), .I1(n36594), .I2(n176), .I3(n118), 
            .O(n41981));   // verilog/coms.v(113[11:16])
    defparam i38_4_lut.LUT_INIT = 16'h1110;
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n29403));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37109_3_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[21] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52901));
    defparam i37109_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n29402));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1059 (.I0(n41981), .I1(n28717), .I2(GND_net), 
            .I3(GND_net), .O(n6223[0]));
    defparam i1_2_lut_adj_1059.LUT_INIT = 16'heeee;
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n29401));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n29400));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1060 (.I0(n45488), .I1(n49010), .I2(\data_in_frame[17] [5]), 
            .I3(GND_net), .O(n45424));
    defparam i1_3_lut_adj_1060.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1061 (.I0(n49420), .I1(n4_c), .I2(n46415), .I3(n49308), 
            .O(n52672));
    defparam i1_4_lut_adj_1061.LUT_INIT = 16'h9669;
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n29396));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n29395));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n29394));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\data_in_frame[17] [3]), .I1(n46462), 
            .I2(GND_net), .I3(GND_net), .O(n46577));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h6666;
    SB_LUT4 i15510_3_lut_4_lut (.I0(n10_adj_4630), .I1(n49999), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n29586));
    defparam i15510_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_4_lut_adj_1063 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[21] [4]), 
            .I2(\data_in_frame[21] [3]), .I3(\data_in_frame[23] [5]), .O(n52666));
    defparam i1_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 n56614_bdd_4_lut (.I0(n56614), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n56617));
    defparam n56614_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n29391));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n29390));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n29389));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n29388));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n29387));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n29386));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n29385));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n29384));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15511_3_lut_4_lut (.I0(n10_adj_4630), .I1(n49999), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n29587));
    defparam i15511_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n29378));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n29377));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1064 (.I0(\data_in_frame[20] [7]), .I1(\data_in_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49105));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1065 (.I0(\data_in_frame[20] [2]), .I1(\data_in_frame[21] [5]), 
            .I2(\data_in_frame[20] [3]), .I3(\data_in_frame[21] [6]), .O(n52226));
    defparam i1_4_lut_adj_1065.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1066 (.I0(n49105), .I1(\data_in_frame[20] [4]), 
            .I2(\data_in_frame[21] [1]), .I3(\data_in_frame[20] [5]), .O(n52228));
    defparam i1_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i37071_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52863));
    defparam i37071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1067 (.I0(n49127), .I1(n49318), .I2(n52228), 
            .I3(n52226), .O(n52234));
    defparam i1_4_lut_adj_1067.LUT_INIT = 16'h6996;
    SB_LUT4 i37072_4_lut (.I0(n52863), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n52864));
    defparam i37072_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i37070_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52862));
    defparam i37070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1068 (.I0(n49248), .I1(n46429), .I2(n48781), 
            .I3(n52234), .O(n52240));
    defparam i1_4_lut_adj_1068.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n52202));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h6666;
    SB_LUT4 i15447_3_lut_4_lut (.I0(n10), .I1(n49999), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n29523));
    defparam i15447_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_3_lut_adj_1070 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[17] [1]), 
            .I2(\data_in_frame[21] [7]), .I3(GND_net), .O(n52204));
    defparam i1_3_lut_adj_1070.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_40744 (.I0(byte_transmit_counter[3]), 
            .I1(n56431), .I2(n54301), .I3(byte_transmit_counter[4]), .O(n56584));
    defparam byte_transmit_counter_3__bdd_4_lut_40744.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(n52204), .I1(\data_in_frame[19] [7]), 
            .I2(n52202), .I3(\data_in_frame[19] [5]), .O(n52208));
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1072 (.I0(n46393), .I1(n45137), .I2(n49272), 
            .I3(n52208), .O(n52214));
    defparam i1_4_lut_adj_1072.LUT_INIT = 16'h9669;
    SB_LUT4 i37112_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52904));
    defparam i37112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37113_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52905));
    defparam i37113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37224_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53016));
    defparam i37224_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n2_adj_4704), .S(n3_adj_4628));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37223_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53015));
    defparam i37223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37136_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52928));
    defparam i37136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37137_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52929));
    defparam i37137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37143_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52935));
    defparam i37143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1073 (.I0(n48681), .I1(n49426), .I2(n46481), 
            .I3(n52214), .O(n52220));
    defparam i1_4_lut_adj_1073.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1074 (.I0(\data_in_frame[19] [1]), .I1(n49406), 
            .I2(n52220), .I3(n45510), .O(n50753));
    defparam i1_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n29376));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15496_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48658), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n29572));
    defparam i15496_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1075 (.I0(n46407), .I1(n50753), .I2(n48881), 
            .I3(n52244), .O(n46363));
    defparam i1_4_lut_adj_1075.LUT_INIT = 16'h9669;
    SB_LUT4 i37142_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52934));
    defparam i37142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37157_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52949));
    defparam i37157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37158_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52950));
    defparam i37158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37167_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52959));
    defparam i37167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37166_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52958));
    defparam i37166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37163_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52955));
    defparam i37163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1076 (.I0(\data_in_frame[22] [1]), .I1(\data_in_frame[19] [7]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n7_adj_4705));
    defparam i2_3_lut_adj_1076.LUT_INIT = 16'h9696;
    SB_LUT4 i37164_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52956));
    defparam i37164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37131_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52923));
    defparam i37131_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n29375));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37130_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52922));
    defparam i37130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15497_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48658), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n29573));
    defparam i15497_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15498_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48658), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n29574));
    defparam i15498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(\data_in_frame[15] [5]), .I1(n45384), 
            .I2(GND_net), .I3(GND_net), .O(n45492));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h6666;
    SB_LUT4 i15499_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48658), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n29575));
    defparam i15499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15500_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48658), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n29576));
    defparam i15500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1078 (.I0(n49363), .I1(n49305), .I2(\data_in_frame[19] [1]), 
            .I3(\data_in_frame[16] [5]), .O(n14_adj_4706));
    defparam i6_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i15501_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48658), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n29577));
    defparam i15501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_40769 (.I0(byte_transmit_counter[3]), 
            .I1(n56389), .I2(n54307), .I3(byte_transmit_counter[4]), .O(n56608));
    defparam byte_transmit_counter_3__bdd_4_lut_40769.LUT_INIT = 16'he4aa;
    SB_LUT4 n56608_bdd_4_lut (.I0(n56608), .I1(n56497), .I2(n7_adj_4707), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n56608_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15502_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48658), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n29578));
    defparam i15502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1079 (.I0(n1), .I1(\FRAME_MATCHER.state [1]), .I2(\FRAME_MATCHER.state [2]), 
            .I3(\FRAME_MATCHER.state_31__N_2943 [3]), .O(n13));
    defparam i1_4_lut_adj_1079.LUT_INIT = 16'ha0ac;
    SB_LUT4 i15503_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48658), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n29579));
    defparam i15503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(n46407), .I3(GND_net), .O(n49333));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i39822_4_lut (.I0(n144), .I1(n48641), .I2(n13), .I3(n11_adj_4702), 
            .O(n48644));
    defparam i39822_4_lut.LUT_INIT = 16'h0313;
    SB_LUT4 i5_4_lut (.I0(\data_in_frame[21] [2]), .I1(n48986), .I2(\data_in_frame[23] [3]), 
            .I3(n49096), .O(n13_adj_4708));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1080 (.I0(n25573), .I1(n52252), .I2(n8_adj_4696), 
            .I3(\data_in_frame[22] [4]), .O(n52254));   // verilog/coms.v(269[9:85])
    defparam i1_4_lut_adj_1080.LUT_INIT = 16'hedde;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n28649), .D(n9046[1]), .R(n29210));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i4_4_lut_adj_1081 (.I0(\data_in_frame[11] [1]), .I1(Kp_23__N_1587), 
            .I2(\data_in_frame[16] [0]), .I3(n6_adj_4709), .O(n49248));
    defparam i4_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49351));
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1083 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49403));
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[18] [0]), .I3(n49173), .O(n52184));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15488_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48658), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n29564));
    defparam i15488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1084 (.I0(n49151), .I1(n48728), .I2(n49403), 
            .I3(n49351), .O(n52644));
    defparam i1_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1085 (.I0(n27969), .I1(n49423), .I2(n48742), 
            .I3(n52644), .O(n50425));
    defparam i1_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i15489_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48658), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n29565));
    defparam i15489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1086 (.I0(\data_in_frame[15] [3]), .I1(n50425), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n51116));
    defparam i1_3_lut_adj_1086.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1087 (.I0(n46429), .I1(n49248), .I2(\data_in_frame[17] [7]), 
            .I3(GND_net), .O(n46448));
    defparam i2_3_lut_adj_1087.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1088 (.I0(n46393), .I1(n49010), .I2(\data_in_frame[17] [6]), 
            .I3(GND_net), .O(n49296));
    defparam i2_3_lut_adj_1088.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_adj_1089 (.I0(\data_in_frame[13] [2]), .I1(n50394), 
            .I2(\data_in_frame[13] [3]), .I3(GND_net), .O(n45524));
    defparam i1_3_lut_adj_1089.LUT_INIT = 16'h6969;
    SB_LUT4 i15490_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48658), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n29566));
    defparam i15490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27608));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1091 (.I0(\data_in_frame[13] [5]), .I1(Kp_23__N_1536), 
            .I2(Kp_23__N_1539), .I3(n27608), .O(n27631));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n2_adj_4711), .S(n3));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49052));
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1093 (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49400));
    defparam i1_2_lut_adj_1093.LUT_INIT = 16'h6666;
    SB_LUT4 n56572_bdd_4_lut (.I0(n56572), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n56575));
    defparam n56572_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(n45514), .I1(\data_in_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n48960));
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1095 (.I0(n49010), .I1(n49400), .I2(n49318), 
            .I3(\data_in_frame[18] [0]), .O(n50005));
    defparam i3_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1096 (.I0(n7_adj_4705), .I1(n46577), .I2(n48992), 
            .I3(n49296), .O(n50581));
    defparam i4_4_lut_adj_1096.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1097 (.I0(n50581), .I1(n52254), .I2(n13_adj_4708), 
            .I3(n14_adj_4706), .O(n52258));   // verilog/coms.v(269[9:85])
    defparam i1_4_lut_adj_1097.LUT_INIT = 16'heffe;
    SB_LUT4 i1_2_lut_adj_1098 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27961));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1099 (.I0(\data_in_frame[14] [5]), .I1(n46415), 
            .I2(GND_net), .I3(GND_net), .O(n46426));
    defparam i1_2_lut_adj_1099.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1100 (.I0(\data_in_frame[19] [0]), .I1(n46426), 
            .I2(n28010), .I3(\data_in_frame[16] [6]), .O(n49266));
    defparam i3_4_lut_adj_1100.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1101 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27549));   // verilog/coms.v(74[16:34])
    defparam i1_2_lut_adj_1101.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n2_adj_4712), .S(n3_adj_4713));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n2_adj_4714), .S(n3_adj_4715));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15491_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48658), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n29567));
    defparam i15491_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n29374));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1102 (.I0(n26308), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n27822));
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1103 (.I0(\data_in_frame[2] [6]), .I1(n28335), 
            .I2(\data_in_frame[5] [1]), .I3(GND_net), .O(n48811));
    defparam i1_3_lut_adj_1103.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1104 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n49204));   // verilog/coms.v(86[17:70])
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n29373));   // verilog/coms.v(128[12] 303[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk16MHz), 
            .E(n28649), .D(n9046[2]), .R(n29210));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_3_lut (.I0(n46389), .I1(\data_in_frame[22] [0]), .I2(n48992), 
            .I3(GND_net), .O(n8_adj_4716));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n28649), .D(n9046[3]), .R(n29210));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15492_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48658), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n29568));
    defparam i15492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n28649), .D(n9046[4]), .R(n29210));   // verilog/coms.v(128[12] 303[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk16MHz), 
            .E(n28649), .D(n9046[5]), .R(n29210));   // verilog/coms.v(128[12] 303[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk16MHz), 
            .E(n28649), .D(n9046[6]), .R(n29210));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n29372));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1105 (.I0(n52258), .I1(n48942), .I2(n48986), 
            .I3(\data_in_frame[23] [2]), .O(n52260));   // verilog/coms.v(269[9:85])
    defparam i1_4_lut_adj_1105.LUT_INIT = 16'hbeeb;
    SB_LUT4 i1_4_lut_adj_1106 (.I0(\data_in_frame[21] [6]), .I1(n52260), 
            .I2(n8_adj_4716), .I3(\data_in_frame[19] [6]), .O(n52262));   // verilog/coms.v(269[9:85])
    defparam i1_4_lut_adj_1106.LUT_INIT = 16'hdeed;
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n29371));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1107 (.I0(\data_in_frame[21] [5]), .I1(n49127), 
            .I2(n48681), .I3(\data_in_frame[23] [6]), .O(n50588));
    defparam i3_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n29370));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n29369));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n29368));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i4_4_lut_adj_1108 (.I0(\data_in_frame[23] [7]), .I1(n56717), 
            .I2(n46389), .I3(n6_adj_4699), .O(n50811));   // verilog/coms.v(86[17:28])
    defparam i4_4_lut_adj_1108.LUT_INIT = 16'h9669;
    SB_DFF data_in_0___i8 (.Q(\data_in[0]_c [7]), .C(clk16MHz), .D(n29367));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n29366));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1][1] ), .C(clk16MHz), .D(n29365));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1][2] ), .C(clk16MHz), .D(n29364));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1][3] ), .C(clk16MHz), .D(n29363));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n29362));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n29361));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1109 (.I0(n49204), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[7] [3]), .O(n52360));   // verilog/coms.v(72[16:69])
    defparam i1_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1110 (.I0(n48811), .I1(n27822), .I2(Kp_23__N_1098), 
            .I3(n52360), .O(n45470));   // verilog/coms.v(72[16:69])
    defparam i1_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(n27913), .I1(n45470), .I2(GND_net), 
            .I3(GND_net), .O(n46436));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i15 (.Q(\data_in[1][6] ), .C(clk16MHz), .D(n29360));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15493_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48658), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n29569));
    defparam i15493_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1112 (.I0(n52666), .I1(n52672), .I2(\data_in_frame[19] [1]), 
            .I3(n45510), .O(n50405));
    defparam i1_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1113 (.I0(n28051), .I1(n49230), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[4] [3]), .O(Kp_23__N_1206));   // verilog/coms.v(74[16:42])
    defparam i1_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i16 (.Q(\data_in[1]_c [7]), .C(clk16MHz), .D(n29359));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2][0] ), .C(clk16MHz), .D(n29358));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2][1] ), .C(clk16MHz), .D(n29356));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n29355));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2][3] ), .C(clk16MHz), .D(n29354));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_40730 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n56566));
    defparam byte_transmit_counter_0__bdd_4_lut_40730.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1114 (.I0(n49007), .I1(n49173), .I2(\data_in_frame[19] [6]), 
            .I3(\data_in_frame[22] [2]), .O(n52436));
    defparam i1_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1115 (.I0(\data_in_frame[21] [0]), .I1(\data_in_frame[22] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n52328));
    defparam i1_2_lut_adj_1115.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1116 (.I0(n49266), .I1(n27961), .I2(n52328), 
            .I3(\data_in_frame[20] [5]), .O(n52334));
    defparam i1_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i15494_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48658), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n29570));
    defparam i15494_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1117 (.I0(\data_in_frame[20] [2]), .I1(\data_in_frame[20] [1]), 
            .I2(\data_in_frame[22] [3]), .I3(\data_in_frame[19] [7]), .O(n52450));
    defparam i1_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1118 (.I0(n50405), .I1(n50811), .I2(n50588), 
            .I3(n52262), .O(n52268));   // verilog/coms.v(269[9:85])
    defparam i1_4_lut_adj_1118.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1119 (.I0(Kp_23__N_1206), .I1(n27590), .I2(\data_in_frame[6] [4]), 
            .I3(\data_in_frame[8] [6]), .O(n28032));   // verilog/coms.v(77[16:43])
    defparam i1_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i15495_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48658), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n29571));
    defparam i15495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_in_frame[8] [7]), .I1(n28032), 
            .I2(GND_net), .I3(GND_net), .O(n28477));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1121 (.I0(n49296), .I1(n46448), .I2(n52436), 
            .I3(n51116), .O(n52442));
    defparam i1_4_lut_adj_1121.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1122 (.I0(n50005), .I1(n48960), .I2(n52450), 
            .I3(GND_net), .O(n52454));
    defparam i1_3_lut_adj_1122.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_in_frame[8] [1]), .I1(Kp_23__N_1324), 
            .I2(GND_net), .I3(GND_net), .O(n49207));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1124 (.I0(n52454), .I1(n52442), .I2(n52268), 
            .I3(n49045), .O(n52272));   // verilog/coms.v(269[9:85])
    defparam i1_4_lut_adj_1124.LUT_INIT = 16'hf7fe;
    SB_LUT4 i1_4_lut_adj_1125 (.I0(n49336), .I1(n46363), .I2(n48960), 
            .I3(n52334), .O(n50889));
    defparam i1_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n29353));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1126 (.I0(n48942), .I1(n52272), .I2(n45486), 
            .I3(\data_in_frame[23] [0]), .O(n52274));   // verilog/coms.v(269[9:85])
    defparam i1_4_lut_adj_1126.LUT_INIT = 16'hedde;
    SB_LUT4 i1_4_lut_adj_1127 (.I0(n52274), .I1(\data_in_frame[23] [1]), 
            .I2(n50889), .I3(n45486), .O(n31_adj_4679));   // verilog/coms.v(269[9:85])
    defparam i1_4_lut_adj_1127.LUT_INIT = 16'hefbf;
    SB_LUT4 i15480_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48658), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n29556));
    defparam i15480_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(n27916), .I1(n27946), .I2(GND_net), 
            .I3(GND_net), .O(n28295));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1129 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[9] [2]), .I3(\data_in_frame[8] [3]), .O(n52580));
    defparam i1_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1130 (.I0(n49245), .I1(n52580), .I2(\data_in_frame[9] [1]), 
            .I3(\data_in_frame[8] [2]), .O(n52584));
    defparam i1_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i37127_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52919));
    defparam i37127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37128_3_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52920));
    defparam i37128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15481_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48658), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n29557));
    defparam i15481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i22 (.Q(\data_in[2][5] ), .C(clk16MHz), .D(n29352));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2][6] ), .C(clk16MHz), .D(n29351));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2]_c [7]), .C(clk16MHz), .D(n35692));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n29349));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3]_c [1]), .C(clk16MHz), .D(n29348));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n29347));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3][3] ), .C(clk16MHz), .D(n29346));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n29345));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3][5] ), .C(clk16MHz), .D(n35686));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3][6] ), .C(clk16MHz), .D(n29343));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3]_c [7]), .C(clk16MHz), .D(n35689));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
           .D(n29341));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
           .D(n29340));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
           .D(n29339));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
           .D(n29338));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
           .D(n29337));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
           .D(n29336));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
           .D(n29335));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
           .D(n29334));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
           .D(n29333));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
           .D(n29332));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
           .D(n29331));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
           .D(n29330));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
           .D(n29329));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
           .D(n29328));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
           .D(n29327));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1131 (.I0(n28105), .I1(n49207), .I2(n48817), 
            .I3(n52584), .O(n52590));
    defparam i1_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
           .D(n29326));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
           .D(n29325));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
           .D(n29323));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1132 (.I0(n28477), .I1(n52590), .I2(\data_in_frame[12] [0]), 
            .I3(n45442), .O(n49257));
    defparam i1_4_lut_adj_1132.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
           .D(n29322));   // verilog/coms.v(128[12] 303[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk16MHz), 
            .E(n28649), .D(n9046[7]), .R(n29210));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56566_bdd_4_lut (.I0(n56566), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n56569));
    defparam n56566_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_40725 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n56560));
    defparam byte_transmit_counter_0__bdd_4_lut_40725.LUT_INIT = 16'he4aa;
    SB_LUT4 n56560_bdd_4_lut (.I0(n56560), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n56563));
    defparam n56560_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n28717), .D(n48773));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37212_3_lut (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53004));
    defparam i37212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37211_3_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[21] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53003));
    defparam i37211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1133 (.I0(n49358), .I1(n49406), .I2(n49333), 
            .I3(GND_net), .O(n49045));
    defparam i1_3_lut_adj_1133.LUT_INIT = 16'h9696;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n28717), .D(n50782));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n28717), .D(n50686));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n28717), .D(n50306));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n28717), .D(n50411));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n28717), .D(n50065));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15482_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48658), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n29558));
    defparam i15482_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37103_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52895));
    defparam i37103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37104_3_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52896));
    defparam i37104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15483_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48658), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n29559));
    defparam i15483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n28717), .D(n50541));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n28717), .D(n50073));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n28717), .D(n50544));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n28717), .D(n50966));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n28717), .D(n49279));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1134 (.I0(\data_in_frame[11] [7]), .I1(n45470), 
            .I2(GND_net), .I3(GND_net), .O(n48945));
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1135 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27615));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_adj_1135.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1136 (.I0(n48945), .I1(n49198), .I2(\data_in_frame[14] [1]), 
            .I3(\data_in_frame[11] [5]), .O(n12_adj_4718));
    defparam i5_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n52913), .I2(n52914), .I3(byte_transmit_counter[2]), .O(n56530));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n56530_bdd_4_lut (.I0(n56530), .I1(n52908), .I2(n52907), .I3(byte_transmit_counter[2]), 
            .O(n56533));
    defparam n56530_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n28717), .D(n50662));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37254_3_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53046));
    defparam i37254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37253_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[21] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53045));
    defparam i37253_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n28717), .D(n50903));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i6_4_lut_adj_1137 (.I0(\data_in_frame[13] [7]), .I1(n12_adj_4718), 
            .I2(n49257), .I3(n28295), .O(n46444));
    defparam i6_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i15484_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48658), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n29560));
    defparam i15484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1138 (.I0(\data_in_frame[11] [5]), .I1(n46436), 
            .I2(\data_in_frame[9] [3]), .I3(n6_adj_4719), .O(Kp_23__N_1587));
    defparam i4_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\data_in_frame[12] [5]), .I1(n27669), 
            .I2(GND_net), .I3(GND_net), .O(n48820));
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n28717), .D(n50534));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15485_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48658), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n29561));
    defparam i15485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n52426));   // verilog/coms.v(264[5:27])
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_1141 (.I0(n27119), .I1(n31_adj_4679), .I2(n24561), 
            .I3(n52426), .O(n50602));   // verilog/coms.v(264[5:27])
    defparam i1_4_lut_adj_1141.LUT_INIT = 16'hfffe;
    SB_LUT4 i38620_2_lut (.I0(n56641), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54306));
    defparam i38620_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n28717), .D(n50504));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n28717), .D(n51075));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n2_adj_4720), .S(n3_adj_4721));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n2_adj_4722), .S(n3_adj_4723));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1142 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n48768));
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(\data_in_frame[12] [1]), .I1(n45569), 
            .I2(GND_net), .I3(GND_net), .O(n49093));
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1144 (.I0(n48971), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[12] [5]), .I3(\data_in_frame[12] [0]), .O(n52472));
    defparam i1_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1145 (.I0(n52472), .I1(n27608), .I2(n48736), 
            .I3(n49351), .O(n52478));
    defparam i1_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1146 (.I0(n48916), .I1(n48922), .I2(n52478), 
            .I3(n49157), .O(n52484));
    defparam i1_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1147 (.I0(n49170), .I1(n49093), .I2(n49260), 
            .I3(n52484), .O(n52490));
    defparam i1_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1148 (.I0(n46432), .I1(n49004), .I2(n45436), 
            .I3(n52490), .O(n46409));
    defparam i1_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1149 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n48728));
    defparam i1_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1150 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n48704));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49384));
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i21734_3_lut (.I0(n63_adj_4653), .I1(n63_c), .I2(\FRAME_MATCHER.state [2]), 
            .I3(GND_net), .O(n122));   // verilog/coms.v(140[4] 142[7])
    defparam i21734_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_751_Select_2_i5_4_lut (.I0(n122), .I1(\FRAME_MATCHER.i_31__N_2843 ), 
            .I2(n3303), .I3(n63), .O(n5));
    defparam select_751_Select_2_i5_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i15486_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48658), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n29562));
    defparam i15486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21730_rep_443_2_lut (.I0(n122), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n57092));   // verilog/coms.v(143[4] 145[7])
    defparam i21730_rep_443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15487_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48658), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n29563));
    defparam i15487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(n27556), .I1(n28047), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1130));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n2_adj_4725), .S(n3_adj_4726));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_adj_1153 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n27556));   // verilog/coms.v(167[9:87])
    defparam i1_3_lut_adj_1153.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1154 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n28051));   // verilog/coms.v(76[16:43])
    defparam i1_3_lut_adj_1154.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n2_adj_4727), .S(n3_adj_4728));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n2_adj_4729), .S(n3_adj_4730));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37089_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52881));
    defparam i37089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1155 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n52528));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1155.LUT_INIT = 16'h6666;
    SB_LUT4 i37090_4_lut (.I0(n52881), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n52882));
    defparam i37090_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i37088_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52880));
    defparam i37088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1156 (.I0(\data_in_frame[1] [7]), .I1(n49087), 
            .I2(n52528), .I3(\data_in_frame[0] [0]), .O(n27590));   // verilog/coms.v(75[16:43])
    defparam i1_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1157 (.I0(n28051), .I1(n27556), .I2(\data_in_frame[4] [4]), 
            .I3(GND_net), .O(n27506));   // verilog/coms.v(76[16:43])
    defparam i1_3_lut_adj_1157.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1158 (.I0(n27506), .I1(n27590), .I2(\data_in_frame[4] [5]), 
            .I3(\data_in_frame[6] [6]), .O(Kp_23__N_1324));   // verilog/coms.v(76[16:43])
    defparam i1_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1159 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[4] [5]), 
            .I2(\data_in_frame[7] [1]), .I3(GND_net), .O(n52552));   // verilog/coms.v(71[16:27])
    defparam i1_3_lut_adj_1159.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1160 (.I0(n49069), .I1(Kp_23__N_1130), .I2(n28335), 
            .I3(n52552), .O(n27913));   // verilog/coms.v(71[16:27])
    defparam i1_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_in_frame[9] [2]), .I1(n27913), 
            .I2(GND_net), .I3(GND_net), .O(n48922));   // verilog/coms.v(73[16:41])
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1162 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_1324), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4678));
    defparam i2_2_lut_adj_1162.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1163 (.I0(n7_adj_4678), .I1(n48922), .I2(\data_in_frame[9] [1]), 
            .I3(GND_net), .O(Kp_23__N_1536));   // verilog/coms.v(73[16:41])
    defparam i3_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1164 (.I0(\data_in_frame[13] [7]), .I1(n48728), 
            .I2(n46409), .I3(\data_in_frame[13] [1]), .O(n10_adj_4731));
    defparam i4_4_lut_adj_1164.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1165 (.I0(\data_in_frame[15] [7]), .I1(n10_adj_4731), 
            .I2(n27661), .I3(GND_net), .O(n48905));
    defparam i5_3_lut_adj_1165.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1166 (.I0(Kp_23__N_1587), .I1(\data_in_frame[16] [2]), 
            .I2(n46444), .I3(n27615), .O(n12_adj_4732));
    defparam i5_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1167 (.I0(n48905), .I1(n12_adj_4732), .I2(n49192), 
            .I3(\data_in_frame[16] [1]), .O(n45514));
    defparam i6_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1168 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n49173));
    defparam i1_2_lut_adj_1168.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(n45514), .I1(\data_in_frame[20] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n49007));
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n52544));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1171 (.I0(n48866), .I1(n49230), .I2(n52544), 
            .I3(\data_in_frame[0] [0]), .O(Kp_23__N_1203));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1172 (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_1203), 
            .I2(\data_in_frame[8] [4]), .I3(GND_net), .O(n49245));   // verilog/coms.v(75[16:43])
    defparam i1_3_lut_adj_1172.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1173 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n48866));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1173.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\data_in_frame[7] [7]), .I1(n48878), 
            .I2(GND_net), .I3(GND_net), .O(n28387));
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1175 (.I0(\data_in_frame[4] [0]), .I1(n48866), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[6] [1]), .O(n48710));   // verilog/coms.v(76[16:27])
    defparam i1_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1176 (.I0(n48710), .I1(n28387), .I2(\data_in_frame[10] [3]), 
            .I3(n49201), .O(n10_adj_4733));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1177 (.I0(\data_in_frame[8] [2]), .I1(n10_adj_4733), 
            .I2(\data_in_frame[8] [1]), .I3(GND_net), .O(n27669));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1178 (.I0(\data_in_frame[9] [5]), .I1(n27922), 
            .I2(\data_in_frame[9] [1]), .I3(Kp_23__N_1416), .O(n48731));
    defparam i3_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_in_frame[11] [1]), .I1(n28032), 
            .I2(GND_net), .I3(GND_net), .O(n48742));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(n48731), .I1(n49423), .I2(GND_net), 
            .I3(GND_net), .O(n49154));
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(n48896), .I1(n49245), .I2(GND_net), 
            .I3(GND_net), .O(n27601));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1182 (.I0(n49154), .I1(n45132), .I2(n48742), 
            .I3(n52080), .O(n50394));
    defparam i1_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1183 (.I0(n27669), .I1(n45522), .I2(GND_net), 
            .I3(GND_net), .O(n45571));
    defparam i1_2_lut_adj_1183.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1184 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[4] [0]), .I3(GND_net), .O(n49167));   // verilog/coms.v(79[16:27])
    defparam i1_3_lut_adj_1184.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1185 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[6] [2]), .O(n52700));   // verilog/coms.v(79[16:27])
    defparam i1_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1186 (.I0(\data_in_frame[15] [0]), .I1(n28353), 
            .I2(\data_in_frame[14] [7]), .I3(GND_net), .O(n49387));
    defparam i2_3_lut_adj_1186.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49284));
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(n4_adj_4669), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n48916));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1189 (.I0(n48896), .I1(n27583), .I2(\data_in_frame[8] [3]), 
            .I3(GND_net), .O(n28075));   // verilog/coms.v(74[16:42])
    defparam i1_3_lut_adj_1189.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_in_frame[11] [4]), .I1(Kp_23__N_1539), 
            .I2(GND_net), .I3(GND_net), .O(n27621));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1191 (.I0(n48974), .I1(n49084), .I2(n27615), 
            .I3(\data_in_frame[13] [5]), .O(n46500));
    defparam i1_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1192 (.I0(Kp_23__N_1206), .I1(Kp_23__N_1203), .I2(n27564), 
            .I3(\data_in_frame[8] [5]), .O(n28078));
    defparam i1_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1193 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n52300));
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1194 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[11] [4]), .O(n52314));
    defparam i1_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1195 (.I0(n28353), .I1(n49354), .I2(n28078), 
            .I3(n52314), .O(n52320));
    defparam i1_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1196 (.I0(n48967), .I1(n27969), .I2(n52300), 
            .I3(\data_in_frame[15] [1]), .O(n52306));
    defparam i1_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1197 (.I0(n49012), .I1(n46500), .I2(Kp_23__N_1539), 
            .I3(n52320), .O(n52326));
    defparam i1_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1198 (.I0(n45571), .I1(n52326), .I2(n52306), 
            .I3(n50394), .O(n46367));
    defparam i1_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
           .D(n29321));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40695 (.I0(byte_transmit_counter[1]), 
            .I1(n52898), .I2(n52899), .I3(byte_transmit_counter[2]), .O(n56494));
    defparam byte_transmit_counter_1__bdd_4_lut_40695.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n48919));
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1200 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n52344));
    defparam i1_2_lut_adj_1200.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1201 (.I0(n28328), .I1(n49189), .I2(n28468), 
            .I3(n52344), .O(n48925));
    defparam i1_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1202 (.I0(\data_in_frame[5] [4]), .I1(n28468), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n27445));
    defparam i1_3_lut_adj_1202.LUT_INIT = 16'h9696;
    SB_LUT4 n56494_bdd_4_lut (.I0(n56494), .I1(n52965), .I2(n52964), .I3(byte_transmit_counter[2]), 
            .O(n56497));
    defparam n56494_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15472_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48658), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n29548));
    defparam i15472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1203 (.I0(n27685), .I1(n27445), .I2(\data_in_frame[7] [6]), 
            .I3(GND_net), .O(n27649));
    defparam i1_3_lut_adj_1203.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1204 (.I0(n4_adj_4735), .I1(n48925), .I2(GND_net), 
            .I3(GND_net), .O(n27639));
    defparam i1_2_lut_adj_1204.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1416));   // verilog/coms.v(86[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n52458));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1206 (.I0(n48958), .I1(n49263), .I2(n27649), 
            .I3(n52458), .O(n45522));
    defparam i1_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n48971));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i15473_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48658), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n29549));
    defparam i15473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28129));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_LUT4 i15474_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48658), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n29550));
    defparam i15474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n27570));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1210 (.I0(n28129), .I1(n49201), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[1] [4]), .O(n28384));
    defparam i1_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1211 (.I0(n27570), .I1(n48817), .I2(n27515), 
            .I3(n28129), .O(n27552));   // verilog/coms.v(76[16:27])
    defparam i1_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4736));
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1213 (.I0(n27552), .I1(n45422), .I2(n28384), 
            .I3(n6_adj_4736), .O(n45569));
    defparam i4_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1214 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[16] [7]), 
            .I2(n49393), .I3(GND_net), .O(n49096));   // verilog/coms.v(79[16:27])
    defparam i2_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1215 (.I0(\data_in_frame[14] [4]), .I1(n48971), 
            .I2(n45436), .I3(n45522), .O(n28010));
    defparam i3_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(\data_in_frame[19] [2]), .I1(n46389), 
            .I2(GND_net), .I3(GND_net), .O(n48681));
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h9999;
    SB_LUT4 i37172_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52964));
    defparam i37172_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
           .D(n29957));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
           .D(n29956));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
           .D(n29955));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
           .D(n29954));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
           .D(n29953));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
           .D(n29952));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
           .D(n29951));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
           .D(n29950));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
           .D(n29949));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
           .D(n29948));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
           .D(n29947));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
           .D(n29946));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
           .D(n29945));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37173_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52965));
    defparam i37173_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
           .D(n29944));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
           .D(n29943));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
           .D(n29942));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
           .D(n29941));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
           .D(n29940));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
           .D(n29939));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
           .D(n29938));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
           .D(n29937));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
           .D(n29936));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
           .D(n29935));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
           .D(n29934));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
           .D(n29933));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
           .D(n29932));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_in_frame[21] [4]), .I1(n28010), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4737));
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
           .D(n29931));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i4_4_lut_adj_1218 (.I0(n46507), .I1(\data_in_frame[17] [1]), 
            .I2(n49096), .I3(n6_adj_4737), .O(n49127));
    defparam i4_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
           .D(n29930));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
           .D(n29929));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
           .D(n29928));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
           .D(n29927));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
           .D(n29926));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
           .D(n29925));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
           .D(n29924));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
           .D(n29923));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
           .D(n29922));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
           .D(n29921));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
           .D(n29920));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
           .D(n29919));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
           .D(n29918));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
           .D(n29917));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
           .D(n29916));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
           .D(n29915));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
           .D(n29914));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
           .D(n29913));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
           .D(n29912));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
           .D(n29911));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
           .D(n29910));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
           .D(n29909));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
           .D(n29908));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
           .D(n29907));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
           .D(n29906));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1219 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27515));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1219.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
           .D(n29905));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
           .D(n29904));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
           .D(n29903));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
           .D(n29902));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
           .D(n29901));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
           .D(n29900));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
           .D(n29899));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
           .D(n29898));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
           .D(n29897));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
           .D(n29896));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
           .D(n29895));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
           .D(n29894));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
           .D(n29893));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
           .D(n29892));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
           .D(n29891));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
           .D(n29890));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
           .D(n29889));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
           .D(n29888));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
           .D(n29887));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
           .D(n29886));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
           .D(n29885));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
           .D(n29884));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
           .D(n29883));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_4114_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n43271), .O(n9046[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4114_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n43270), .O(n9046[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_8 (.CI(n43270), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n43271));
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
           .D(n29882));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_4114_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n43269), .O(n9046[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_7 (.CI(n43269), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n43270));
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n28649), .D(n9046[0]), .R(n29210));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15475_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48658), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n29551));
    defparam i15475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n171), .D(n27278), 
            .R(n124));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15476_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48658), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n29552));
    defparam i15476_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n48644), .D(n29040), 
            .R(n49607));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40665 (.I0(byte_transmit_counter[1]), 
            .I1(n52922), .I2(n52923), .I3(byte_transmit_counter[2]), .O(n56488));
    defparam byte_transmit_counter_1__bdd_4_lut_40665.LUT_INIT = 16'he4aa;
    SB_LUT4 n56488_bdd_4_lut (.I0(n56488), .I1(n52956), .I2(n52955), .I3(byte_transmit_counter[2]), 
            .O(n56491));
    defparam n56488_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40660 (.I0(byte_transmit_counter[1]), 
            .I1(n52958), .I2(n52959), .I3(byte_transmit_counter[2]), .O(n56482));
    defparam byte_transmit_counter_1__bdd_4_lut_40660.LUT_INIT = 16'he4aa;
    SB_LUT4 n56482_bdd_4_lut (.I0(n56482), .I1(n52950), .I2(n52949), .I3(byte_transmit_counter[2]), 
            .O(n56485));
    defparam n56482_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40655 (.I0(byte_transmit_counter[1]), 
            .I1(n52934), .I2(n52935), .I3(byte_transmit_counter[2]), .O(n56476));
    defparam byte_transmit_counter_1__bdd_4_lut_40655.LUT_INIT = 16'he4aa;
    SB_LUT4 n56476_bdd_4_lut (.I0(n56476), .I1(n52929), .I2(n52928), .I3(byte_transmit_counter[2]), 
            .O(n56479));
    defparam n56476_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40650 (.I0(byte_transmit_counter[1]), 
            .I1(n53015), .I2(n53016), .I3(byte_transmit_counter[2]), .O(n56470));
    defparam byte_transmit_counter_1__bdd_4_lut_40650.LUT_INIT = 16'he4aa;
    SB_LUT4 n56470_bdd_4_lut (.I0(n56470), .I1(n52905), .I2(n52904), .I3(byte_transmit_counter[2]), 
            .O(n56473));
    defparam n56470_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
           .D(n29319));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
           .D(n29318));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
           .D(n29316));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
           .D(n29315));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
           .D(n29314));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
           .D(n29313));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
           .D(n29312));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
           .D(n29311));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
           .D(n29310));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
           .D(n29307));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
           .D(n29306));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
           .D(n29305));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
           .D(n29304));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
           .D(n29300));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
           .D(n29299));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
           .D(n29298));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
           .D(n29297));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
           .D(n29296));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
           .D(n29881));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15477_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48658), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n29553));
    defparam i15477_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15478_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48658), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n29554));
    defparam i15478_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15479_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48658), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n29555));
    defparam i15479_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1220 (.I0(n28078), .I1(n48731), .I2(GND_net), 
            .I3(GND_net), .O(n49151));
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1221 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[3] [3]), 
            .I2(\data_in_frame[5] [4]), .I3(\data_in_frame[7] [5]), .O(n52678));   // verilog/coms.v(86[17:63])
    defparam i1_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1222 (.I0(n48796), .I1(n49189), .I2(n52678), 
            .I3(GND_net), .O(n45422));   // verilog/coms.v(86[17:63])
    defparam i1_3_lut_adj_1222.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
           .D(n29880));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
           .D(n29879));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
           .D(n29878));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
           .D(n29877));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
           .D(n29876));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
           .D(n29875));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
           .D(n29874));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
           .D(n29873));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
           .D(n29872));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40645 (.I0(byte_transmit_counter[1]), 
            .I1(n52901), .I2(n52902), .I3(byte_transmit_counter[2]), .O(n56434));
    defparam byte_transmit_counter_1__bdd_4_lut_40645.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
           .D(n29871));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56434_bdd_4_lut (.I0(n56434), .I1(n53043), .I2(n53042), .I3(byte_transmit_counter[2]), 
            .O(n56437));
    defparam n56434_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
           .D(n29870));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_4114_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n43268), .O(n9046[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
           .D(n29869));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40616 (.I0(byte_transmit_counter[1]), 
            .I1(n52997), .I2(n52998), .I3(byte_transmit_counter[2]), .O(n56428));
    defparam byte_transmit_counter_1__bdd_4_lut_40616.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
           .D(n29868));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_4114_6 (.CI(n43268), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n43269));
    SB_LUT4 n56428_bdd_4_lut (.I0(n56428), .I1(n52917), .I2(n52916), .I3(byte_transmit_counter[2]), 
            .O(n56431));
    defparam n56428_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
           .D(n29867));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n29866));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40611 (.I0(byte_transmit_counter[1]), 
            .I1(n52982), .I2(n52983), .I3(byte_transmit_counter[2]), .O(n56422));
    defparam byte_transmit_counter_1__bdd_4_lut_40611.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n29865));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56422_bdd_4_lut (.I0(n56422), .I1(n52947), .I2(n52946), .I3(byte_transmit_counter[2]), 
            .O(n56425));
    defparam n56422_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n29864));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n29863));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40606 (.I0(byte_transmit_counter[1]), 
            .I1(n52943), .I2(n52944), .I3(byte_transmit_counter[2]), .O(n56416));
    defparam byte_transmit_counter_1__bdd_4_lut_40606.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n29862));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56416_bdd_4_lut (.I0(n56416), .I1(n52953), .I2(n52952), .I3(byte_transmit_counter[2]), 
            .O(n56419));
    defparam n56416_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29861));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n29860));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29859));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29858));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n29857));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n29856));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n29855));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n29854));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40601 (.I0(byte_transmit_counter[1]), 
            .I1(n52910), .I2(n52911), .I3(byte_transmit_counter[2]), .O(n56398));
    defparam byte_transmit_counter_1__bdd_4_lut_40601.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n29853));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56398_bdd_4_lut (.I0(n56398), .I1(n52962), .I2(n52961), .I3(byte_transmit_counter[2]), 
            .O(n56401));
    defparam n56398_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n29852));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29851));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
           .D(n29295));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n29850));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n29849));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 select_713_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4738));
    defparam select_713_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n29848));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n29847));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n29846));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n29845));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
           .D(n29294));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n29844));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
           .D(n29293));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n29843));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n29842));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n29841));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n29840));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i37107_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52899));
    defparam i37107_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
           .D(n29292));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_4_lut_adj_1223 (.I0(n49207), .I1(n52284), .I2(n28295), 
            .I3(Kp_23__N_1398), .O(n52288));
    defparam i1_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i37106_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52898));
    defparam i37106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_in_frame[16] [4]), .I1(n46475), 
            .I2(GND_net), .I3(GND_net), .O(n49305));
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1225 (.I0(n48933), .I1(n49263), .I2(n46436), 
            .I3(n52288), .O(n46432));
    defparam i1_4_lut_adj_1225.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
           .D(n29291));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
           .D(n29290));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
           .D(n29288));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
           .D(n29287));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
           .D(n29286));   // verilog/coms.v(128[12] 303[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk16MHz), 
           .D(n48016));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29284));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n29283));   // verilog/coms.v(128[12] 303[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n29282));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
           .D(n29281));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29280));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29279));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29278));   // verilog/coms.v(128[12] 303[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n29277));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n29276));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
           .D(n29275));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
           .D(n29274));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
           .D(n29273));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n29839));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n29838));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_4114_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n43267), .O(n9046[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n29837));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_4114_5 (.CI(n43267), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n43268));
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n29836));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_40759 (.I0(byte_transmit_counter[3]), 
            .I1(n56401), .I2(n54305), .I3(byte_transmit_counter[4]), .O(n56602));
    defparam byte_transmit_counter_3__bdd_4_lut_40759.LUT_INIT = 16'he4aa;
    SB_LUT4 add_4114_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n43266), .O(n9046[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n29835));   // verilog/coms.v(128[12] 303[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n29834));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1226 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [10]), .O(n48086));
    defparam i1_2_lut_4_lut_adj_1226.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_4_lut_adj_1227 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [11]), .O(n48084));
    defparam i1_2_lut_4_lut_adj_1227.LUT_INIT = 16'hec00;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40586 (.I0(byte_transmit_counter[1]), 
            .I1(n52883), .I2(n52884), .I3(byte_transmit_counter[2]), .O(n56386));
    defparam byte_transmit_counter_1__bdd_4_lut_40586.LUT_INIT = 16'he4aa;
    SB_LUT4 n56386_bdd_4_lut (.I0(n56386), .I1(n52974), .I2(n52973), .I3(byte_transmit_counter[2]), 
            .O(n56389));
    defparam n56386_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40576 (.I0(byte_transmit_counter[1]), 
            .I1(n52892), .I2(n52893), .I3(byte_transmit_counter[2]), .O(n56374));
    defparam byte_transmit_counter_1__bdd_4_lut_40576.LUT_INIT = 16'he4aa;
    SB_LUT4 n56374_bdd_4_lut (.I0(n56374), .I1(n52989), .I2(n52988), .I3(byte_transmit_counter[2]), 
            .O(n56377));
    defparam n56374_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_751_Select_1_i5_4_lut (.I0(n63), .I1(\FRAME_MATCHER.i_31__N_2843 ), 
            .I2(n3303), .I3(n92[1]), .O(n5_adj_4739));
    defparam select_751_Select_1_i5_4_lut.LUT_INIT = 16'hccc4;
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n28627), 
            .D(n7696));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n28627), 
            .D(n7695));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n28627), 
            .D(n7694));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n28627), 
            .D(n7693));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n28627), 
            .D(n7692));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n28627), 
            .D(n7691));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n28627), 
            .D(n7690));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_4114_4 (.CI(n43266), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n43267));
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n28627), 
            .D(n7689));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n28627), 
            .D(n7688));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1228 (.I0(n63_adj_6), .I1(n44910), .I2(n5_adj_4739), 
            .I3(n1_adj_4741), .O(n56701));
    defparam i3_4_lut_adj_1228.LUT_INIT = 16'hfffd;
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n28627), 
            .D(n7687));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n28627), 
            .D(n7686));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n28627), 
            .D(n7685));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n28627), 
            .D(n7684));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n28627), 
            .D(n7683));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n28627), .D(n7682));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n28627), .D(n7681));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n28627), .D(n7680));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n28627), .D(n7679));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n28627), .D(n7678));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n28627), .D(n7677));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n28627), .D(n7676));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n28627), .D(n7675));   // verilog/coms.v(128[12] 303[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n28627), .D(n7674));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk16MHz), 
            .D(n48110), .S(n48102));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1229 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [12]), .O(n48082));
    defparam i1_2_lut_4_lut_adj_1229.LUT_INIT = 16'hec00;
    SB_LUT4 add_4114_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n43265), .O(n9046[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4114_3 (.CI(n43265), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n43266));
    SB_LUT4 i1_2_lut_4_lut_adj_1230 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [13]), .O(n48080));
    defparam i1_2_lut_4_lut_adj_1230.LUT_INIT = 16'hec00;
    SB_LUT4 select_713_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4730));
    defparam select_713_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4728));
    defparam select_713_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4726));
    defparam select_713_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4114_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3748), .I3(GND_net), .O(n9046[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4114_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1231 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [14]), .O(n48078));
    defparam i1_2_lut_4_lut_adj_1231.LUT_INIT = 16'hec00;
    SB_CARRY add_4114_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3748), 
            .CO(n43265));
    SB_LUT4 add_43_33_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n43264), .O(n2_adj_4711)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n29833));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_32_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n43263), .O(n2_adj_4712)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_32 (.CI(n43263), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n43264));
    SB_LUT4 add_43_31_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n43262), .O(n2_adj_4714)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_31 (.CI(n43262), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n43263));
    SB_LUT4 add_43_30_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n43261), .O(n2_adj_4720)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_30 (.CI(n43261), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n43262));
    SB_LUT4 add_43_29_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n43260), .O(n2_adj_4722)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_29 (.CI(n43260), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n43261));
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n29832));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_28_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n43259), .O(n2_adj_4725)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_28 (.CI(n43259), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n43260));
    SB_LUT4 add_43_27_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n43258), .O(n2_adj_4727)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1232 (.I0(\FRAME_MATCHER.state [3]), .I1(n22902), 
            .I2(n4_adj_4742), .I3(n9), .O(n7_adj_4744));
    defparam i1_4_lut_adj_1232.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_4_lut_adj_1233 (.I0(n27119), .I1(n7_adj_4744), .I2(n27244), 
            .I3(\FRAME_MATCHER.state_31__N_2943 [3]), .O(n48114));
    defparam i1_4_lut_adj_1233.LUT_INIT = 16'hcdcc;
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n29831));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 select_713_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4723));
    defparam select_713_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4721));
    defparam select_713_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1234 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [15]), .O(n48076));
    defparam i1_2_lut_4_lut_adj_1234.LUT_INIT = 16'hec00;
    SB_LUT4 i5_4_lut_adj_1235 (.I0(n46498), .I1(n46440), .I2(\data_out_frame[25] [6]), 
            .I3(\data_out_frame[23] [6]), .O(n12_adj_4745));
    defparam i5_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1236 (.I0(\FRAME_MATCHER.state [3]), .I1(n22902), 
            .I2(n2_adj_4627), .I3(n4599), .O(n48012));
    defparam i1_4_lut_adj_1236.LUT_INIT = 16'ha8a0;
    SB_LUT4 i6_4_lut_adj_1237 (.I0(\data_out_frame[23] [4]), .I1(n12_adj_4745), 
            .I2(n49074), .I3(\data_out_frame[25] [7]), .O(n51075));
    defparam i6_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1238 (.I0(\FRAME_MATCHER.state [4]), .I1(n5_adj_4746), 
            .I2(GND_net), .I3(GND_net), .O(n48014));
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h8888;
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n29830));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i5_4_lut_adj_1239 (.I0(n46052), .I1(n48995), .I2(n45453), 
            .I3(n50908), .O(n12_adj_4747));
    defparam i5_4_lut_adj_1239.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1240 (.I0(n46477), .I1(n12_adj_4747), .I2(n49278), 
            .I3(\data_out_frame[25] [7]), .O(n50504));
    defparam i6_4_lut_adj_1240.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1241 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [16]), .O(n48074));
    defparam i1_2_lut_4_lut_adj_1241.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_adj_1242 (.I0(\FRAME_MATCHER.state [5]), .I1(n5_adj_4746), 
            .I2(GND_net), .I3(GND_net), .O(n48096));
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_1243 (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[21] [6]), 
            .I2(n49114), .I3(n6_adj_4748), .O(n50534));
    defparam i4_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n29829));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_27 (.CI(n43258), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n43259));
    SB_LUT4 add_43_26_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n43257), .O(n2_adj_4729)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i9_4_lut_adj_1244 (.I0(\data_out_frame[22] [1]), .I1(n49275), 
            .I2(n49375), .I3(n49217), .O(n22));
    defparam i9_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n29828));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\FRAME_MATCHER.state [6]), .I1(n5_adj_4746), 
            .I2(GND_net), .I3(GND_net), .O(n48094));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h8888;
    SB_LUT4 i7_3_lut (.I0(n51165), .I1(n49293), .I2(n45480), .I3(GND_net), 
            .O(n20_adj_4749));
    defparam i7_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i11_4_lut (.I0(n15_adj_4750), .I1(n22), .I2(n49269), .I3(n50160), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'h9669;
    SB_CARRY add_43_26 (.CI(n43257), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n43258));
    SB_LUT4 i12_4_lut (.I0(\data_out_frame[21] [6]), .I1(n24), .I2(n20_adj_4749), 
            .I3(\data_out_frame[19] [7]), .O(n46477));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
           .D(n29260));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1246 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [17]), .O(n48072));
    defparam i1_2_lut_4_lut_adj_1246.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\FRAME_MATCHER.state [7]), .I1(n5_adj_4746), 
            .I2(GND_net), .I3(GND_net), .O(n48092));
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_25_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n43256), .O(n2_adj_4751)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_25 (.CI(n43256), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n43257));
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\FRAME_MATCHER.state [8]), .I1(n5_adj_4746), 
            .I2(GND_net), .I3(GND_net), .O(n48090));
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_24_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n43255), .O(n2_adj_4752)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_24 (.CI(n43255), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n43256));
    SB_LUT4 add_43_23_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n43254), .O(n2_adj_4753)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_23 (.CI(n43254), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n43255));
    SB_LUT4 i37115_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52907));
    defparam i37115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37116_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52908));
    defparam i37116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37122_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52914));
    defparam i37122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_22_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n43253), .O(n2_adj_4754)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i37121_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52913));
    defparam i37121_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_22 (.CI(n43253), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n43254));
    SB_LUT4 add_43_21_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n43252), .O(n2_adj_4684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(\FRAME_MATCHER.state [9]), .I1(n5_adj_4746), 
            .I2(GND_net), .I3(GND_net), .O(n48088));
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h8888;
    SB_CARRY add_43_21 (.CI(n43252), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n43253));
    SB_LUT4 add_43_20_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n43251), .O(n2_adj_4685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n43251), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n43252));
    SB_LUT4 i1_2_lut_4_lut_adj_1250 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [18]), .O(n48018));
    defparam i1_2_lut_4_lut_adj_1250.LUT_INIT = 16'hec00;
    SB_LUT4 i5_4_lut_adj_1251 (.I0(n27448), .I1(n49020), .I2(n50561), 
            .I3(\data_out_frame[21] [7]), .O(n12_adj_4755));
    defparam i5_4_lut_adj_1251.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1252 (.I0(n51086), .I1(n12_adj_4755), .I2(n49118), 
            .I3(n50784), .O(n46456));
    defparam i6_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1253 (.I0(\data_out_frame[20] [2]), .I1(n51199), 
            .I2(\data_out_frame[20] [0]), .I3(GND_net), .O(n49118));
    defparam i2_3_lut_adj_1253.LUT_INIT = 16'h6969;
    SB_LUT4 add_43_19_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n43250), .O(n2_adj_4686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1254 (.I0(n50467), .I1(n49118), .I2(\data_out_frame[22] [3]), 
            .I3(GND_net), .O(n50101));
    defparam i2_3_lut_adj_1254.LUT_INIT = 16'h6969;
    SB_DFF deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29259));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n29827));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_out_frame[24] [5]), .I1(n46052), 
            .I2(GND_net), .I3(GND_net), .O(n49064));
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n29826));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1256 (.I0(\data_out_frame[25] [0]), .I1(n49287), 
            .I2(n49064), .I3(n49075), .O(n50544));
    defparam i3_4_lut_adj_1256.LUT_INIT = 16'h9669;
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n29825));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56590_bdd_4_lut (.I0(n56590), .I1(n56479), .I2(n7_adj_4756), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n56590_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15432_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48665), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n29508));
    defparam i15432_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n29824));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_19 (.CI(n43250), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n43251));
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n29823));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15433_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48665), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n29509));
    defparam i15433_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15434_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48665), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n29510));
    defparam i15434_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n29822));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n29821));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15435_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48665), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n29511));
    defparam i15435_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1257 (.I0(n2520), .I1(n49195), .I2(n48995), .I3(n49075), 
            .O(n50073));
    defparam i3_4_lut_adj_1257.LUT_INIT = 16'h9669;
    SB_LUT4 i15436_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48665), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n29512));
    defparam i15436_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n29820));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk16MHz), 
            .D(n48184), .S(n48048));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15437_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48665), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n29513));
    defparam i15437_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15438_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48665), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n29514));
    defparam i15438_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk16MHz), 
            .D(n48182), .S(n48050));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk16MHz), 
            .D(n48180), .S(n48052));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk16MHz), 
            .D(n48178), .S(n48054));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk16MHz), 
            .D(n48176), .S(n48056));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk16MHz), 
            .D(n48174), .S(n48058));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk16MHz), 
            .D(n48172), .S(n48060));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk16MHz), 
            .D(n48170), .S(n48062));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk16MHz), 
            .D(n48168), .S(n48064));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk16MHz), 
            .D(n48166), .S(n48066));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk16MHz), 
            .D(n48164), .S(n48068));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk16MHz), 
            .D(n48162), .S(n48070));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk16MHz), 
            .D(n48160), .S(n48018));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk16MHz), 
            .D(n48158), .S(n48072));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk16MHz), 
            .D(n48156), .S(n48074));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk16MHz), 
            .D(n48150), .S(n48076));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk16MHz), 
            .D(n48142), .S(n48078));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk16MHz), 
            .D(n48134), .S(n48080));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk16MHz), 
            .D(n48132), .S(n48082));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk16MHz), 
            .D(n48130), .S(n48084));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk16MHz), 
            .D(n48128), .S(n48086));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk16MHz), 
            .D(n48126), .S(n48088));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk16MHz), 
            .D(n48124), .S(n48090));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk16MHz), 
            .D(n48122), .S(n48092));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk16MHz), 
            .D(n48120), .S(n48094));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk16MHz), 
            .D(n48118), .S(n48096));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk16MHz), 
            .D(n48116), .S(n48014));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk16MHz), 
            .D(n48012), .S(n48114));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk16MHz), 
            .D(n48010), .S(n56701));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[24] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n48980));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n2_adj_4751), .S(n3_adj_4738));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15439_3_lut_4_lut (.I0(n8_adj_4625), .I1(n48665), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n29515));
    defparam i15439_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n2_adj_4752), .S(n3_adj_4663));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_18_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n43249), .O(n2_adj_4689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n2_adj_4753), .S(n3_adj_4662));   // verilog/coms.v(128[12] 303[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n2_adj_4754), .S(n3_adj_4659));   // verilog/coms.v(128[12] 303[6])
    SB_CARRY add_43_18 (.CI(n43249), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n43250));
    SB_LUT4 i4_4_lut_adj_1259 (.I0(n27421), .I1(n49026), .I2(\data_out_frame[22] [0]), 
            .I3(\data_out_frame[19] [6]), .O(n10_adj_4757));
    defparam i4_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_17_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n43248), .O(n2_adj_4690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_17 (.CI(n43248), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n43249));
    SB_LUT4 add_43_16_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n43247), .O(n2_adj_4703)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_16 (.CI(n43247), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n43248));
    SB_LUT4 add_43_15_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n43246), .O(n2_adj_4704)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1260 (.I0(\data_out_frame[22] [2]), .I1(n27905), 
            .I2(n49269), .I3(n48964), .O(n50467));
    defparam i3_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_CARRY add_43_15 (.CI(n43246), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n43247));
    SB_LUT4 add_43_14_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n43245), .O(n2_adj_4701)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_14 (.CI(n43245), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n43246));
    SB_LUT4 add_43_13_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n43244), .O(n2_adj_4700)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_13 (.CI(n43244), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n43245));
    SB_LUT4 add_43_12_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n43243), .O(n2_adj_4698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_12 (.CI(n43243), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n43244));
    SB_LUT4 add_43_11_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n43242), .O(n2_adj_4697)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15424_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48665), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n29500));
    defparam i15424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_11 (.CI(n43242), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n43243));
    SB_LUT4 add_43_10_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n43241), .O(n2_adj_4695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_10 (.CI(n43241), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n43242));
    SB_LUT4 add_43_9_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n43240), .O(n2_adj_4694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_9 (.CI(n43240), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n43241));
    SB_LUT4 i15425_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48665), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n29501));
    defparam i15425_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_8_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n43239), .O(n2_adj_4693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_8 (.CI(n43239), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n43240));
    SB_LUT4 add_43_7_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n43238), .O(n2_adj_4692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1261 (.I0(n51165), .I1(n50160), .I2(\data_out_frame[21] [5]), 
            .I3(n49061), .O(n49114));
    defparam i3_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_CARRY add_43_7 (.CI(n43238), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n43239));
    SB_LUT4 add_43_6_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n43237), .O(n2_adj_4688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15426_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48665), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n29502));
    defparam i15426_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15427_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48665), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n29503));
    defparam i15427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15428_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48665), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n29504));
    defparam i15428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\FRAME_MATCHER.state [14]), .I1(n4_adj_4758), 
            .I2(GND_net), .I3(GND_net), .O(n48142));
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(n46452), .I1(n49114), .I2(GND_net), 
            .I3(GND_net), .O(n49342));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1264 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [19]), .O(n48070));
    defparam i1_2_lut_4_lut_adj_1264.LUT_INIT = 16'hec00;
    SB_LUT4 i2_2_lut_adj_1265 (.I0(\data_out_frame[20] [6]), .I1(n46387), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4759));
    defparam i2_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1266 (.I0(n7_adj_4759), .I1(\data_out_frame[20] [7]), 
            .I2(n50467), .I3(\data_out_frame[22] [1]), .O(n49020));
    defparam i4_4_lut_adj_1266.LUT_INIT = 16'h9669;
    SB_CARRY add_43_6 (.CI(n43237), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n43238));
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
           .D(n29256));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n29819));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n29818));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n29817));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n29816));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n29815));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 add_43_5_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n43236), .O(n2_adj_4687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1267 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [20]), .O(n48068));
    defparam i1_2_lut_4_lut_adj_1267.LUT_INIT = 16'hec00;
    SB_LUT4 i15429_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48665), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n29505));
    defparam i15429_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_5 (.CI(n43236), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n43237));
    SB_LUT4 i15430_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48665), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n29506));
    defparam i15430_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15431_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48665), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n29507));
    defparam i15431_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_4_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n43235), .O(n2_adj_4683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_4 (.CI(n43235), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n43236));
    SB_LUT4 add_43_3_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n43234), .O(n2_adj_4681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_3_lut_adj_1268 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[19] [7]), 
            .I2(n49214), .I3(GND_net), .O(n8_adj_4760));
    defparam i3_3_lut_adj_1268.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4761));
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_CARRY add_43_3 (.CI(n43234), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n43235));
    SB_LUT4 add_43_2_lut (.I0(n3746), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_4_lut_adj_1270 (.I0(n28257), .I1(n4_adj_4761), .I2(n8_adj_4760), 
            .I3(n48823), .O(n48861));
    defparam i2_4_lut_adj_1270.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(\data_out_frame[19] [3]), .I1(n49130), 
            .I2(GND_net), .I3(GND_net), .O(n49061));
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n43234));
    SB_LUT4 i15416_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48665), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n29492));
    defparam i15416_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1272 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [21]), .O(n48066));
    defparam i1_2_lut_4_lut_adj_1272.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_adj_1273 (.I0(\FRAME_MATCHER.state [15]), .I1(n4_adj_4758), 
            .I2(GND_net), .I3(GND_net), .O(n48150));
    defparam i1_2_lut_adj_1273.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1274 (.I0(n50938), .I1(n48952), .I2(n28410), 
            .I3(GND_net), .O(n50160));
    defparam i2_3_lut_adj_1274.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[13] [0]), .I1(n27969), 
            .I2(\data_in_frame[12] [5]), .I3(n27669), .O(n28107));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15417_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48665), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n29493));
    defparam i15417_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1275 (.I0(\data_out_frame[21] [7]), .I1(n46504), 
            .I2(GND_net), .I3(GND_net), .O(n48707));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1275.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1276 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[3] [4]), .O(n48805));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i15418_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48665), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n29494));
    defparam i15418_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15419_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48665), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n29495));
    defparam i15419_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1277 (.I0(n45389), .I1(n48701), .I2(n49330), 
            .I3(n6_adj_4762), .O(n46387));
    defparam i4_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1278 (.I0(n51086), .I1(n49042), .I2(\data_out_frame[21] [6]), 
            .I3(n46387), .O(n50783));
    defparam i3_4_lut_adj_1278.LUT_INIT = 16'h9669;
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n29814));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n29813));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n29812));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i6_4_lut_adj_1279 (.I0(n50783), .I1(n28094), .I2(n48707), 
            .I3(n46452), .O(n14_adj_4763));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1279.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1280 (.I0(n45480), .I1(n46454), .I2(n49139), 
            .I3(n46440), .O(n13_adj_4764));   // verilog/coms.v(72[16:27])
    defparam i5_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n29811));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n29810));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n29809));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n29808));   // verilog/coms.v(128[12] 303[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n29807));   // verilog/coms.v(128[12] 303[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk16MHz), 
           .D(n56702));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i15420_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48665), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n29496));
    defparam i15420_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1281 (.I0(\FRAME_MATCHER.state [16]), .I1(n4_adj_4758), 
            .I2(GND_net), .I3(GND_net), .O(n48156));
    defparam i1_2_lut_adj_1281.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40567 (.I0(byte_transmit_counter[1]), 
            .I1(n53045), .I2(n53046), .I3(byte_transmit_counter[2]), .O(n56326));
    defparam byte_transmit_counter_1__bdd_4_lut_40567.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_adj_1282 (.I0(n13_adj_4764), .I1(n48861), .I2(n14_adj_4763), 
            .I3(GND_net), .O(n8_adj_4765));
    defparam i1_3_lut_adj_1282.LUT_INIT = 16'h9696;
    SB_LUT4 n56326_bdd_4_lut (.I0(n56326), .I1(n52896), .I2(n52895), .I3(byte_transmit_counter[2]), 
            .O(n56329));
    defparam n56326_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_40528 (.I0(byte_transmit_counter[1]), 
            .I1(n53003), .I2(n53004), .I3(byte_transmit_counter[2]), .O(n56320));
    defparam byte_transmit_counter_1__bdd_4_lut_40528.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_4_lut_adj_1283 (.I0(n49020), .I1(n49342), .I2(n45478), 
            .I3(n48955), .O(n12_adj_4766));
    defparam i5_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i15421_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48665), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n29497));
    defparam i15421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1284 (.I0(n46440), .I1(\data_out_frame[24] [7]), 
            .I2(\data_out_frame[23] [5]), .I3(\data_out_frame[23] [4]), 
            .O(n26));
    defparam i11_4_lut_adj_1284.LUT_INIT = 16'h9669;
    SB_LUT4 n56320_bdd_4_lut (.I0(n56320), .I1(n52920), .I2(n52919), .I3(byte_transmit_counter[2]), 
            .O(n56323));
    defparam n56320_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15422_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48665), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n29498));
    defparam i15422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15423_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48665), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n29499));
    defparam i15423_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n41963), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n27244), .O(\FRAME_MATCHER.i_31__N_2845 ));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i4_4_lut_adj_1285 (.I0(n27894), .I1(\data_out_frame[23] [7]), 
            .I2(n12_adj_4766), .I3(n8_adj_4765), .O(n19_adj_4767));
    defparam i4_4_lut_adj_1285.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1286 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(n41963), .I2(\FRAME_MATCHER.state[0] ), .I3(n27278), .O(\FRAME_MATCHER.i_31__N_2839 ));
    defparam i1_2_lut_3_lut_4_lut_adj_1286.LUT_INIT = 16'h1000;
    SB_LUT4 i36976_3_lut_4_lut (.I0(n4_adj_4735), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[0] [0]), .I3(Kp_23__N_1079), .O(n52716));
    defparam i36976_3_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i9_4_lut_adj_1287 (.I0(\data_out_frame[24] [5]), .I1(n48850), 
            .I2(n45604), .I3(\data_out_frame[24] [2]), .O(n24_adj_4768));
    defparam i9_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_LUT4 i15408_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48665), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29484));
    defparam i15408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut (.I0(n19_adj_4767), .I1(n26), .I2(n48980), .I3(\data_out_frame[23] [1]), 
            .O(n28));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15409_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48665), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29485));
    defparam i15409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_1288 (.I0(\data_out_frame[24] [6]), .I1(n28), 
            .I2(n24_adj_4768), .I3(n16_adj_4769), .O(n45453));
    defparam i14_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i15410_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48665), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n29486));
    defparam i15410_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15411_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48665), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29487));
    defparam i15411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15412_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48665), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29488));
    defparam i15412_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15413_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48665), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29489));
    defparam i15413_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15414_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48665), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29490));
    defparam i15414_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1289 (.I0(n45453), .I1(n49075), .I2(n45604), 
            .I3(\data_out_frame[24] [0]), .O(n50646));
    defparam i3_4_lut_adj_1289.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1290 (.I0(n27153), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n63_adj_6), .O(n29210));   // verilog/coms.v(213[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1290.LUT_INIT = 16'h00bf;
    SB_LUT4 i15415_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48665), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29491));
    defparam i15415_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1291 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [22]), .O(n48064));
    defparam i1_2_lut_4_lut_adj_1291.LUT_INIT = 16'hec00;
    SB_LUT4 i39853_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n11_adj_4702), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n171));   // verilog/coms.v(113[11:16])
    defparam i39853_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i4_4_lut_adj_1292 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[25] [1]), 
            .I2(n48755), .I3(n6_adj_4770), .O(n2520));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(n2520), .I1(n50646), .I2(GND_net), 
            .I3(GND_net), .O(n49287));
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h9999;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n56656));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1294 (.I0(n48989), .I1(n26792), .I2(n49019), 
            .I3(n49287), .O(n10_adj_4771));
    defparam i4_4_lut_adj_1294.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
           .D(n29762));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
           .D(n29761));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
           .D(n29760));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
           .D(n29759));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
           .D(n29758));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
           .D(n29757));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
           .D(n29756));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
           .D(n29755));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
           .D(n29754));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
           .D(n29753));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
           .D(n29752));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
           .D(n29751));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1295 (.I0(n45590), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[17] [7]), .I3(\data_out_frame[18] [0]), 
            .O(n49214));
    defparam i3_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1296 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[13] [4]), .I3(n26789), .O(n49375));
    defparam i3_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
           .D(n29726));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
           .D(n29725));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
           .D(n29724));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
           .D(n29723));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
           .D(n29722));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
           .D(n29721));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56656_bdd_4_lut (.I0(n56656), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n56659));
    defparam n56656_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
           .D(n29720));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
           .D(n29719));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
           .D(n29718));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
           .D(n29717));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
           .D(n29716));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1297 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [23]), .O(n48062));
    defparam i1_2_lut_4_lut_adj_1297.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1298 (.I0(n27916), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[9] [0]), .I3(\data_in_frame[11] [2]), .O(n49354));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
           .D(n29707));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
           .D(n29706));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
           .D(n29705));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
           .D(n29704));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
           .D(n29703));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
           .D(n29702));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1299 (.I0(n49039), .I1(n49375), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4772));
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
           .D(n29701));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i4_4_lut_adj_1300 (.I0(n28318), .I1(n27985), .I2(n49214), 
            .I3(n6_adj_4772), .O(n51199));
    defparam i4_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1301 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [24]), .O(n48060));
    defparam i1_2_lut_4_lut_adj_1301.LUT_INIT = 16'hec00;
    SB_LUT4 n56602_bdd_4_lut (.I0(n56602), .I1(n56491), .I2(n7_adj_4773), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n56602_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
           .D(n29687));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
           .D(n29686));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
           .D(n29685));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29666));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29665));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29664));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29663));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29662));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1302 (.I0(n48896), .I1(n49245), .I2(n28078), 
            .I3(GND_net), .O(Kp_23__N_1398));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1302.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29661));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29660));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29659));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29658));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29657));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29656));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29655));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n29654));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n29653));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n29652));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n29651));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n29650));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n29649));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n29648));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n29646));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n29645));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n29644));   // verilog/coms.v(128[12] 303[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n29643));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
           .D(n29642));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
           .D(n29641));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
           .D(n29640));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
           .D(n29639));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
           .D(n29638));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
           .D(n29637));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
           .D(n29636));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
           .D(n29635));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
           .D(n29634));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk16MHz), 
           .D(n29633));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk16MHz), 
           .D(n29632));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
           .D(n29631));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
           .D(n29630));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
           .D(n29629));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
           .D(n29628));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
           .D(n29627));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
           .D(n29626));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
           .D(n29625));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
           .D(n29624));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
           .D(n29623));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
           .D(n29622));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
           .D(n29621));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
           .D(n29620));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk16MHz), 
           .D(n29619));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1303 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[3] [2]), .O(n28468));
    defparam i1_3_lut_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
           .D(n29618));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk16MHz), 
           .D(n29617));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk16MHz), 
           .D(n29616));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk16MHz), 
           .D(n29615));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk16MHz), 
           .D(n29614));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk16MHz), 
           .D(n29613));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk16MHz), 
           .D(n29612));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
           .D(n29611));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
           .D(n29610));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
           .D(n29609));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
           .D(n29608));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
           .D(n29607));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
           .D(n29606));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
           .D(n29605));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
           .D(n29604));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n29603));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n29602));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
           .D(n29601));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n29600));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n29599));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
           .D(n29598));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
           .D(n29597));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
           .D(n29596));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
           .D(n29595));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
           .D(n29594));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
           .D(n29593));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
           .D(n29592));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
           .D(n29591));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
           .D(n29590));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
           .D(n29589));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
           .D(n29588));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
           .D(n29587));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
           .D(n29586));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
           .D(n29585));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
           .D(n29584));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
           .D(n29583));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
           .D(n29582));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
           .D(n29581));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
           .D(n29580));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
           .D(n29579));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
           .D(n29578));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
           .D(n29577));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
           .D(n29576));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
           .D(n29575));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
           .D(n29574));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
           .D(n29573));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
           .D(n29572));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n29571));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n29570));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n29569));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n29568));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n29567));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n29566));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1304 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[11] [2]), .I3(GND_net), .O(n49157));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1304.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n29565));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_adj_1305 (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[25] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49195));
    defparam i1_2_lut_adj_1305.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n29564));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
           .D(n29563));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
           .D(n29562));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_3_lut_adj_1306 (.I0(n48802), .I1(n49195), .I2(n27894), 
            .I3(GND_net), .O(n50065));
    defparam i2_3_lut_adj_1306.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
           .D(n29561));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i6_4_lut_adj_1307 (.I0(\data_out_frame[18] [1]), .I1(n49180), 
            .I2(n28318), .I3(n49372), .O(n16_adj_4774));
    defparam i6_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
           .D(n29560));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
           .D(n29559));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
           .D(n29558));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n29557));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
           .D(n29556));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n29555));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n29554));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n29553));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n29552));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n29551));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n29550));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n29549));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n29548));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n29547));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n29546));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n29545));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n29544));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n29543));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n29542));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n29541));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n29540));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n29539));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n29538));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n29537));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n29536));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
           .D(n29535));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
           .D(n29534));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
           .D(n29533));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
           .D(n29532));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
           .D(n29531));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
           .D(n29530));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
           .D(n29529));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
           .D(n29528));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
           .D(n29527));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
           .D(n29526));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i7_4_lut_adj_1308 (.I0(n46395), .I1(n49315), .I2(n50720), 
            .I3(n49090), .O(n17_adj_4775));
    defparam i7_4_lut_adj_1308.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
           .D(n29525));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
           .D(n29524));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
           .D(n29523));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
           .D(n29522));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
           .D(n29521));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
           .D(n29520));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
           .D(n29519));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i9_4_lut_adj_1309 (.I0(n17_adj_4775), .I1(n46513), .I2(n16_adj_4774), 
            .I3(\data_out_frame[13] [5]), .O(n49039));
    defparam i9_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1310 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [25]), .O(n48058));
    defparam i1_2_lut_4_lut_adj_1310.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_3_lut_adj_1311 (.I0(\data_out_frame[23] [5]), .I1(n28094), 
            .I2(n46504), .I3(GND_net), .O(n49075));
    defparam i1_2_lut_3_lut_adj_1311.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(n1247), .I3(GND_net), .O(n10_adj_4776));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1312 (.I0(n46138), .I1(n49039), .I2(\data_out_frame[20] [3]), 
            .I3(GND_net), .O(n27448));
    defparam i2_3_lut_adj_1312.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1313 (.I0(n27448), .I1(n48955), .I2(GND_net), 
            .I3(GND_net), .O(n45604));
    defparam i1_2_lut_adj_1313.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1314 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [3]), .I3(\data_out_frame[4] [2]), .O(n49034));
    defparam i1_2_lut_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
           .D(n29518));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
           .D(n29517));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n29516));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
           .D(n29515));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
           .D(n29514));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
           .D(n29513));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n29512));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n29511));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
           .D(n29510));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n29509));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
           .D(n29508));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
           .D(n29507));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n29506));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n29505));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n29504));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n29503));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
           .D(n29502));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
           .D(n29501));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
           .D(n29500));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
           .D(n29499));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n29498));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n29497));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n29496));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n29495));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n29494));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n29493));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n29492));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n29491));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n29490));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n29489));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n29488));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n29487));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
           .D(n29486));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n29485));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
           .D(n29484));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
           .D(n29483));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
           .D(n29482));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n29481));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n29480));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n29479));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n29478));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n29477));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n29476));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n29475));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
           .D(n29474));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
           .D(n29473));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
           .D(n29472));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
           .D(n29471));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
           .D(n29470));   // verilog/coms.v(128[12] 303[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n29469));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n29468));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n29467));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n29466));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n29465));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n29464));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n29463));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i2_2_lut_3_lut_adj_1315 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [2]), .I3(GND_net), .O(n10_adj_4777));   // verilog/coms.v(75[16:27])
    defparam i2_2_lut_3_lut_adj_1315.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n29462));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n29461));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n29460));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n29459));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n29458));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1316 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[12] [2]), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n49220));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1316.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n29457));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1317 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[25] [7]), .I3(GND_net), .O(n6_adj_4770));
    defparam i1_2_lut_3_lut_adj_1317.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1318 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [26]), .O(n48056));
    defparam i1_2_lut_4_lut_adj_1318.LUT_INIT = 16'hec00;
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n29456));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n29455));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n29454));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n29453));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n29452));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n29451));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n29450));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n29449));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n29448));   // verilog/coms.v(128[12] 303[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n29447));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1319 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [6]), 
            .I2(n49019), .I3(GND_net), .O(n48773));
    defparam i1_2_lut_3_lut_adj_1319.LUT_INIT = 16'h6969;
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n29446));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1320 (.I0(\data_out_frame[24] [7]), .I1(n50784), 
            .I2(\data_out_frame[22] [6]), .I3(n45438), .O(n48989));
    defparam i3_4_lut_adj_1320.LUT_INIT = 16'h9669;
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n29445));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[23] [3]), .I1(n46454), .I2(n46498), 
            .I3(n10_adj_4778), .O(n50782));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n29442));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n29441));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n29440));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n29439));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1321 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n28275));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1321.LUT_INIT = 16'h9696;
    SB_DFF deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n29438));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n29437));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_40799 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n56650));
    defparam byte_transmit_counter_0__bdd_4_lut_40799.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1322 (.I0(n48802), .I1(n48989), .I2(\data_out_frame[25] [2]), 
            .I3(GND_net), .O(n50411));
    defparam i2_3_lut_adj_1322.LUT_INIT = 16'h9696;
    SB_DFF deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n29434));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 n56650_bdd_4_lut (.I0(n56650), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n56653));
    defparam n56650_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[4] [2]), .O(n28401));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n29433));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1323 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [3]), .I3(\data_out_frame[4] [1]), .O(n1247));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_DFF deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n29432));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n29431));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n29430));   // verilog/coms.v(128[12] 303[6])
    SB_DFF deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n29429));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i3_4_lut_adj_1324 (.I0(\data_out_frame[16] [0]), .I1(n45590), 
            .I2(\data_out_frame[16] [1]), .I3(n27905), .O(n49372));
    defparam i3_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1325 (.I0(n25317), .I1(n49372), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4779));
    defparam i2_2_lut_adj_1325.LUT_INIT = 16'h6666;
    SB_DFF deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n29428));   // verilog/coms.v(128[12] 303[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1326 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(n27916), .I3(n27946), .O(Kp_23__N_1539));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1327 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[6] [1]), .I3(\data_out_frame[6] [2]), .O(n48687));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1328 (.I0(n49186), .I1(n14_adj_4780), .I2(n10_adj_4779), 
            .I3(\data_out_frame[18] [2]), .O(n46138));
    defparam i7_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1329 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[4] [2]), .I3(GND_net), .O(n27347));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1329.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_3_lut_4_lut (.I0(n28078), .I1(n48731), .I2(\data_in_frame[9] [0]), 
            .I3(n7_adj_4678), .O(n49423));
    defparam i1_3_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1330 (.I0(n28289), .I1(\data_out_frame[18] [5]), 
            .I2(n27848), .I3(n49000), .O(n10_adj_4781));
    defparam i4_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1331 (.I0(\data_out_frame[16] [3]), .I1(n10_adj_4781), 
            .I2(n50826), .I3(GND_net), .O(n49293));
    defparam i5_3_lut_adj_1331.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1332 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[19] [5]), .I3(n6_adj_4782), .O(n50561));
    defparam i4_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1333 (.I0(\data_out_frame[16] [6]), .I1(n48858), 
            .I2(\data_out_frame[19] [2]), .I3(GND_net), .O(n28289));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1333.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1334 (.I0(n48690), .I1(\data_out_frame[9] [6]), 
            .I2(n10_adj_4783), .I3(n28140), .O(n45376));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i22518_3_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n27153), .I3(n27119), .O(n4623));   // verilog/coms.v(128[12] 303[6])
    defparam i22518_3_lut_4_lut_4_lut.LUT_INIT = 16'hf8e8;
    SB_LUT4 i3_4_lut_adj_1335 (.I0(n48823), .I1(n48853), .I2(\data_out_frame[17] [3]), 
            .I3(n27863), .O(n49226));
    defparam i3_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1336 (.I0(n92[1]), .I1(n63), .I2(n4599), 
            .I3(n4_adj_4626), .O(n48010));   // verilog/coms.v(143[4] 145[7])
    defparam i1_2_lut_3_lut_4_lut_adj_1336.LUT_INIT = 16'hbbb0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1337 (.I0(n92[1]), .I1(n63), .I2(\FRAME_MATCHER.i_31__N_2845 ), 
            .I3(n4452), .O(n44910));   // verilog/coms.v(143[4] 145[7])
    defparam i1_2_lut_3_lut_4_lut_adj_1337.LUT_INIT = 16'h00b0;
    SB_LUT4 i2_3_lut_4_lut_adj_1338 (.I0(\data_out_frame[21] [1]), .I1(n45584), 
            .I2(\data_out_frame[20] [7]), .I3(n50826), .O(n49302));
    defparam i2_3_lut_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1339 (.I0(n50561), .I1(\data_out_frame[20] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n45480));
    defparam i1_2_lut_adj_1339.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1340 (.I0(\data_out_frame[16] [6]), .I1(n48858), 
            .I2(n49327), .I3(GND_net), .O(n6_adj_4784));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_LUT4 i21687_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n27153), .I3(n161), .O(n35747));   // verilog/coms.v(128[12] 303[6])
    defparam i21687_2_lut_3_lut_4_lut.LUT_INIT = 16'h0700;
    SB_LUT4 i2_4_lut_adj_1341 (.I0(\data_out_frame[20] [4]), .I1(n45480), 
            .I2(\data_out_frame[20] [7]), .I3(n48834), .O(n8_adj_4785));
    defparam i2_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut (.I0(\data_out_frame[16] [4]), .I1(n27580), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4786));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1342 (.I0(\data_out_frame[16] [5]), .I1(n48858), 
            .I2(n49217), .I3(n48834), .O(n45584));
    defparam i2_3_lut_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1343 (.I0(n9_adj_4786), .I1(n49077), .I2(n8_adj_4785), 
            .I3(n49082), .O(n51086));
    defparam i5_4_lut_adj_1343.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1344 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [27]), .O(n48054));
    defparam i1_2_lut_4_lut_adj_1344.LUT_INIT = 16'hec00;
    SB_LUT4 i2_3_lut_adj_1345 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[19] [4]), .I3(GND_net), .O(n49275));
    defparam i2_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27863));
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1347 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n41963), .I3(GND_net), .O(n27153));   // verilog/coms.v(128[12] 303[6])
    defparam i1_2_lut_3_lut_adj_1347.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_1348 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27421));
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1349 (.I0(n28401), .I1(n49339), .I2(GND_net), 
            .I3(GND_net), .O(n49162));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1349.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1350 (.I0(\data_out_frame[16] [5]), .I1(n48858), 
            .I2(n46403), .I3(GND_net), .O(n48684));
    defparam i1_2_lut_3_lut_adj_1350.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1351 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [28]), .O(n48052));
    defparam i1_2_lut_4_lut_adj_1351.LUT_INIT = 16'hec00;
    SB_LUT4 i4_4_lut_adj_1352 (.I0(\data_out_frame[13] [1]), .I1(n49312), 
            .I2(n48746), .I3(\data_out_frame[8] [3]), .O(n10_adj_4787));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1353 (.I0(n48713), .I1(n48939), .I2(\data_out_frame[11] [1]), 
            .I3(\data_out_frame[13] [3]), .O(n12_adj_4788));
    defparam i5_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1354 (.I0(\data_out_frame[11] [2]), .I1(n12_adj_4788), 
            .I2(n49162), .I3(n28394), .O(n28318));
    defparam i6_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(n28318), .I1(n48823), .I2(GND_net), 
            .I3(GND_net), .O(n49210));
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1356 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n1191), .I3(n48725), .O(n1168));   // verilog/coms.v(74[16:34])
    defparam i2_3_lut_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1357 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[24] [1]), 
            .I2(\data_out_frame[21] [7]), .I3(n46504), .O(n6_adj_4748));
    defparam i1_2_lut_3_lut_4_lut_adj_1357.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1358 (.I0(n49145), .I1(n28401), .I2(\data_out_frame[8] [7]), 
            .I3(n49239), .O(n10_adj_4789));
    defparam i4_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1359 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(\data_out_frame[4] [7]), .O(n28140));   // verilog/coms.v(74[16:34])
    defparam i2_3_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1360 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [29]), .O(n48050));
    defparam i1_2_lut_4_lut_adj_1360.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_4_lut_adj_1361 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [30]), .O(n48048));
    defparam i1_2_lut_4_lut_adj_1361.LUT_INIT = 16'hec00;
    SB_LUT4 i6_3_lut_4_lut (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[7] [5]), .I3(\data_out_frame[5] [3]), .O(n17_adj_4790));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1362 (.I0(\data_out_frame[13] [4]), .I1(n26789), 
            .I2(GND_net), .I3(GND_net), .O(n27905));
    defparam i1_2_lut_adj_1362.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1363 (.I0(n27347), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[10] [5]), .O(n10_adj_4791));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1364 (.I0(\data_out_frame[11] [0]), .I1(n10_adj_4791), 
            .I2(\data_out_frame[12] [7]), .I3(GND_net), .O(n48746));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_adj_1364.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1365 (.I0(n49345), .I1(\data_out_frame[11] [0]), 
            .I2(n48890), .I3(\data_out_frame[9] [0]), .O(n14_adj_4792));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1366 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[9] [7]), .I3(\data_out_frame[9] [4]), .O(n48884));
    defparam i2_3_lut_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1367 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(n1168), .I3(\data_out_frame[7] [0]), .O(n28394));   // verilog/coms.v(86[17:28])
    defparam i2_2_lut_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1368 (.I0(\data_out_frame[13] [2]), .I1(n14_adj_4792), 
            .I2(n10_adj_4793), .I3(\data_out_frame[11] [1]), .O(n27985));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[11] [2]), .I3(\data_out_frame[11] [1]), 
            .O(n10_adj_4794));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1369 (.I0(\data_out_frame[11] [3]), .I1(n28394), 
            .I2(GND_net), .I3(GND_net), .O(n48739));
    defparam i1_2_lut_adj_1369.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1370 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[11] [6]), .I3(n4_adj_4795), .O(n48912));   // verilog/coms.v(86[17:28])
    defparam i2_3_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1371 (.I0(n27208), .I1(n48674), .I2(n4), 
            .I3(\FRAME_MATCHER.state [31]), .O(n48102));
    defparam i1_2_lut_4_lut_adj_1371.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_adj_1372 (.I0(\data_out_frame[13] [0]), .I1(n50938), 
            .I2(GND_net), .I3(GND_net), .O(n46610));
    defparam i1_2_lut_adj_1372.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1373 (.I0(n49082), .I1(n49327), .I2(n49293), 
            .I3(GND_net), .O(n6_adj_4782));
    defparam i1_2_lut_3_lut_adj_1373.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1374 (.I0(n27343), .I1(n46610), .I2(n27848), 
            .I3(\data_out_frame[14] [6]), .O(n28_adj_4796));
    defparam i12_4_lut_adj_1374.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1375 (.I0(n1182), .I1(n48739), .I2(n48841), 
            .I3(\data_out_frame[13] [6]), .O(n26_adj_4797));
    defparam i10_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1376 (.I0(\data_out_frame[14] [1]), .I1(n28398), 
            .I2(\data_out_frame[13] [7]), .I3(n27985), .O(n27));
    defparam i11_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1377 (.I0(\data_out_frame[14] [4]), .I1(n48690), 
            .I2(\data_out_frame[11] [5]), .I3(n48746), .O(n25));
    defparam i9_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1378 (.I0(n25), .I1(n27), .I2(n26_adj_4797), 
            .I3(n28_adj_4796), .O(n51207));
    defparam i15_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(n49082), .I1(n49327), .I2(\data_out_frame[18] [6]), 
            .I3(GND_net), .O(n49217));
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1380 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(\data_out_frame[6] [1]), .O(n49312));
    defparam i1_2_lut_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1381 (.I0(n48930), .I1(n49233), .I2(n51207), 
            .I3(n49378), .O(n16_adj_4798));
    defparam i6_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1382 (.I0(\data_out_frame[14] [2]), .I1(n27905), 
            .I2(n49251), .I3(n49108), .O(n17_adj_4799));
    defparam i7_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1383 (.I0(n17_adj_4799), .I1(n49210), .I2(n16_adj_4798), 
            .I3(n49079), .O(n51208));
    defparam i9_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1384 (.I0(\data_out_frame[15] [7]), .I1(n27421), 
            .I2(n51208), .I3(\data_out_frame[15] [6]), .O(n10_adj_4800));
    defparam i4_4_lut_adj_1384.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1385 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[7] [7]), .I3(\data_out_frame[7] [6]), .O(n49324));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1386 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(n49145), .O(n6_adj_4801));
    defparam i2_2_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1387 (.I0(\data_out_frame[21] [0]), .I1(n49111), 
            .I2(n48850), .I3(n46498), .O(n25447));
    defparam i2_3_lut_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1388 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n49315));
    defparam i1_2_lut_3_lut_adj_1388.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1389 (.I0(n49048), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[17] [7]), .I3(n49315), .O(n10_adj_4802));
    defparam i4_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1390 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [6]), 
            .I2(n46361), .I3(GND_net), .O(n6_adj_4803));
    defparam i1_2_lut_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_4_lut (.I0(n27208), .I1(n4_adj_4626), .I2(\FRAME_MATCHER.i_31__N_2845 ), 
            .I3(n4452), .O(n4_adj_4758));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h88a8;
    SB_LUT4 i3_4_lut_adj_1391 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[17] [6]), .I3(\data_out_frame[19] [7]), 
            .O(n48964));
    defparam i3_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1392 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n48701));
    defparam i1_2_lut_adj_1392.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1393 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[17] [1]), .I3(\data_out_frame[18] [0]), 
            .O(n28_adj_4804));
    defparam i12_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1394 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[17] [2]), 
            .I2(n48964), .I3(n50720), .O(n26_adj_4805));
    defparam i10_4_lut_adj_1394.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1395 (.I0(\data_out_frame[17] [0]), .I1(n48701), 
            .I2(n48977), .I3(\data_out_frame[17] [3]), .O(n27_adj_4806));
    defparam i11_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1396 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[16] [0]), 
            .I2(n49275), .I3(\data_out_frame[18] [1]), .O(n25_adj_4807));
    defparam i9_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1397 (.I0(\data_out_frame[7] [0]), .I1(n1168), 
            .I2(n4_adj_4795), .I3(n48930), .O(n25317));   // verilog/coms.v(86[17:70])
    defparam i2_3_lut_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_40754 (.I0(byte_transmit_counter[3]), 
            .I1(n56419), .I2(n54303), .I3(byte_transmit_counter[4]), .O(n56596));
    defparam byte_transmit_counter_3__bdd_4_lut_40754.LUT_INIT = 16'he4aa;
    SB_LUT4 i15_4_lut_adj_1398 (.I0(n25_adj_4807), .I1(n27_adj_4806), .I2(n26_adj_4805), 
            .I3(n28_adj_4804), .O(n49000));
    defparam i15_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1399 (.I0(n26997), .I1(\data_out_frame[11] [5]), 
            .I2(\data_out_frame[15] [7]), .I3(GND_net), .O(n46395));
    defparam i1_2_lut_3_lut_adj_1399.LUT_INIT = 16'h9696;
    SB_LUT4 i37083_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52875));
    defparam i37083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_2_lut_3_lut (.I0(n49026), .I1(n49226), .I2(n46520), .I3(GND_net), 
            .O(n13_adj_4808));
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1400 (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[22] [6]), 
            .I2(n51086), .I3(GND_net), .O(n45478));
    defparam i2_3_lut_adj_1400.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1401 (.I0(n49026), .I1(n49226), .I2(\data_out_frame[19] [5]), 
            .I3(GND_net), .O(n49077));
    defparam i1_2_lut_3_lut_adj_1401.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1402 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [3]), 
            .I2(n28381), .I3(\data_out_frame[20] [2]), .O(n27580));   // verilog/coms.v(79[16:27])
    defparam i3_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i37084_4_lut (.I0(n52875), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n52876));
    defparam i37084_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i5_3_lut_adj_1403 (.I0(n45584), .I1(n27580), .I2(\data_out_frame[20] [0]), 
            .I3(GND_net), .O(n14_adj_4809));
    defparam i5_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1404 (.I0(n49111), .I1(\data_out_frame[19] [2]), 
            .I2(n45478), .I3(n49000), .O(n15_adj_4810));
    defparam i6_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1405 (.I0(\data_out_frame[23] [0]), .I1(n15_adj_4810), 
            .I2(n13_adj_4808), .I3(n14_adj_4809), .O(n49121));
    defparam i1_4_lut_adj_1405.LUT_INIT = 16'h9669;
    SB_LUT4 i37082_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52874));
    defparam i37082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1406 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n48725));   // verilog/coms.v(72[16:62])
    defparam i1_2_lut_3_lut_adj_1406.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1407 (.I0(n49139), .I1(n49429), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4811));
    defparam i1_2_lut_adj_1407.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1408 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(n27985), .I3(n46391), .O(n49026));
    defparam i2_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1409 (.I0(n46395), .I1(n49121), .I2(n49348), 
            .I3(n6_adj_4811), .O(n45438));
    defparam i4_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1410 (.I0(\data_out_frame[25] [2]), .I1(\data_out_frame[25] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n48755));
    defparam i1_2_lut_adj_1410.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1411 (.I0(n49029), .I1(\data_in_frame[16] [4]), 
            .I2(n46475), .I3(n48749), .O(n49165));
    defparam i1_2_lut_3_lut_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1412 (.I0(n49183), .I1(n49366), .I2(n49082), 
            .I3(n46138), .O(n46520));
    defparam i1_2_lut_4_lut_adj_1412.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1413 (.I0(n49183), .I1(n49366), .I2(n49082), 
            .I3(n46361), .O(n49042));
    defparam i1_2_lut_4_lut_adj_1413.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1414 (.I0(\data_out_frame[13] [6]), .I1(n48789), 
            .I2(\data_out_frame[16] [2]), .I3(\data_out_frame[18] [3]), 
            .O(n49348));
    defparam i3_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1415 (.I0(\data_out_frame[20] [4]), .I1(n46520), 
            .I2(\data_out_frame[22] [5]), .I3(GND_net), .O(n48955));
    defparam i1_2_lut_3_lut_adj_1415.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1416 (.I0(\data_out_frame[20] [4]), .I1(n46520), 
            .I2(n49042), .I3(\data_out_frame[20] [5]), .O(n50784));
    defparam i2_3_lut_4_lut_adj_1416.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1417 (.I0(\data_out_frame[16] [3]), .I1(n49220), 
            .I2(n10_adj_4783), .I3(n28140), .O(n45389));
    defparam i1_2_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1418 (.I0(n46395), .I1(n49348), .I2(GND_net), 
            .I3(GND_net), .O(n49183));
    defparam i1_2_lut_adj_1418.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1419 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n48939));
    defparam i1_2_lut_adj_1419.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1420 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[19] [1]), 
            .I2(n49023), .I3(GND_net), .O(n46498));
    defparam i1_2_lut_3_lut_adj_1420.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1421 (.I0(\data_out_frame[11] [3]), .I1(n28143), 
            .I2(n6_adj_4801), .I3(n48939), .O(n49180));
    defparam i1_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1422 (.I0(n49180), .I1(\data_out_frame[13] [5]), 
            .I2(n48789), .I3(GND_net), .O(n45590));
    defparam i2_3_lut_adj_1422.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1423 (.I0(\data_out_frame[16] [1]), .I1(n45590), 
            .I2(GND_net), .I3(GND_net), .O(n49366));
    defparam i1_2_lut_adj_1423.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1424 (.I0(n45604), .I1(n49121), .I2(n25447), 
            .I3(n10_adj_4771), .O(n50541));
    defparam i5_3_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1425 (.I0(n48834), .I1(\data_out_frame[23] [1]), 
            .I2(n49048), .I3(\data_out_frame[22] [7]), .O(n49429));
    defparam i3_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1426 (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[13] [6]), 
            .I2(n49330), .I3(GND_net), .O(n7_adj_4812));
    defparam i2_2_lut_3_lut_adj_1426.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1427 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28381));
    defparam i1_2_lut_adj_1427.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1428 (.I0(n49302), .I1(n28381), .I2(\data_out_frame[23] [2]), 
            .I3(n49429), .O(n10_adj_4813));
    defparam i4_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1429 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n48977));
    defparam i1_2_lut_adj_1429.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1430 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n49142));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1430.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1431 (.I0(n27448), .I1(\data_out_frame[22] [4]), 
            .I2(n48861), .I3(GND_net), .O(n46052));
    defparam i1_2_lut_3_lut_adj_1431.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1432 (.I0(n48713), .I1(n49142), .I2(\data_out_frame[9] [2]), 
            .I3(GND_net), .O(n28143));
    defparam i2_3_lut_adj_1432.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1433 (.I0(\data_out_frame[9] [3]), .I1(n48713), 
            .I2(n49142), .I3(\data_out_frame[9] [2]), .O(n48930));
    defparam i1_2_lut_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1434 (.I0(n26792), .I1(\data_out_frame[25] [4]), 
            .I2(n25447), .I3(\data_out_frame[25] [3]), .O(n50686));
    defparam i2_3_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1435 (.I0(\data_out_frame[11] [4]), .I1(n25317), 
            .I2(GND_net), .I3(GND_net), .O(n48789));
    defparam i1_2_lut_adj_1435.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1436 (.I0(n46395), .I1(n49348), .I2(n10_adj_4813), 
            .I3(\data_out_frame[19] [0]), .O(n26792));
    defparam i5_3_lut_4_lut_adj_1436.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1437 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [1]), 
            .I2(n45590), .I3(GND_net), .O(n49048));
    defparam i1_2_lut_3_lut_adj_1437.LUT_INIT = 16'h9696;
    SB_LUT4 i15464_3_lut_4_lut (.I0(n10), .I1(n48645), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n29540));
    defparam i15464_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1438 (.I0(n27448), .I1(\data_out_frame[22] [4]), 
            .I2(\data_out_frame[20] [2]), .I3(n51199), .O(n27894));
    defparam i2_3_lut_4_lut_adj_1438.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1439 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27576));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1439.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1440 (.I0(\data_out_frame[14] [0]), .I1(n48912), 
            .I2(GND_net), .I3(GND_net), .O(n49251));
    defparam i1_2_lut_adj_1440.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1441 (.I0(\data_out_frame[9] [5]), .I1(n49251), 
            .I2(\data_out_frame[9] [4]), .I3(\data_out_frame[5] [2]), .O(n10_adj_4814));
    defparam i4_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1442 (.I0(n27448), .I1(n48955), .I2(n49121), 
            .I3(\data_out_frame[25] [1]), .O(n48802));
    defparam i1_2_lut_3_lut_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1443 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[7] [4]), 
            .I2(n10_adj_4814), .I3(\data_out_frame[5] [3]), .O(n49330));
    defparam i1_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1444 (.I0(\data_out_frame[13] [6]), .I1(n49330), 
            .I2(GND_net), .I3(GND_net), .O(n49186));
    defparam i1_2_lut_adj_1444.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1445 (.I0(n7_adj_4812), .I1(n27576), .I2(n49082), 
            .I3(n49369), .O(n46361));
    defparam i4_4_lut_adj_1445.LUT_INIT = 16'h9669;
    SB_LUT4 i15465_3_lut_4_lut (.I0(n10), .I1(n48645), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n29541));
    defparam i15465_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1446 (.I0(n26792), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[25] [3]), .I3(n45438), .O(n50306));
    defparam i2_3_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1447 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(n28318), .I3(n48823), .O(n15_adj_4750));
    defparam i2_2_lut_3_lut_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1448 (.I0(\data_out_frame[20] [6]), .I1(n46599), 
            .I2(n46403), .I3(n6_adj_4803), .O(n49111));
    defparam i4_4_lut_adj_1448.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_3_lut_4_lut (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4780));
    defparam i6_4_lut_3_lut_4_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1449 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n48850));
    defparam i1_2_lut_adj_1449.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1450 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(n10_adj_4802), .I3(n46513), .O(n50720));
    defparam i5_3_lut_4_lut_adj_1450.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(\data_out_frame[25] [4]), .I1(n25447), 
            .I2(GND_net), .I3(GND_net), .O(n48844));
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1452 (.I0(n48844), .I1(\data_out_frame[23] [4]), 
            .I2(\data_out_frame[25] [5]), .I3(n28094), .O(n10_adj_4778));
    defparam i4_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1453 (.I0(\data_out_frame[21] [0]), .I1(n49111), 
            .I2(\data_out_frame[20] [6]), .I3(\data_out_frame[20] [5]), 
            .O(n49139));
    defparam i1_2_lut_3_lut_4_lut_adj_1453.LUT_INIT = 16'h9669;
    SB_LUT4 i15466_3_lut_4_lut (.I0(n10), .I1(n48645), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n29542));
    defparam i15466_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1454 (.I0(\data_out_frame[15] [0]), .I1(n10_adj_4800), 
            .I2(\data_out_frame[15] [1]), .I3(\data_out_frame[15] [2]), 
            .O(n46513));
    defparam i5_3_lut_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1455 (.I0(n49082), .I1(n49327), .I2(\data_out_frame[11] [4]), 
            .I3(n25317), .O(n49369));
    defparam i1_2_lut_3_lut_4_lut_adj_1455.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1456 (.I0(\data_out_frame[14] [6]), .I1(n1519), 
            .I2(n1516), .I3(n27356), .O(n28410));
    defparam i3_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1457 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27711));
    defparam i1_2_lut_adj_1457.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1458 (.I0(\data_out_frame[10] [7]), .I1(n1247), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n49339));
    defparam i2_3_lut_adj_1458.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1459 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n27343));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1459.LUT_INIT = 16'h9696;
    SB_LUT4 i22408_1_lut_2_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n165), .O(n3746));   // verilog/coms.v(128[12] 303[6])
    defparam i22408_1_lut_2_lut_4_lut.LUT_INIT = 16'h0070;
    SB_LUT4 i2_2_lut_4_lut_adj_1460 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[4] [5]), .I3(n27343), .O(n10_adj_4793));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1461 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n48902));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1461.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1462 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n49108));
    defparam i1_2_lut_adj_1462.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1463 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[4] [5]), 
            .I2(n1168), .I3(\data_out_frame[5] [0]), .O(n48713));   // verilog/coms.v(86[17:70])
    defparam i3_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1464 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n49239));
    defparam i1_2_lut_adj_1464.LUT_INIT = 16'h6666;
    SB_LUT4 i394_2_lut (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1182));   // verilog/coms.v(76[16:27])
    defparam i394_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1465 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[8] [4]), .I3(GND_net), .O(n48890));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1465.LUT_INIT = 16'h9696;
    SB_LUT4 i16_4_lut_adj_1466 (.I0(n49242), .I1(n27891), .I2(\data_out_frame[7] [1]), 
            .I3(\data_out_frame[4] [6]), .O(n40_adj_4815));
    defparam i16_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1467 (.I0(n1247), .I1(n48725), .I2(\data_out_frame[9] [3]), 
            .I3(n49324), .O(n38));
    defparam i14_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1468 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[7] [0]), 
            .I2(n48890), .I3(\data_out_frame[7] [2]), .O(n39_adj_4816));
    defparam i15_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1469 (.I0(\data_out_frame[9] [1]), .I1(n1182), 
            .I2(n48884), .I3(n49239), .O(n37));
    defparam i13_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1470 (.I0(\data_out_frame[11] [3]), .I1(n28394), 
            .I2(n10_adj_4789), .I3(\data_out_frame[11] [2]), .O(n26789));
    defparam i5_3_lut_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1471 (.I0(n49034), .I1(\data_out_frame[6] [4]), 
            .I2(n48713), .I3(\data_out_frame[4] [7]), .O(n42_adj_4817));
    defparam i18_4_lut_adj_1471.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n37), .I1(n39_adj_4816), .I2(n38), .I3(n40_adj_4815), 
            .O(n46));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1472 (.I0(n48902), .I1(\data_out_frame[6] [6]), 
            .I2(n49312), .I3(\data_out_frame[5] [5]), .O(n41_adj_4818));
    defparam i17_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1473 (.I0(\data_out_frame[10] [5]), .I1(n41_adj_4818), 
            .I2(n46), .I3(n42_adj_4817), .O(n12_adj_4819));
    defparam i4_4_lut_adj_1473.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1474 (.I0(n49029), .I1(n49305), .I2(\data_in_frame[18] [4]), 
            .I3(n50466), .O(n49336));
    defparam i2_3_lut_4_lut_adj_1474.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1475 (.I0(\data_out_frame[10] [0]), .I1(n49108), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[10] [2]), 
            .O(n13_adj_4820));
    defparam i5_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1476 (.I0(n13_adj_4820), .I1(n49339), .I2(n12_adj_4819), 
            .I3(\data_out_frame[10] [1]), .O(n46355));
    defparam i7_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i15467_3_lut_4_lut (.I0(n10), .I1(n48645), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n29543));
    defparam i15467_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1477 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(n1168), .I3(GND_net), .O(n49145));   // verilog/coms.v(72[16:69])
    defparam i2_3_lut_adj_1477.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1478 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27356));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_adj_1478.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1479 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28398));
    defparam i1_2_lut_adj_1479.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1480 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(\data_out_frame[12] [2]), 
            .O(n14_adj_4821));
    defparam i6_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1481 (.I0(\data_out_frame[19] [4]), .I1(n49226), 
            .I2(\data_out_frame[21] [5]), .I3(n49061), .O(n46440));
    defparam i2_3_lut_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1482 (.I0(\data_out_frame[19] [4]), .I1(n49226), 
            .I2(n49077), .I3(n50160), .O(n46452));
    defparam i2_3_lut_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1483 (.I0(\data_out_frame[12] [1]), .I1(n14_adj_4821), 
            .I2(n10_adj_4794), .I3(n27356), .O(n48872));
    defparam i7_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1484 (.I0(\data_out_frame[12] [0]), .I1(n46355), 
            .I2(GND_net), .I3(GND_net), .O(n49233));
    defparam i1_2_lut_adj_1484.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1485 (.I0(\data_out_frame[9] [4]), .I1(n49145), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4822));
    defparam i1_2_lut_adj_1485.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1486 (.I0(n28140), .I1(\data_out_frame[9] [3]), 
            .I2(n48713), .I3(n6_adj_4822), .O(n26997));
    defparam i4_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1487 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[24] [1]), 
            .I2(\data_out_frame[23] [0]), .I3(GND_net), .O(n16_adj_4769));
    defparam i1_2_lut_3_lut_adj_1487.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1488 (.I0(n26997), .I1(\data_out_frame[11] [7]), 
            .I2(n49233), .I3(n48872), .O(n10_adj_4823));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1489 (.I0(\data_out_frame[11] [4]), .I1(n10_adj_4823), 
            .I2(\data_out_frame[11] [6]), .I3(GND_net), .O(n50291));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_adj_1489.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1490 (.I0(n46355), .I1(\data_out_frame[11] [6]), 
            .I2(n50291), .I3(\data_out_frame[13] [7]), .O(n18_adj_4824));
    defparam i7_4_lut_adj_1490.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(n22902), .I1(n4_adj_4626), .I2(\FRAME_MATCHER.i_31__N_2839 ), 
            .I3(n771), .O(n4_adj_4742));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h88a8;
    SB_LUT4 i5_3_lut_4_lut_adj_1491 (.I0(n28401), .I1(n49339), .I2(n10_adj_4787), 
            .I3(\data_out_frame[4] [0]), .O(n48823));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_4_lut_adj_1491.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1492 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(Kp_23__N_1098), .I3(\data_in_frame[3] [0]), .O(n28328));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_4_lut_adj_1492.LUT_INIT = 16'h6996;
    SB_LUT4 i15468_3_lut_4_lut (.I0(n10), .I1(n48645), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n29544));
    defparam i15468_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1493 (.I0(n48872), .I1(\data_out_frame[5] [4]), 
            .I2(n28140), .I3(n27711), .O(n19_adj_4825));
    defparam i8_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1494 (.I0(\data_out_frame[14] [1]), .I1(n19_adj_4825), 
            .I2(n17_adj_4790), .I3(n18_adj_4824), .O(n49082));
    defparam i1_4_lut_adj_1494.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1495 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[13] [0]), 
            .I2(n50938), .I3(GND_net), .O(n46391));
    defparam i1_2_lut_3_lut_adj_1495.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1496 (.I0(\data_out_frame[23] [3]), .I1(n46454), 
            .I2(\data_out_frame[23] [5]), .I3(n49074), .O(n49019));
    defparam i1_2_lut_3_lut_4_lut_adj_1496.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1497 (.I0(\data_out_frame[18] [5]), .I1(n45389), 
            .I2(GND_net), .I3(GND_net), .O(n48834));
    defparam i1_2_lut_adj_1497.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1498 (.I0(\data_out_frame[20] [7]), .I1(n50826), 
            .I2(GND_net), .I3(GND_net), .O(n46599));
    defparam i1_2_lut_adj_1498.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1499 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n105));   // verilog/coms.v(113[11:16])
    defparam i1_2_lut_adj_1499.LUT_INIT = 16'h8888;
    SB_LUT4 i39838_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27278));
    defparam i39838_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i15469_3_lut_4_lut (.I0(n10), .I1(n48645), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n29545));
    defparam i15469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1500 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n49254));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1500.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1501 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [4]), .I3(\data_out_frame[13] [6]), 
            .O(n49090));
    defparam i2_3_lut_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1502 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4795));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1502.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1503 (.I0(n27576), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[13] [6]), .I3(n49369), .O(n6_adj_4762));
    defparam i1_2_lut_4_lut_adj_1503.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1504 (.I0(\data_out_frame[12] [0]), .I1(n48884), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4826));   // verilog/coms.v(72[16:27])
    defparam i2_2_lut_adj_1504.LUT_INIT = 16'h6666;
    SB_LUT4 select_713_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4624));
    defparam select_713_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1505 (.I0(n771), .I1(n22902), .I2(\FRAME_MATCHER.i_31__N_2839 ), 
            .I3(n48674), .O(n5_adj_4746));   // verilog/coms.v(158[6] 160[9])
    defparam i1_2_lut_4_lut_adj_1505.LUT_INIT = 16'hff40;
    SB_LUT4 i6_4_lut_adj_1506 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[10] [0]), 
            .I2(n48912), .I3(\data_out_frame[7] [6]), .O(n14_adj_4827));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1507 (.I0(\data_out_frame[14] [2]), .I1(n14_adj_4827), 
            .I2(n10_adj_4826), .I3(n49254), .O(n49327));   // verilog/coms.v(72[16:27])
    defparam i7_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i15470_3_lut_4_lut (.I0(n10), .I1(n48645), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n29546));
    defparam i15470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_40794 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n56644));
    defparam byte_transmit_counter_0__bdd_4_lut_40794.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1508 (.I0(\data_out_frame[24] [2]), .I1(n46477), 
            .I2(n46456), .I3(\data_out_frame[24] [3]), .O(n50662));
    defparam i2_3_lut_4_lut_adj_1508.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1509 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[18] [6]), 
            .I2(n46403), .I3(n6_adj_4784), .O(n50826));
    defparam i4_4_lut_adj_1509.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1510 (.I0(\data_out_frame[24] [2]), .I1(n46477), 
            .I2(n50908), .I3(\data_out_frame[24] [1]), .O(n50903));
    defparam i2_3_lut_4_lut_adj_1510.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1511 (.I0(n28410), .I1(n48684), .I2(\data_out_frame[17] [0]), 
            .I3(\data_out_frame[16] [7]), .O(n50278));
    defparam i3_4_lut_adj_1511.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1512 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[15] [3]), .I3(GND_net), .O(n28257));
    defparam i1_2_lut_3_lut_adj_1512.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_4_lut_adj_1513 (.I0(n63), .I1(n771), .I2(n4_adj_4626), 
            .I3(\FRAME_MATCHER.i_31__N_2839 ), .O(n5_adj_7));   // verilog/coms.v(158[6] 160[9])
    defparam i1_4_lut_4_lut_adj_1513.LUT_INIT = 16'ha2a0;
    SB_LUT4 i2_3_lut_adj_1514 (.I0(\data_out_frame[21] [2]), .I1(n50278), 
            .I2(n50826), .I3(GND_net), .O(n49023));
    defparam i2_3_lut_adj_1514.LUT_INIT = 16'h9696;
    SB_LUT4 i15471_3_lut_4_lut (.I0(n10), .I1(n48645), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n29547));
    defparam i15471_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_751_Select_1_i1_3_lut_4_lut (.I0(n63), .I1(n771), .I2(\FRAME_MATCHER.i_31__N_2839 ), 
            .I3(n92[1]), .O(n1_adj_4741));   // verilog/coms.v(158[6] 160[9])
    defparam select_751_Select_1_i1_3_lut_4_lut.LUT_INIT = 16'hf0d0;
    SB_LUT4 i1_2_lut_4_lut_adj_1515 (.I0(n45422), .I1(n49151), .I2(\data_in_frame[9] [0]), 
            .I3(n46432), .O(n45442));
    defparam i1_2_lut_4_lut_adj_1515.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1516 (.I0(\data_out_frame[15] [2]), .I1(n46610), 
            .I2(\data_out_frame[15] [5]), .I3(n27421), .O(n49269));
    defparam i1_2_lut_4_lut_adj_1516.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1517 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[11] [7]), .I3(\data_out_frame[14] [3]), 
            .O(n49378));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1518 (.I0(\data_out_frame[17] [5]), .I1(n10_adj_4757), 
            .I2(n28318), .I3(n48823), .O(n51165));
    defparam i5_3_lut_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1519 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [4]), .I3(n27515), .O(n48796));   // verilog/coms.v(79[16:27])
    defparam i1_3_lut_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1520 (.I0(n49378), .I1(n49136), .I2(\data_out_frame[9] [5]), 
            .I3(n49412), .O(n10_adj_4783));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1521 (.I0(n45376), .I1(\data_out_frame[18] [7]), 
            .I2(n27848), .I3(GND_net), .O(n46403));
    defparam i2_3_lut_adj_1521.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1522 (.I0(n27894), .I1(n50646), .I2(n27448), 
            .I3(n48955), .O(n48995));
    defparam i2_3_lut_4_lut_adj_1522.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1523 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n49230));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_3_lut_adj_1523.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1524 (.I0(\data_in_frame[12] [3]), .I1(n45569), 
            .I2(n45424), .I3(n51116), .O(n49426));
    defparam i1_2_lut_3_lut_4_lut_adj_1524.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1525 (.I0(\data_in_frame[12] [3]), .I1(n45569), 
            .I2(n27669), .I3(\data_in_frame[12] [4]), .O(n46415));
    defparam i2_3_lut_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1526 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[24] [5]), 
            .I2(n46052), .I3(n50101), .O(n50966));
    defparam i2_3_lut_4_lut_adj_1526.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1527 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49136));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1527.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1528 (.I0(\data_in_frame[12] [3]), .I1(n45569), 
            .I2(n49272), .I3(GND_net), .O(n46507));
    defparam i1_2_lut_3_lut_adj_1528.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1529 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [6]), .I3(GND_net), .O(n6_adj_4829));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1529.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1530 (.I0(n49056), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [0]), .I3(n49324), .O(n10_adj_4830));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1531 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n4_adj_4735));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1531.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1532 (.I0(\data_in_frame[16] [3]), .I1(n46475), 
            .I2(n46444), .I3(GND_net), .O(n48749));
    defparam i1_3_lut_adj_1532.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_4_lut_adj_1533 (.I0(\data_in_frame[17] [1]), .I1(n46367), 
            .I2(n52170), .I3(n49426), .O(n49358));
    defparam i1_3_lut_4_lut_adj_1533.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1534 (.I0(\data_out_frame[10] [2]), .I1(n10_adj_4830), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n1516));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_adj_1534.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1535 (.I0(n63_adj_4653), .I1(n63_c), .I2(n63), 
            .I3(GND_net), .O(n27208));   // verilog/coms.v(140[4] 142[7])
    defparam i1_2_lut_3_lut_adj_1535.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1536 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n49242));   // verilog/coms.v(72[16:62])
    defparam i1_2_lut_adj_1536.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1537 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n49056));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1537.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1538 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49079));
    defparam i1_2_lut_adj_1538.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1539 (.I0(\data_in_frame[17] [1]), .I1(n46367), 
            .I2(n46507), .I3(\data_in_frame[19] [3]), .O(n45510));
    defparam i1_3_lut_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1540 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[24] [3]), 
            .I2(n49278), .I3(GND_net), .O(n49279));
    defparam i1_2_lut_3_lut_adj_1540.LUT_INIT = 16'h9696;
    SB_LUT4 i22118_2_lut_3_lut (.I0(n63_adj_4653), .I1(n63_c), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n92[1]));   // verilog/coms.v(140[4] 142[7])
    defparam i22118_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1541 (.I0(n48687), .I1(n49242), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4831));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1541.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1542 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[10] [3]), 
            .I2(n49136), .I3(n6_adj_4831), .O(n1519));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1543 (.I0(n1519), .I1(n48687), .I2(n49079), .I3(GND_net), 
            .O(n14_adj_4832));
    defparam i5_3_lut_adj_1543.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1544 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[12] [6]), .I3(n49133), .O(n15_adj_4833));
    defparam i6_4_lut_adj_1544.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1545 (.I0(n15_adj_4833), .I1(\data_out_frame[10] [5]), 
            .I2(n14_adj_4832), .I3(\data_out_frame[6] [3]), .O(n48853));
    defparam i8_4_lut_adj_1545.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1546 (.I0(\data_out_frame[14] [5]), .I1(n48838), 
            .I2(\data_out_frame[12] [4]), .I3(n1516), .O(n27848));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1546.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1547 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4834));
    defparam i1_2_lut_adj_1547.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1548 (.I0(n50467), .I1(n49118), .I2(\data_out_frame[22] [3]), 
            .I3(n46456), .O(n49278));
    defparam i1_2_lut_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1549 (.I0(\data_out_frame[21] [7]), .I1(n46452), 
            .I2(n49114), .I3(\data_out_frame[23] [7]), .O(n50908));
    defparam i2_3_lut_4_lut_adj_1549.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1550 (.I0(n27848), .I1(\data_out_frame[16] [7]), 
            .I2(n48853), .I3(n6_adj_4834), .O(n49130));
    defparam i4_4_lut_adj_1550.LUT_INIT = 16'h6996;
    SB_LUT4 n56644_bdd_4_lut (.I0(n56644), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n56647));
    defparam n56644_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1551 (.I0(n28107), .I1(n46500), .I2(\data_in_frame[9] [4]), 
            .I3(GND_net), .O(n6_adj_4719));
    defparam i1_2_lut_3_lut_adj_1551.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1552 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n49412));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1552.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1553 (.I0(\data_out_frame[6] [0]), .I1(n49412), 
            .I2(\data_out_frame[8] [1]), .I3(\data_out_frame[7] [5]), .O(n48841));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1554 (.I0(n28107), .I1(n46500), .I2(n27621), 
            .I3(\data_in_frame[14] [7]), .O(n49012));
    defparam i1_3_lut_4_lut_adj_1554.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1555 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(n52700), .I3(n49167), .O(n48896));   // verilog/coms.v(79[16:27])
    defparam i1_3_lut_4_lut_adj_1555.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1556 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(n27556), .I3(GND_net), .O(n10_adj_4673));   // verilog/coms.v(79[16:27])
    defparam i2_2_lut_3_lut_adj_1556.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1557 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n27922));   // verilog/coms.v(74[16:42])
    defparam i1_2_lut_3_lut_adj_1557.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1558 (.I0(\data_out_frame[12] [3]), .I1(n49223), 
            .I2(\data_out_frame[10] [2]), .I3(\data_out_frame[5] [3]), .O(n10_adj_4835));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1558.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1559 (.I0(n48841), .I1(n10_adj_4835), .I2(\data_out_frame[5] [7]), 
            .I3(GND_net), .O(n48838));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_adj_1559.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1560 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n48690));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1560.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1561 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49223));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1561.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53035), .I3(n53033), .O(n7_adj_4836));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n52870), .I3(n52868), .O(n7_adj_4837));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53026), .I3(n53024), .O(n7_adj_4838));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1562 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27891));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1562.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n52864), .I3(n52862), .O(n7_adj_4773));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n52876), .I3(n52874), .O(n7_adj_4756));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i6_4_lut_adj_1563 (.I0(n49220), .I1(n28275), .I2(\data_out_frame[10] [0]), 
            .I3(\data_out_frame[10] [1]), .O(n14_adj_4839));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1563.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1564 (.I0(\data_out_frame[14] [4]), .I1(n14_adj_4839), 
            .I2(n10_adj_4777), .I3(n48838), .O(n48858));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_40789 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n56638));
    defparam byte_transmit_counter_0__bdd_4_lut_40789.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_4_lut_adj_1565 (.I0(n4_adj_4669), .I1(\data_in_frame[8] [7]), 
            .I2(n28032), .I3(n28075), .O(n52284));
    defparam i1_3_lut_4_lut_adj_1565.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n52882), .I3(n52880), .O(n7));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n52891), .I3(n52889), .O(n7_adj_4668));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n53050), .I3(n53048), .O(n7_adj_4707));   // verilog/coms.v(107[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1566 (.I0(\data_in_frame[5] [3]), .I1(n26308), 
            .I2(\data_in_frame[2] [7]), .I3(GND_net), .O(n49189));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_3_lut_adj_1566.LUT_INIT = 16'h9696;
    SB_LUT4 i880_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1668));   // verilog/coms.v(86[17:28])
    defparam i880_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15456_3_lut_4_lut (.I0(n8), .I1(n48658), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n29532));
    defparam i15456_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(72[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1567 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49345));
    defparam i1_2_lut_adj_1567.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1568 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [31]), .O(n48110));
    defparam i1_2_lut_4_lut_adj_1568.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_adj_1569 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n49133));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1569.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1570 (.I0(n48799), .I1(n49192), .I2(n27615), 
            .I3(n45132), .O(n45384));   // verilog/coms.v(72[16:27])
    defparam i1_3_lut_4_lut_adj_1570.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1571 (.I0(n48799), .I1(n49192), .I2(n27631), 
            .I3(n49052), .O(n49318));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1572 (.I0(n49345), .I1(n1191), .I2(n49034), .I3(n1668), 
            .O(n14_adj_4840));
    defparam i6_4_lut_adj_1572.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1573 (.I0(\data_out_frame[8] [3]), .I1(n14_adj_4840), 
            .I2(n10_adj_4776), .I3(\data_out_frame[10] [4]), .O(n50938));
    defparam i7_4_lut_adj_1573.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1574 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[17] [2]), .I3(\data_out_frame[13] [0]), 
            .O(n48952));
    defparam i3_4_lut_adj_1574.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1575 (.I0(\data_out_frame[16] [7]), .I1(n48952), 
            .I2(n50938), .I3(GND_net), .O(n8_adj_4841));
    defparam i2_3_lut_adj_1575.LUT_INIT = 16'h9696;
    SB_LUT4 i15457_3_lut_4_lut (.I0(n8), .I1(n48658), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n29533));
    defparam i15457_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1576 (.I0(n28289), .I1(\data_out_frame[21] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4842));
    defparam i1_2_lut_adj_1576.LUT_INIT = 16'h6666;
    SB_LUT4 i15458_3_lut_4_lut (.I0(n8), .I1(n48658), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n29534));
    defparam i15458_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1577 (.I0(\data_out_frame[17] [0]), .I1(n7_adj_4842), 
            .I2(\data_out_frame[19] [3]), .I3(n8_adj_4841), .O(n46504));
    defparam i5_4_lut_adj_1577.LUT_INIT = 16'h6996;
    SB_LUT4 i15459_3_lut_4_lut (.I0(n8), .I1(n48658), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n29535));
    defparam i15459_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1578 (.I0(\data_out_frame[19] [1]), .I1(n49130), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4843));
    defparam i1_2_lut_adj_1578.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1579 (.I0(\data_out_frame[21] [3]), .I1(n28289), 
            .I2(n48684), .I3(n6_adj_4843), .O(n28094));
    defparam i4_4_lut_adj_1579.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1580 (.I0(n28094), .I1(n46504), .I2(GND_net), 
            .I3(GND_net), .O(n49074));
    defparam i1_2_lut_adj_1580.LUT_INIT = 16'h6666;
    SB_LUT4 n56638_bdd_4_lut (.I0(n56638), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n56641));
    defparam n56638_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15460_3_lut_4_lut (.I0(n8), .I1(n48658), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n29536));
    defparam i15460_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15461_3_lut_4_lut (.I0(n8), .I1(n48658), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n29537));
    defparam i15461_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1581 (.I0(n49023), .I1(n49302), .I2(\data_out_frame[19] [1]), 
            .I3(GND_net), .O(n46454));
    defparam i2_3_lut_adj_1581.LUT_INIT = 16'h9696;
    SB_LUT4 i15462_3_lut_4_lut (.I0(n8), .I1(n48658), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n29538));
    defparam i15462_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15463_3_lut_4_lut (.I0(n8), .I1(n48658), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n29539));
    defparam i15463_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1582 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[12] [4]), 
            .I2(n49387), .I3(n49397), .O(n49272));
    defparam i1_2_lut_4_lut_adj_1582.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1583 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[7] [7]), 
            .I2(n48878), .I3(GND_net), .O(n48817));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1583.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1584 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n48933), .I3(\data_in_frame[10] [0]), .O(n45436));
    defparam i1_2_lut_4_lut_adj_1584.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1585 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n48933), .I3(GND_net), .O(n28105));
    defparam i1_2_lut_3_lut_adj_1585.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1586 (.I0(n4_adj_4735), .I1(n48925), .I2(n27649), 
            .I3(GND_net), .O(n48933));
    defparam i1_2_lut_3_lut_adj_1586.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1587 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n27685));
    defparam i1_2_lut_3_lut_adj_1587.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1588 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27564));   // verilog/coms.v(86[17:28])
    defparam i1_2_lut_adj_1588.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1589 (.I0(n45988), .I1(n27552), .I2(GND_net), 
            .I3(GND_net), .O(n49263));
    defparam i1_2_lut_adj_1589.LUT_INIT = 16'h6666;
    SB_LUT4 i37243_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n53035));
    defparam i37243_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i37241_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53033));
    defparam i37241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22911133_i1_3_lut (.I0(n56617), .I1(n56293), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4844));
    defparam i22911133_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38671_2_lut (.I0(n56569), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54289));
    defparam i38671_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i38631_2_lut (.I0(n56653), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54302));
    defparam i38631_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i37077_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52869));
    defparam i37077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37078_4_lut (.I0(n52869), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n52870));
    defparam i37078_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i15448_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48658), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n29524));
    defparam i15448_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37076_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n52868));
    defparam i37076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1590 (.I0(n48896), .I1(n49245), .I2(n28075), 
            .I3(\data_in_frame[10] [5]), .O(n28353));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1590.LUT_INIT = 16'h6996;
    SB_LUT4 i15449_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48658), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n29525));
    defparam i15449_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n56323), .I2(n54300), .I3(byte_transmit_counter[4]), .O(n56626));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1591 (.I0(n51116), .I1(n45424), .I2(\data_in_frame[21] [7]), 
            .I3(GND_net), .O(n48992));
    defparam i1_2_lut_3_lut_adj_1591.LUT_INIT = 16'h6969;
    SB_LUT4 i15450_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48658), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n29526));
    defparam i15450_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i40487_2_lut_4_lut (.I0(n27278), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n11_adj_4702), .I3(\FRAME_MATCHER.state [3]), .O(n49607));
    defparam i40487_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i15451_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48658), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n29527));
    defparam i15451_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1592 (.I0(n27278), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n11_adj_4702), .I3(\FRAME_MATCHER.state [3]), .O(n28717));
    defparam i1_2_lut_4_lut_adj_1592.LUT_INIT = 16'h0200;
    SB_LUT4 i15552_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48649), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29628));
    defparam i15552_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15553_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48649), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n29629));
    defparam i15553_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15452_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48658), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n29528));
    defparam i15452_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15554_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48649), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29630));
    defparam i15554_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15555_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48649), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29631));
    defparam i15555_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37233_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53025));
    defparam i37233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37234_4_lut (.I0(n53025), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n53026));
    defparam i37234_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i37232_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n53024));
    defparam i37232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15556_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48649), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n29632));
    defparam i15556_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1593 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[12] [4]), 
            .I2(n49387), .I3(GND_net), .O(n48967));
    defparam i1_2_lut_3_lut_adj_1593.LUT_INIT = 16'h9696;
    SB_LUT4 i15557_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48649), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n29633));
    defparam i15557_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i38773_2_lut (.I0(n56575), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54300));
    defparam i38773_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15558_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48649), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n29634));
    defparam i15558_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15559_3_lut_4_lut (.I0(n8_adj_4710), .I1(n48649), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n29635));
    defparam i15559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1594 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n6_adj_4671));   // verilog/coms.v(167[9:87])
    defparam i1_2_lut_3_lut_adj_1594.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1595 (.I0(n28075), .I1(n4_adj_4669), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n27969));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1595.LUT_INIT = 16'h9696;
    SB_LUT4 i38625_2_lut (.I0(n56659), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n54303));
    defparam i38625_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1596 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n28335));   // verilog/coms.v(167[9:87])
    defparam i1_2_lut_3_lut_adj_1596.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1597 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(n48710), .I3(Kp_23__N_1174), .O(n27583));   // verilog/coms.v(79[16:27])
    defparam i1_3_lut_4_lut_adj_1597.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1598 (.I0(n31), .I1(n24561), .I2(n105), 
            .I3(n27119), .O(n50620));
    defparam i2_3_lut_4_lut_adj_1598.LUT_INIT = 16'hffef;
    SB_LUT4 i2112_2_lut_3_lut (.I0(n31), .I1(n24561), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n7672));
    defparam i2112_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i15453_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48658), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n29529));
    defparam i15453_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1599 (.I0(n48896), .I1(n49245), .I2(\data_in_frame[11] [0]), 
            .I3(\data_in_frame[10] [6]), .O(n52080));
    defparam i1_3_lut_4_lut_adj_1599.LUT_INIT = 16'h6996;
    SB_LUT4 i15544_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48649), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29620));
    defparam i15544_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15545_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48649), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n29621));
    defparam i15545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15546_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48649), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n29622));
    defparam i15546_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15454_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48658), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n29530));
    defparam i15454_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15547_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48649), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n29623));
    defparam i15547_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15548_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48649), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n29624));
    defparam i15548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1600 (.I0(\data_in_frame[11] [1]), .I1(n28032), 
            .I2(n46429), .I3(n49354), .O(n45132));   // verilog/coms.v(72[16:27])
    defparam i1_3_lut_4_lut_adj_1600.LUT_INIT = 16'h9669;
    SB_LUT4 i15455_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48658), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n29531));
    defparam i15455_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1601 (.I0(n22902), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [4]), .O(n48116));
    defparam i1_2_lut_4_lut_adj_1601.LUT_INIT = 16'hf800;
    SB_LUT4 i15549_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48649), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n29625));
    defparam i15549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15550_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48649), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n29626));
    defparam i15550_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15551_3_lut_4_lut (.I0(n8_adj_4717), .I1(n48649), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29627));
    defparam i15551_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1602 (.I0(n22902), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [5]), .O(n48118));
    defparam i1_2_lut_4_lut_adj_1602.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut_adj_1603 (.I0(\FRAME_MATCHER.state [3]), .I1(n11_adj_4702), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n48641));   // verilog/coms.v(113[11:16])
    defparam i1_2_lut_3_lut_adj_1603.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_345_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4717));   // verilog/coms.v(155[7:23])
    defparam equal_345_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_336_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4734));   // verilog/coms.v(155[7:23])
    defparam equal_336_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 n56626_bdd_4_lut (.I0(n56626), .I1(n56473), .I2(n7_adj_4838), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n56626_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1604 (.I0(n27153), .I1(n105), .I2(n21), 
            .I3(n41963), .O(n4599));   // verilog/coms.v(213[5:16])
    defparam i1_3_lut_4_lut_adj_1604.LUT_INIT = 16'hbbb0;
    SB_LUT4 i1_2_lut_4_lut_adj_1605 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[1] [3]), .I3(n48919), .O(n49201));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_4_lut_adj_1605.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1606 (.I0(n27153), .I1(n105), .I2(n35749), 
            .I3(tx_transmit_N_3748), .O(n4_adj_4626));   // verilog/coms.v(213[5:16])
    defparam i1_3_lut_4_lut_adj_1606.LUT_INIT = 16'h4440;
    SB_LUT4 i1_2_lut_4_lut_adj_1607 (.I0(n22902), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [6]), .O(n48120));
    defparam i1_2_lut_4_lut_adj_1607.LUT_INIT = 16'hf800;
    SB_LUT4 i39809_3_lut_4_lut (.I0(n27153), .I1(n105), .I2(n63_adj_6), 
            .I3(n35749), .O(n28649));   // verilog/coms.v(213[5:16])
    defparam i39809_3_lut_4_lut.LUT_INIT = 16'h0f4f;
    SB_LUT4 i15536_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48649), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n29612));
    defparam i15536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1608 (.I0(n22902), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [7]), .O(n48122));
    defparam i1_2_lut_4_lut_adj_1608.LUT_INIT = 16'hf800;
    SB_LUT4 i15537_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48649), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n29613));
    defparam i15537_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1609 (.I0(n22902), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [8]), .O(n48124));
    defparam i1_2_lut_4_lut_adj_1609.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_4_lut_adj_1610 (.I0(\data_in_frame[11] [3]), .I1(n7_adj_4678), 
            .I2(n48922), .I3(\data_in_frame[9] [1]), .O(n49192));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_4_lut_adj_1610.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1611 (.I0(n22902), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [9]), .O(n48126));
    defparam i1_2_lut_4_lut_adj_1611.LUT_INIT = 16'hf800;
    SB_LUT4 i15538_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48649), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n29614));
    defparam i15538_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15539_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48649), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n29615));
    defparam i15539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1612 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [10]), .O(n48128));
    defparam i1_2_lut_4_lut_adj_1612.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_4_lut_adj_1613 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [11]), .O(n48130));
    defparam i1_2_lut_4_lut_adj_1613.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_adj_1614 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_1079), 
            .I2(GND_net), .I3(GND_net), .O(n48899));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1614.LUT_INIT = 16'h6666;
    SB_LUT4 i15540_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48649), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n29616));
    defparam i15540_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1615 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [3]), 
            .I2(n48704), .I3(n6_adj_4829), .O(Kp_23__N_1079));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1615.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1616 (.I0(\FRAME_MATCHER.state [2]), .I1(n48641), 
            .I2(GND_net), .I3(GND_net), .O(n57));
    defparam i1_2_lut_adj_1616.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1617 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_1079), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[2] [1]), .O(n23));
    defparam i6_4_lut_adj_1617.LUT_INIT = 16'h2184;
    SB_LUT4 i9_3_lut (.I0(n24561), .I1(\data_in_frame[1] [3]), .I2(\data_in_frame[1] [2]), 
            .I3(GND_net), .O(n26_adj_4845));
    defparam i9_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i15541_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48649), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n29617));
    defparam i15541_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1618 (.I0(n23), .I1(n27556), .I2(\data_in_frame[0] [6]), 
            .I3(n48722), .O(n29));
    defparam i12_4_lut_adj_1618.LUT_INIT = 16'h2002;
    SB_LUT4 i5_4_lut_adj_1619 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n48758), .I3(n48899), .O(n22_adj_4846));
    defparam i5_4_lut_adj_1619.LUT_INIT = 16'h1248;
    SB_LUT4 i1_2_lut_4_lut_adj_1620 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [12]), .O(n48132));
    defparam i1_2_lut_4_lut_adj_1620.LUT_INIT = 16'hf800;
    SB_LUT4 i15_4_lut_adj_1621 (.I0(n29), .I1(n6_adj_4671), .I2(n26_adj_4845), 
            .I3(n28051), .O(n32));
    defparam i15_4_lut_adj_1621.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_4_lut_adj_1622 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [13]), .O(n48134));
    defparam i1_2_lut_4_lut_adj_1622.LUT_INIT = 16'hf800;
    SB_LUT4 i15542_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48649), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n29618));
    defparam i15542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1623 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(n28047), .I3(\data_in_frame[1] [5]), .O(n27_adj_4847));
    defparam i10_4_lut_adj_1623.LUT_INIT = 16'h0800;
    SB_LUT4 i16_4_lut_adj_1624 (.I0(n27_adj_4847), .I1(n32), .I2(n52716), 
            .I3(n22_adj_4846), .O(\FRAME_MATCHER.state_31__N_2943 [3]));
    defparam i16_4_lut_adj_1624.LUT_INIT = 16'h0800;
    SB_LUT4 i15543_3_lut_4_lut (.I0(n8_adj_4734), .I1(n48649), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n29619));
    defparam i15543_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1625 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [17]), .O(n48158));
    defparam i1_2_lut_4_lut_adj_1625.LUT_INIT = 16'hf800;
    SB_LUT4 i2_4_lut_adj_1626 (.I0(\FRAME_MATCHER.state_31__N_2943 [3]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n57), .I3(n28717), .O(n24373));
    defparam i2_4_lut_adj_1626.LUT_INIT = 16'h8808;
    SB_LUT4 i21628_3_lut (.I0(\data_in[3]_c [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n35689));   // verilog/coms.v(91[7:20])
    defparam i21628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1627 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [18]), .O(n48160));
    defparam i1_2_lut_4_lut_adj_1627.LUT_INIT = 16'hf800;
    SB_LUT4 i21625_3_lut (.I0(\data_in[3][5] ), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n35686));   // verilog/coms.v(91[7:20])
    defparam i21625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1628 (.I0(n165), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state [1]), 
            .O(\FRAME_MATCHER.i_31__N_2843 ));
    defparam i2_3_lut_4_lut_adj_1628.LUT_INIT = 16'h0040;
    SB_LUT4 i21626_3_lut (.I0(\data_in[3]_c [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29348));   // verilog/coms.v(91[7:20])
    defparam i21626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1629 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [19]), .O(n48162));
    defparam i1_2_lut_4_lut_adj_1629.LUT_INIT = 16'hf800;
    SB_LUT4 i21631_3_lut (.I0(\data_in[2]_c [7]), .I1(\data_in[3]_c [7]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n35692));   // verilog/coms.v(91[7:20])
    defparam i21631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1630 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [20]), .O(n48164));
    defparam i1_2_lut_4_lut_adj_1630.LUT_INIT = 16'hf800;
    SB_LUT4 equal_330_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4710));   // verilog/coms.v(155[7:23])
    defparam equal_330_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_4_lut_adj_1631 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [21]), .O(n48166));
    defparam i1_2_lut_4_lut_adj_1631.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_4_lut_adj_1632 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [22]), .O(n48168));
    defparam i1_2_lut_4_lut_adj_1632.LUT_INIT = 16'hf800;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_40720 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n56296));
    defparam byte_transmit_counter_0__bdd_4_lut_40720.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1633 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[5] [0]), .I3(GND_net), .O(n49069));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1633.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1634 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n28047));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1634.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1635 (.I0(n4_adj_4735), .I1(n48925), .I2(\data_in_frame[9] [5]), 
            .I3(\data_in_frame[11] [6]), .O(n49170));
    defparam i1_2_lut_4_lut_adj_1635.LUT_INIT = 16'h6996;
    SB_LUT4 equal_331_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4625));   // verilog/coms.v(155[7:23])
    defparam equal_331_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15784_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48665), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n29860));
    defparam i15784_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15785_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48665), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n29861));
    defparam i15785_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1636 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[11] [7]), 
            .I2(n45470), .I3(GND_net), .O(n49260));
    defparam i1_2_lut_3_lut_adj_1636.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1637 (.I0(\data_in_frame[12] [4]), .I1(n27669), 
            .I2(n45522), .I3(GND_net), .O(n49004));
    defparam i1_2_lut_3_lut_adj_1637.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1638 (.I0(n48781), .I1(n49266), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4848));
    defparam i1_2_lut_adj_1638.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1639 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[20] [7]), 
            .I2(n49165), .I3(n6_adj_4848), .O(n46365));
    defparam i4_4_lut_adj_1639.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1640 (.I0(n46365), .I1(n46363), .I2(GND_net), 
            .I3(GND_net), .O(n45486));
    defparam i1_2_lut_adj_1640.LUT_INIT = 16'h6666;
    SB_LUT4 i15786_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48665), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n29862));
    defparam i15786_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1641 (.I0(\FRAME_MATCHER.state [5]), .I1(\FRAME_MATCHER.state [12]), 
            .I2(\FRAME_MATCHER.state [10]), .I3(\FRAME_MATCHER.state [7]), 
            .O(n16_adj_4849));   // verilog/coms.v(128[12] 303[6])
    defparam i6_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 i15787_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48665), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n29863));
    defparam i15787_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n56296_bdd_4_lut (.I0(n56296), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n56299));
    defparam n56296_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_40505 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n56290));
    defparam byte_transmit_counter_0__bdd_4_lut_40505.LUT_INIT = 16'he4aa;
    SB_LUT4 i7_4_lut_adj_1642 (.I0(\FRAME_MATCHER.state [11]), .I1(\FRAME_MATCHER.state [15]), 
            .I2(\FRAME_MATCHER.state [8]), .I3(\FRAME_MATCHER.state [14]), 
            .O(n17_adj_4850));   // verilog/coms.v(128[12] 303[6])
    defparam i7_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1643 (.I0(n17_adj_4850), .I1(\FRAME_MATCHER.state [9]), 
            .I2(n16_adj_4849), .I3(\FRAME_MATCHER.state [13]), .O(n48560));   // verilog/coms.v(128[12] 303[6])
    defparam i9_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 n56290_bdd_4_lut (.I0(n56290), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n56293));
    defparam n56290_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15788_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48665), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n29864));
    defparam i15788_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n56596_bdd_4_lut (.I0(n56596), .I1(n56485), .I2(n7_adj_4837), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n56596_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1644 (.I0(\FRAME_MATCHER.state [30]), .I1(\FRAME_MATCHER.state [29]), 
            .I2(\FRAME_MATCHER.state [23]), .I3(\FRAME_MATCHER.state [27]), 
            .O(n50821));   // verilog/coms.v(128[12] 303[6])
    defparam i3_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 i15789_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48665), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n29865));
    defparam i15789_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21627_3_lut (.I0(\data_in[2][1] ), .I1(\data_in[3]_c [1]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n29356));   // verilog/coms.v(91[7:20])
    defparam i21627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_40749 (.I0(byte_transmit_counter[3]), 
            .I1(n56425), .I2(n54302), .I3(byte_transmit_counter[4]), .O(n56590));
    defparam byte_transmit_counter_3__bdd_4_lut_40749.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_4_lut_adj_1645 (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [18]), 
            .I2(\FRAME_MATCHER.state [17]), .I3(\FRAME_MATCHER.state [24]), 
            .O(n12_adj_4851));   // verilog/coms.v(128[12] 303[6])
    defparam i5_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1646 (.I0(\FRAME_MATCHER.state [19]), .I1(n12_adj_4851), 
            .I2(n50821), .I3(\FRAME_MATCHER.state [20]), .O(n46240));   // verilog/coms.v(128[12] 303[6])
    defparam i6_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1647 (.I0(\FRAME_MATCHER.state [26]), .I1(\FRAME_MATCHER.state [22]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4852));
    defparam i2_2_lut_adj_1647.LUT_INIT = 16'heeee;
    SB_LUT4 i15790_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48665), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n29866));
    defparam i15790_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1648 (.I0(\FRAME_MATCHER.state [16]), .I1(\FRAME_MATCHER.state [6]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [28]), 
            .O(n14_adj_4853));
    defparam i6_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i15338_3_lut_4_lut (.I0(n8_adj_4631), .I1(n48665), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n29414));
    defparam i15338_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1649 (.I0(\FRAME_MATCHER.state [25]), .I1(n14_adj_4853), 
            .I2(n10_adj_4852), .I3(\FRAME_MATCHER.state [4]), .O(n48679));
    defparam i7_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i15528_3_lut_4_lut (.I0(n10_adj_4630), .I1(n48645), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n29604));
    defparam i15528_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21629_3_lut (.I0(\data_in[1]_c [7]), .I1(\data_in[2]_c [7]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n29359));   // verilog/coms.v(91[7:20])
    defparam i21629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1650 (.I0(n48679), .I1(n46240), .I2(n48560), 
            .I3(GND_net), .O(n41963));   // verilog/coms.v(128[12] 303[6])
    defparam i2_3_lut_adj_1650.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1651 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n41963), .I3(GND_net), .O(n27119));   // verilog/coms.v(128[12] 303[6])
    defparam i1_2_lut_3_lut_adj_1651.LUT_INIT = 16'hfefe;
    SB_LUT4 i15529_3_lut_4_lut (.I0(n10_adj_4630), .I1(n48645), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n29605));
    defparam i15529_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1652 (.I0(n28075), .I1(n48916), .I2(\data_in_frame[12] [5]), 
            .I3(n27669), .O(n27661));
    defparam i1_2_lut_4_lut_adj_1652.LUT_INIT = 16'h6996;
    SB_LUT4 i15530_3_lut_4_lut (.I0(n10_adj_4630), .I1(n48645), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n29606));
    defparam i15530_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15531_3_lut_4_lut (.I0(n10_adj_4630), .I1(n48645), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n29607));
    defparam i15531_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15532_3_lut_4_lut (.I0(n10_adj_4630), .I1(n48645), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n29608));
    defparam i15532_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15533_3_lut_4_lut (.I0(n10_adj_4630), .I1(n48645), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n29609));
    defparam i15533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1653 (.I0(n27556), .I1(n28047), .I2(n49149), 
            .I3(GND_net), .O(n49198));   // verilog/coms.v(79[16:27])
    defparam i1_2_lut_3_lut_adj_1653.LUT_INIT = 16'h6969;
    SB_LUT4 i21630_3_lut (.I0(\data_in[0]_c [7]), .I1(\data_in[1]_c [7]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n29367));   // verilog/coms.v(91[7:20])
    defparam i21630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1654 (.I0(\FRAME_MATCHER.state [3]), .I1(n41963), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/coms.v(128[12] 303[6])
    defparam i1_2_lut_adj_1654.LUT_INIT = 16'heeee;
    SB_LUT4 i15534_3_lut_4_lut (.I0(n10_adj_4630), .I1(n48645), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n29610));
    defparam i15534_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15535_3_lut_4_lut (.I0(n10_adj_4630), .I1(n48645), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n29611));
    defparam i15535_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1655 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n35747), .O(n49999));
    defparam i2_3_lut_4_lut_adj_1655.LUT_INIT = 16'h8000;
    SB_LUT4 equal_333_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4631));
    defparam equal_333_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1656 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n35747), .O(n48665));   // verilog/coms.v(155[7:23])
    defparam i1_2_lut_4_lut_adj_1656.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_1657 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n48645), .O(n48646));   // verilog/coms.v(155[7:23])
    defparam i1_2_lut_4_lut_adj_1657.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1658 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(n48796), .I3(GND_net), .O(Kp_23__N_1098));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_3_lut_adj_1658.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1659 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n49999), .O(n48638));   // verilog/coms.v(155[7:23])
    defparam i1_2_lut_4_lut_adj_1659.LUT_INIT = 16'hfbff;
    SB_LUT4 i15393_3_lut_4_lut (.I0(n8), .I1(n48665), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n29469));
    defparam i15393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1660 (.I0(\data_in_frame[0] [5]), .I1(n27549), 
            .I2(n48796), .I3(\data_in_frame[1] [0]), .O(n26308));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_4_lut_adj_1660.LUT_INIT = 16'h6996;
    SB_LUT4 i15394_3_lut_4_lut (.I0(n8), .I1(n48665), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n29470));
    defparam i15394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15395_3_lut_4_lut (.I0(n8), .I1(n48665), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n29471));
    defparam i15395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1661 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [23]), .O(n48170));
    defparam i1_2_lut_4_lut_adj_1661.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_4_lut_adj_1662 (.I0(\data_in_frame[13] [2]), .I1(n50394), 
            .I2(\data_in_frame[13] [3]), .I3(\data_in_frame[15] [4]), .O(n49010));
    defparam i1_2_lut_4_lut_adj_1662.LUT_INIT = 16'h9669;
    SB_LUT4 i15440_3_lut_4_lut (.I0(n10), .I1(n49999), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n29516));
    defparam i15440_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15441_3_lut_4_lut (.I0(n10), .I1(n49999), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n29517));
    defparam i15441_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15442_3_lut_4_lut (.I0(n10), .I1(n49999), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n29518));
    defparam i15442_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15396_3_lut_4_lut (.I0(n8), .I1(n48665), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n29472));
    defparam i15396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1663 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [24]), .O(n48172));
    defparam i1_2_lut_4_lut_adj_1663.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut_adj_1664 (.I0(n28032), .I1(n27916), .I2(n49157), 
            .I3(GND_net), .O(n48799));   // verilog/coms.v(86[17:63])
    defparam i1_2_lut_3_lut_adj_1664.LUT_INIT = 16'h9696;
    SB_LUT4 i15397_3_lut_4_lut (.I0(n8), .I1(n48665), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n29473));
    defparam i15397_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1665 (.I0(\data_in_frame[10] [7]), .I1(n48731), 
            .I2(n49423), .I3(GND_net), .O(n46429));
    defparam i1_2_lut_3_lut_adj_1665.LUT_INIT = 16'h9696;
    SB_LUT4 i15398_3_lut_4_lut (.I0(n8), .I1(n48665), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n29474));
    defparam i15398_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15399_3_lut_4_lut (.I0(n8), .I1(n48665), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n29475));
    defparam i15399_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15443_3_lut_4_lut (.I0(n10), .I1(n49999), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n29519));
    defparam i15443_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15337_3_lut_4_lut (.I0(n8), .I1(n48665), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n29413));
    defparam i15337_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_40774 (.I0(byte_transmit_counter[3]), 
            .I1(n56329), .I2(n54289), .I3(byte_transmit_counter[4]), .O(n56620));
    defparam byte_transmit_counter_3__bdd_4_lut_40774.LUT_INIT = 16'he4aa;
    SB_LUT4 n56620_bdd_4_lut (.I0(n56620), .I1(n14_adj_4844), .I2(n7_adj_4836), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n56620_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1666 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n35747), .O(n48645));   // verilog/coms.v(155[7:23])
    defparam i2_3_lut_4_lut_adj_1666.LUT_INIT = 16'hfbff;
    SB_LUT4 equal_342_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(155[7:23])
    defparam equal_342_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i39851_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n48641), .I3(GND_net), .O(n124));
    defparam i39851_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i39800_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n29040));
    defparam i39800_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i15444_3_lut_4_lut (.I0(n10), .I1(n49999), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n29520));
    defparam i15444_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15520_3_lut_4_lut (.I0(n8), .I1(n48649), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n29596));
    defparam i15520_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1667 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[15] [7]), 
            .I2(n10_adj_4731), .I3(n27661), .O(n6_adj_4709));
    defparam i1_2_lut_4_lut_adj_1667.LUT_INIT = 16'h6996;
    SB_LUT4 i22391_2_lut_4_lut (.I0(n24561), .I1(n31_adj_4679), .I2(n31), 
            .I3(\FRAME_MATCHER.state [1]), .O(n1));
    defparam i22391_2_lut_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_2_lut_3_lut_adj_1668 (.I0(\data_in_frame[20] [0]), .I1(\data_in_frame[15] [5]), 
            .I2(n45384), .I3(GND_net), .O(n46393));
    defparam i1_2_lut_3_lut_adj_1668.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1669 (.I0(n45137), .I1(n45514), .I2(\data_in_frame[20] [1]), 
            .I3(n52240), .O(n52244));
    defparam i1_3_lut_4_lut_adj_1669.LUT_INIT = 16'h6996;
    SB_LUT4 i15521_3_lut_4_lut (.I0(n8), .I1(n48649), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n29597));
    defparam i15521_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1670 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n7936));
    defparam i1_2_lut_3_lut_adj_1670.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_4_lut_adj_1671 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [25]), .O(n48174));
    defparam i1_2_lut_4_lut_adj_1671.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_4_lut_adj_1672 (.I0(\data_in_frame[18] [5]), .I1(n49029), 
            .I2(\data_in_frame[16] [5]), .I3(n28010), .O(n48781));
    defparam i1_2_lut_4_lut_adj_1672.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1673 (.I0(\data_in_frame[17] [3]), .I1(n46462), 
            .I2(n51116), .I3(GND_net), .O(n46481));
    defparam i1_2_lut_3_lut_adj_1673.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1674 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [1]), 
            .I2(n48736), .I3(\data_in_frame[15] [3]), .O(n52522));   // verilog/coms.v(72[16:27])
    defparam i1_3_lut_4_lut_adj_1674.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1675 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n144));
    defparam i1_2_lut_3_lut_adj_1675.LUT_INIT = 16'hfefe;
    SB_LUT4 i15522_3_lut_4_lut (.I0(n8), .I1(n48649), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n29598));
    defparam i15522_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1676 (.I0(n46240), .I1(n48679), .I2(n48560), 
            .I3(GND_net), .O(n11_adj_4702));
    defparam i1_2_lut_3_lut_adj_1676.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1677 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n46409), .I3(GND_net), .O(n49084));
    defparam i1_2_lut_3_lut_adj_1677.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1678 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [26]), .O(n48176));
    defparam i1_2_lut_4_lut_adj_1678.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_4_lut_adj_1679 (.I0(\data_in_frame[16] [5]), .I1(n28010), 
            .I2(\data_in_frame[16] [4]), .I3(n46475), .O(n45137));
    defparam i1_2_lut_4_lut_adj_1679.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1680 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[4] [0]), .I3(n27515), .O(n52116));
    defparam i1_2_lut_4_lut_adj_1680.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1681 (.I0(\data_in_frame[17] [3]), .I1(n46462), 
            .I2(n46367), .I3(\data_in_frame[19] [4]), .O(n46389));
    defparam i1_3_lut_4_lut_adj_1681.LUT_INIT = 16'h9669;
    SB_LUT4 i15523_3_lut_4_lut (.I0(n8), .I1(n48649), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n29599));
    defparam i15523_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15445_3_lut_4_lut (.I0(n10), .I1(n49999), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n29521));
    defparam i15445_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_3_lut_4_lut_adj_1682 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[2] [3]), 
            .I2(n48704), .I3(\data_in_frame[4] [4]), .O(n49087));   // verilog/coms.v(75[16:43])
    defparam i1_3_lut_4_lut_adj_1682.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1683 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [27]), .O(n48178));
    defparam i1_2_lut_4_lut_adj_1683.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_4_lut_adj_1684 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[9] [4]), .I3(n49260), .O(n6_adj_4670));
    defparam i1_2_lut_4_lut_adj_1684.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1685 (.I0(n48983), .I1(n46475), .I2(\data_in_frame[16] [3]), 
            .I3(n25573), .O(n46407));
    defparam i1_2_lut_4_lut_adj_1685.LUT_INIT = 16'h9669;
    SB_LUT4 i29_3_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n11));
    defparam i29_3_lut_3_lut.LUT_INIT = 16'h8181;
    SB_LUT4 select_713_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4715));
    defparam select_713_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_713_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n4623), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4713));
    defparam select_713_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1686 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n27325), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_4654));
    defparam i1_3_lut_4_lut_adj_1686.LUT_INIT = 16'hfefc;
    SB_LUT4 i2_2_lut_3_lut_adj_1687 (.I0(\data_in_frame[20] [7]), .I1(\data_in_frame[20] [6]), 
            .I2(n49336), .I3(GND_net), .O(n7_adj_4629));
    defparam i2_2_lut_3_lut_adj_1687.LUT_INIT = 16'h9696;
    SB_LUT4 i15524_3_lut_4_lut (.I0(n8), .I1(n48649), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n29600));
    defparam i15524_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15525_3_lut_4_lut (.I0(n8), .I1(n48649), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n29601));
    defparam i15525_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_40784 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n56614));
    defparam byte_transmit_counter_0__bdd_4_lut_40784.LUT_INIT = 16'he4aa;
    SB_LUT4 i15526_3_lut_4_lut (.I0(n8), .I1(n48649), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n29602));
    defparam i15526_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1688 (.I0(n49029), .I1(\data_in_frame[16] [5]), 
            .I2(n28010), .I3(GND_net), .O(n50318));
    defparam i2_2_lut_3_lut_adj_1688.LUT_INIT = 16'h9696;
    SB_LUT4 i37054_3_lut_4_lut (.I0(n22902), .I1(\FRAME_MATCHER.i_31__N_2843 ), 
            .I2(n3303), .I3(n4599), .O(n48674));
    defparam i37054_3_lut_4_lut.LUT_INIT = 16'haa08;
    SB_LUT4 i1_2_lut_3_lut_adj_1689 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [5]), 
            .I2(\data_in_frame[16] [7]), .I3(GND_net), .O(n49397));
    defparam i1_2_lut_3_lut_adj_1689.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1690 (.I0(n41963), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n27278), .I3(\FRAME_MATCHER.state [3]), .O(n63_adj_6));   // verilog/coms.v(128[12] 303[6])
    defparam i2_3_lut_4_lut_adj_1690.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_4_lut_adj_1691 (.I0(n27208), .I1(n4_adj_4626), .I2(n2_adj_4627), 
            .I3(\FRAME_MATCHER.state [28]), .O(n48180));
    defparam i1_2_lut_4_lut_adj_1691.LUT_INIT = 16'hf800;
    SB_LUT4 i15446_3_lut_4_lut (.I0(n10), .I1(n49999), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n29522));
    defparam i15446_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_2_lut_3_lut_adj_1692 (.I0(\data_in_frame[12] [1]), .I1(n45569), 
            .I2(n46531), .I3(GND_net), .O(n6));
    defparam i2_2_lut_3_lut_adj_1692.LUT_INIT = 16'h9696;
    uart_tx tx (.GND_net(GND_net), .n28758(n28758), .clk16MHz(clk16MHz), 
            .n29184(n29184), .\r_Bit_Index[0] (\r_Bit_Index[0] ), .\r_SM_Main_2__N_3851[0] (r_SM_Main_2__N_3851[0]), 
            .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3848[1] (\r_SM_Main_2__N_3848[1] ), 
            .VCC_net(VCC_net), .tx_o(tx_o), .tx_data({tx_data}), .n29324(n29324), 
            .tx_active(tx_active), .n29732(n29732), .n56700(n56700), .n4(n4_adj_8), 
            .tx_enable(tx_enable), .n19731(n19731)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(108[10:70])
    uart_rx rx (.n28762(n28762), .clk16MHz(clk16MHz), .n29186(n29186), 
            .n29420(n29420), .rx_data({rx_data}), .r_SM_Main({r_SM_Main_adj_16}), 
            .r_Rx_Data(r_Rx_Data), .GND_net(GND_net), .\r_SM_Main_2__N_3777[2] (\r_SM_Main_2__N_3777[2] ), 
            .n35837(n35837), .VCC_net(VCC_net), .RX_N_10(RX_N_10), .n4(n4_adj_12), 
            .n4_adj_4(n4_adj_13), .n29735(n29735), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_14 ), 
            .n48270(n48270), .rx_data_ready(rx_data_ready), .n29261(n29261), 
            .n4_adj_5(n4_adj_15), .n29769(n29769), .n29767(n29767), .n29766(n29766), 
            .n48565(n48565), .n29749(n29749), .n29748(n29748), .n29740(n29740), 
            .n27227(n27227), .n27232(n27232)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(94[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (GND_net, n28758, clk16MHz, n29184, \r_Bit_Index[0] , 
            \r_SM_Main_2__N_3851[0] , r_SM_Main, \r_SM_Main_2__N_3848[1] , 
            VCC_net, tx_o, tx_data, n29324, tx_active, n29732, n56700, 
            n4, tx_enable, n19731) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n28758;
    input clk16MHz;
    output n29184;
    output \r_Bit_Index[0] ;
    input \r_SM_Main_2__N_3851[0] ;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3848[1] ;
    input VCC_net;
    output tx_o;
    input [7:0]tx_data;
    input n29324;
    output tx_active;
    input n29732;
    input n56700;
    output n4;
    output tx_enable;
    output n19731;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [8:0]n41;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n44172, n44171;
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n1, n29083, n44170, n44169;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n52967, n52968, n52971, n52970, n44168, n36449, n21947, 
        n21948, o_Tx_Serial_N_3879, n3, n44167, n44166, n44165, 
        n26737, n3_adj_4623, n56380, n50757, n10;
    
    SB_LUT4 r_Clock_Count_2292_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n44172), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2292_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n44171), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_9 (.CI(n44171), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n44172));
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n28758), 
            .D(n307[1]), .R(n29184));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n28758), 
            .D(n307[2]), .R(n29184));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_2292__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n29083));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 r_Clock_Count_2292_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n44170), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_8 (.CI(n44170), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n44171));
    SB_LUT4 r_Clock_Count_2292_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n44169), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_7 (.CI(n44169), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n44170));
    SB_LUT4 i37175_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n52967));
    defparam i37175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37176_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n52968));
    defparam i37176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37179_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n52971));
    defparam i37179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37178_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n52970));
    defparam i37178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_2292_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n44168), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7988_4_lut (.I0(\r_SM_Main_2__N_3851[0] ), .I1(n36449), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3848[1] ), .O(n21947));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7988_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7989_3_lut (.I0(n21947), .I1(\r_SM_Main_2__N_3848[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n21948));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7989_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3879), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_CARRY r_Clock_Count_2292_add_4_6 (.CI(n44168), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n44169));
    SB_LUT4 r_Clock_Count_2292_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n44167), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_5 (.CI(n44167), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n44168));
    SB_LUT4 r_Clock_Count_2292_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n44166), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_4 (.CI(n44166), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n44167));
    SB_LUT4 r_Clock_Count_2292_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n44165), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_3 (.CI(n44165), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n44166));
    SB_LUT4 r_Clock_Count_2292_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2292_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2292_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n44165));
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n26737), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n21948), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_2292__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n29083));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n29083));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n29083));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n29083));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n29083));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n29083));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n29083));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2292__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n29083));   // verilog/uart_tx.v(118[34:51])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk16MHz), .D(n29324));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29732));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n56700));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_4623), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n26737), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n26737), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n26737), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n26737), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n26737), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n26737), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n26737), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n52970), 
            .I2(n52971), .I3(r_Bit_Index[2]), .O(n56380));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n56380_bdd_4_lut (.I0(n56380), .I1(n52968), .I2(n52967), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3879));
    defparam n56380_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i39845_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3848[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n29083));
    defparam i39845_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2474_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i2474_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[2]), .O(n50757));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), .I2(n50757), 
            .I3(r_Clock_Count[8]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3848[1] ));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n36449));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i15108_3_lut (.I0(n28758), .I1(n36449), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n29184));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15108_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i10001_2_lut_3_lut (.I0(\r_SM_Main_2__N_3848[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4623));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i10001_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2467_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i2467_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3851[0] ), 
            .I3(r_SM_Main[1]), .O(n26737));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3848[1] ), .O(n28758));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3848[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5781_2_lut (.I0(\r_SM_Main_2__N_3851[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n19731));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5781_2_lut.LUT_INIT = 16'h2222;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n28762, clk16MHz, n29186, n29420, rx_data, r_SM_Main, 
            r_Rx_Data, GND_net, \r_SM_Main_2__N_3777[2] , n35837, VCC_net, 
            RX_N_10, n4, n4_adj_4, n29735, \r_Bit_Index[0] , n48270, 
            rx_data_ready, n29261, n4_adj_5, n29769, n29767, n29766, 
            n48565, n29749, n29748, n29740, n27227, n27232) /* synthesis syn_module_defined=1 */ ;
    output n28762;
    input clk16MHz;
    output n29186;
    input n29420;
    output [7:0]rx_data;
    output [2:0]r_SM_Main;
    output r_Rx_Data;
    input GND_net;
    output \r_SM_Main_2__N_3777[2] ;
    output n35837;
    input VCC_net;
    input RX_N_10;
    output n4;
    output n4_adj_4;
    input n29735;
    output \r_Bit_Index[0] ;
    input n48270;
    output rx_data_ready;
    input n29261;
    output n4_adj_5;
    input n29769;
    input n29767;
    input n29766;
    input n48565;
    input n29749;
    input n29748;
    input n29740;
    output n27227;
    output n27232;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [7:0]n37;
    
    wire n28712;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n29092;
    wire [2:0]r_SM_Main_2__N_3783;
    
    wire n54256, n36620, n36447, n36574, n1, n3, n44164, n44163, 
        n44162, n44161, n44160, n44159, n44158, r_Rx_Data_R, n9, 
        n27112, n54316, n54314, n6, n6_adj_4621, n6_adj_4622;
    
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n28762), 
            .D(n326[1]), .R(n29186));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n28762), 
            .D(n326[2]), .R(n29186));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29420));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_2290__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n28712), .D(n37[0]), .R(n29092));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i38610_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3783[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n54256));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i38610_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n54256), .I1(\r_SM_Main_2__N_3777[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n36620));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_LUT4 i21777_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35837));
    defparam i21777_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n36447), .I1(\r_SM_Main_2__N_3777[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n36574));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3783[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n36574), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_Clock_Count_2290_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n44164), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2290_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n44163), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_8 (.CI(n44163), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n44164));
    SB_LUT4 r_Clock_Count_2290_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n44162), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_7 (.CI(n44162), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n44163));
    SB_LUT4 r_Clock_Count_2290_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n44161), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_6 (.CI(n44161), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n44162));
    SB_LUT4 r_Clock_Count_2290_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n44160), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_5 (.CI(n44160), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n44161));
    SB_DFFESR r_Clock_Count_2290__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n28712), .D(n37[1]), .R(n29092));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_2290_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n44159), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_4 (.CI(n44159), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n44160));
    SB_LUT4 r_Clock_Count_2290_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n44158), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2290_add_4_3 (.CI(n44158), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n44159));
    SB_LUT4 r_Clock_Count_2290_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2290_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_CARRY r_Clock_Count_2290_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n44158));
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_2290__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n28712), .D(n37[2]), .R(n29092));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2290__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n28712), .D(n37[3]), .R(n29092));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2290__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n28712), .D(n37[4]), .R(n29092));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2290__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n28712), .D(n37[5]), .R(n29092));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2290__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n28712), .D(n37[6]), .R(n29092));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2290__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n28712), .D(n37[7]), .R(n29092));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 equal_379_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_379_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_377_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_377_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29735));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk16MHz), .D(n48270));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n29261));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n36620), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i4_4_lut (.I0(n9), .I1(n27112), .I2(r_Clock_Count[3]), .I3(r_Clock_Count[1]), 
            .O(r_SM_Main_2__N_3783[0]));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i3_2_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(GND_net), .O(n9));
    defparam i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38592_4_lut (.I0(r_Rx_Data), .I1(r_Clock_Count[1]), .I2(n27112), 
            .I3(r_Clock_Count[3]), .O(n54316));
    defparam i38592_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i38855_3_lut (.I0(n54316), .I1(r_SM_Main[0]), .I2(n9), .I3(GND_net), 
            .O(n54314));
    defparam i38855_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n54314), .I2(\r_SM_Main_2__N_3777[2] ), 
            .I3(r_SM_Main[1]), .O(n29092));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_2__N_3783[0]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i39798_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_Rx_Data), .O(n28712));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i39798_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 equal_375_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5));   // verilog/uart_rx.v(97[17:39])
    defparam equal_375_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29769));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29767));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29766));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n48565));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n29749));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29748));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n29740));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2452_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i2452_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_3_lut_4_lut (.I0(\r_SM_Main_2__N_3777[2] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n28762));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0203;
    SB_LUT4 i1_2_lut_4_lut (.I0(n6_adj_4621), .I1(\r_SM_Main_2__N_3777[2] ), 
            .I2(r_SM_Main[1]), .I3(\r_Bit_Index[0] ), .O(n27227));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_4_lut_adj_953 (.I0(n6_adj_4621), .I1(\r_SM_Main_2__N_3777[2] ), 
            .I2(r_SM_Main[1]), .I3(\r_Bit_Index[0] ), .O(n27232));
    defparam i1_2_lut_4_lut_adj_953.LUT_INIT = 16'hffbf;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[5]), .O(n27112));   // verilog/uart_rx.v(118[17:47])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_954 (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4621));
    defparam i2_2_lut_adj_954.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_955 (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4622));
    defparam i2_2_lut_adj_955.LUT_INIT = 16'h8888;
    SB_LUT4 i22383_4_lut (.I0(r_Clock_Count[0]), .I1(n27112), .I2(n6_adj_4622), 
            .I3(r_Clock_Count[1]), .O(\r_SM_Main_2__N_3777[2] ));
    defparam i22383_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n36447));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i15110_3_lut (.I0(n28762), .I1(n36447), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n29186));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15110_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2445_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i2445_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (\state[0] , \state[1] , state_7__N_4499, GND_net, \data[12] , 
            clk16MHz, VCC_net, \data[15] , n28640, n35803, n15, 
            n35841, n6, n5, n29966, \data[10] , n5_adj_1, n29965, 
            \data[9] , n29959, \data[8] , n29958, \data[7] , n29320, 
            n29317, \data[11] , n9, clk_out, n29308, CS_c, n29301, 
            \current[0] , n6_adj_2, n5_adj_3, n7, \current[15] , CS_CLK_c, 
            n29805, \data[6] , n29781, \data[5] , n29780, \current[1] , 
            n29779, \current[2] , n29778, \current[3] , n29777, \current[4] , 
            n29776, \current[5] , n29775, \current[6] , n29774, \current[7] , 
            n29773, \current[8] , n29772, \current[9] , n29771, \current[10] , 
            n29770, \current[11] , n29768, \data[4] , n29763, \data[3] , 
            n29750, \data[2] , n29741, \data[0] , n29736, \data[1] , 
            n29647, n27222, n27287, n27281, n27294, n27256) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[0] ;
    output \state[1] ;
    output state_7__N_4499;
    input GND_net;
    output \data[12] ;
    input clk16MHz;
    input VCC_net;
    output \data[15] ;
    output n28640;
    output n35803;
    output n15;
    output n35841;
    output n6;
    output n5;
    input n29966;
    output \data[10] ;
    output n5_adj_1;
    input n29965;
    output \data[9] ;
    input n29959;
    output \data[8] ;
    input n29958;
    output \data[7] ;
    input n29320;
    input n29317;
    output \data[11] ;
    input n9;
    output clk_out;
    input n29308;
    output CS_c;
    input n29301;
    output \current[0] ;
    output n6_adj_2;
    output n5_adj_3;
    output n7;
    output \current[15] ;
    output CS_CLK_c;
    input n29805;
    output \data[6] ;
    input n29781;
    output \data[5] ;
    input n29780;
    output \current[1] ;
    input n29779;
    output \current[2] ;
    input n29778;
    output \current[3] ;
    input n29777;
    output \current[4] ;
    input n29776;
    output \current[5] ;
    input n29775;
    output \current[6] ;
    input n29774;
    output \current[7] ;
    input n29773;
    output \current[8] ;
    input n29772;
    output \current[9] ;
    input n29771;
    output \current[10] ;
    input n29770;
    output \current[11] ;
    input n29768;
    output \data[4] ;
    input n29763;
    output \data[3] ;
    input n29750;
    output \data[2] ;
    input n29741;
    output \data[0] ;
    input n29736;
    output \data[1] ;
    input n29647;
    output n27222;
    output n27287;
    output n27281;
    output n27294;
    output n27256;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n28709;
    wire [13:0]n241;
    
    wire n7796;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n6_c, clk_slow_N_4413, clk_slow_N_4412, n54291, n24139;
    wire [4:0]n25;
    
    wire n44157, n44156, n44155, n44154;
    wire [13:0]n61;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n44153, n44152, n44151, n44150, n44149, n44148, n44147, 
        n44146, n44145, n44144, n44143, n44142, n44141;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    wire [7:0]n37;
    
    wire n29079, n36267, n24108, n24110, n24112, delay_counter_15__N_4494, 
        n10898, n28785, n29060, n6_adj_4617, n44215, n44214, n44213, 
        n44212, n54245, n44211, n54244, n44210, n54243, n44209, 
        n6_adj_4618, n51100, n49889, n49957;
    
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4499));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14888_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28709));
    defparam i14888_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2419_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2151_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n7796));   // verilog/tli4970.v(35[10] 68[6])
    defparam i2151_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6_c));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2392_4_lut (.I0(counter[0]), .I1(counter[4]), .I2(n6_c), 
            .I3(counter[3]), .O(clk_slow_N_4413));
    defparam i2392_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4413), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4412));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10089_3_lut (.I0(\state[0] ), .I1(n54291), .I2(\state[1] ), 
            .I3(GND_net), .O(n24139));   // verilog/tli4970.v(55[24:39])
    defparam i10089_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4412));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 counter_2287_2288_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n44157), .O(n25[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2287_2288_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2287_2288_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n44156), .O(n25[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2287_2288_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2287_2288_add_4_5 (.CI(n44156), .I0(GND_net), .I1(counter[3]), 
            .CO(n44157));
    SB_LUT4 counter_2287_2288_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n44155), .O(n25[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2287_2288_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2287_2288_add_4_4 (.CI(n44155), .I0(GND_net), .I1(counter[2]), 
            .CO(n44156));
    SB_LUT4 counter_2287_2288_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n44154), .O(n25[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2287_2288_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2287_2288_add_4_3 (.CI(n44154), .I0(GND_net), .I1(counter[1]), 
            .CO(n44155));
    SB_LUT4 counter_2287_2288_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n25[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2287_2288_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2287_2288_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n44154));
    SB_LUT4 delay_counter_2285_2286_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[13]), .I3(n44153), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2285_2286_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[12]), .I3(n44152), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_14 (.CI(n44152), .I0(GND_net), 
            .I1(delay_counter[12]), .CO(n44153));
    SB_LUT4 delay_counter_2285_2286_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n44151), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_13 (.CI(n44151), .I0(GND_net), 
            .I1(delay_counter[11]), .CO(n44152));
    SB_LUT4 delay_counter_2285_2286_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n44150), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_12 (.CI(n44150), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n44151));
    SB_LUT4 delay_counter_2285_2286_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n44149), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_11 (.CI(n44149), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n44150));
    SB_LUT4 delay_counter_2285_2286_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n44148), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_10 (.CI(n44148), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n44149));
    SB_LUT4 delay_counter_2285_2286_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n44147), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_9 (.CI(n44147), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n44148));
    SB_LUT4 delay_counter_2285_2286_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n44146), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_8 (.CI(n44146), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n44147));
    SB_LUT4 delay_counter_2285_2286_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n44145), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_7 (.CI(n44145), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n44146));
    SB_LUT4 delay_counter_2285_2286_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n44144), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_6 (.CI(n44144), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n44145));
    SB_LUT4 delay_counter_2285_2286_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n44143), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_5 (.CI(n44143), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n44144));
    SB_LUT4 delay_counter_2285_2286_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n44142), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_4 (.CI(n44142), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n44143));
    SB_LUT4 delay_counter_2285_2286_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n44141), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_3 (.CI(n44141), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n44142));
    SB_LUT4 delay_counter_2285_2286_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2285_2286_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2285_2286_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n44141));
    SB_LUT4 i39811_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n28640));
    defparam i39811_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i21743_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n35803));
    defparam i21743_2_lut.LUT_INIT = 16'h8888;
    SB_DFFNESR bit_counter_2296__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n28709), 
            .D(n37[4]), .R(n29079));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2296__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n28709), 
            .D(n37[5]), .R(n29079));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2296__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n28709), 
            .D(n37[6]), .R(n29079));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2296__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n28709), 
            .D(n37[7]), .R(n29079));   // verilog/tli4970.v(55[24:39])
    SB_LUT4 i40443_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n36267));
    defparam i40443_2_lut.LUT_INIT = 16'h1111;
    SB_DFFNE bit_counter_2296__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n28709), 
            .D(n24108));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2296__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n28709), 
            .D(n24110));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2296__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n28709), 
            .D(n24112));   // verilog/tli4970.v(55[24:39])
    SB_DFFSR counter_2287_2288__i5 (.Q(counter[4]), .C(clk16MHz), .D(n25[4]), 
            .R(clk_slow_N_4413));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2287_2288__i4 (.Q(counter[3]), .C(clk16MHz), .D(n25[3]), 
            .R(clk_slow_N_4413));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2287_2288__i3 (.Q(counter[2]), .C(clk16MHz), .D(n25[2]), 
            .R(clk_slow_N_4413));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2287_2288__i2 (.Q(counter[1]), .C(clk16MHz), .D(n25[1]), 
            .R(clk_slow_N_4413));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_2285_2286__i14 (.Q(delay_counter[13]), .C(clk_slow), 
            .D(n61[13]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i13 (.Q(delay_counter[12]), .C(clk_slow), 
            .D(n61[12]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n61[11]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n61[10]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n61[9]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n61[8]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n61[7]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n61[6]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n61[5]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n61[4]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n61[3]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n61[2]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2285_2286__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n61[1]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_LUT4 i21781_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n35841));
    defparam i21781_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_364_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_364_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n28785), .D(n10898), 
            .R(n29060));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_358_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_358_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n29966));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_361_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_1));   // verilog/tli4970.v(54[9:26])
    defparam equal_361_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29965));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29959));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29958));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n28785), .D(n36267), 
            .S(n29060));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n29320));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n29317));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29308));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29301));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_371_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_2));   // verilog/tli4970.v(54[9:26])
    defparam equal_371_i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_363_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3));   // verilog/tli4970.v(54[9:26])
    defparam equal_363_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4617));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n7), 
            .I3(n6_adj_4617), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFNSR delay_counter_2285_2286__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n61[0]), .R(delay_counter_15__N_4494));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2287_2288__i1 (.Q(counter[0]), .C(clk16MHz), .D(n25[0]), 
            .R(clk_slow_N_4413));   // verilog/tli4970.v(14[16:27])
    SB_DFFNE bit_counter_2296__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n28709), 
            .D(n24139));   // verilog/tli4970.v(55[24:39])
    SB_LUT4 mux_2388_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n10898));
    defparam mux_2388_i2_3_lut.LUT_INIT = 16'h3535;
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n28640), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29805));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29781));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n29780));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n29779));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n29778));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n29777));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n29776));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n29775));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n29774));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n29773));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n29772));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n29771));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n29770));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29768));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29763));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29750));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n29741));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29736));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29647));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 bit_counter_2296_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n44215), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2296_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n44214), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2296_add_4_8 (.CI(n44214), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n44215));
    SB_LUT4 bit_counter_2296_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n44213), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2296_add_4_7 (.CI(n44213), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n44214));
    SB_LUT4 bit_counter_2296_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n44212), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2296_add_4_6 (.CI(n44212), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n44213));
    SB_LUT4 bit_counter_2296_add_4_5_lut (.I0(n7796), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n44211), .O(n54245)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2296_add_4_5 (.CI(n44211), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n44212));
    SB_LUT4 bit_counter_2296_add_4_4_lut (.I0(n7796), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n44210), .O(n54244)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2296_add_4_4 (.CI(n44210), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n44211));
    SB_LUT4 bit_counter_2296_add_4_3_lut (.I0(n7796), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n44209), .O(n54243)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2296_add_4_3 (.CI(n44209), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n44210));
    SB_LUT4 bit_counter_2296_add_4_2_lut (.I0(n7796), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n54291)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2296_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2296_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n44209));
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4494), .O(n28785));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfff4;
    SB_LUT4 i14984_2_lut_4_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4494), .O(n29060));
    defparam i14984_2_lut_4_lut.LUT_INIT = 16'h0b00;
    SB_LUT4 equal_371_i7_2_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n7));   // verilog/tli4970.v(54[9:26])
    defparam equal_371_i7_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n27222));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_946 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27287));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_946.LUT_INIT = 16'hbfff;
    SB_LUT4 i2_2_lut_adj_947 (.I0(delay_counter[5]), .I1(delay_counter[6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4618));
    defparam i2_2_lut_adj_947.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(delay_counter[0]), .I1(delay_counter[1]), .I2(delay_counter[3]), 
            .I3(delay_counter[2]), .O(n51100));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_948 (.I0(n51100), .I1(n6_adj_4618), .I2(delay_counter[7]), 
            .I3(delay_counter[4]), .O(n49889));
    defparam i3_4_lut_adj_948.LUT_INIT = 16'hfefc;
    SB_LUT4 i3_4_lut_adj_949 (.I0(n49889), .I1(delay_counter[8]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n49957));
    defparam i3_4_lut_adj_949.LUT_INIT = 16'h8000;
    SB_LUT4 i2397_4_lut (.I0(n49957), .I1(delay_counter[13]), .I2(delay_counter[12]), 
            .I3(delay_counter[11]), .O(delay_counter_15__N_4494));
    defparam i2397_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_2_lut_4_lut_adj_950 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27281));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_950.LUT_INIT = 16'hfbff;
    SB_LUT4 i10069_3_lut (.I0(\state[0] ), .I1(n54243), .I2(\state[1] ), 
            .I3(GND_net), .O(n24112));   // verilog/tli4970.v(55[24:39])
    defparam i10069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10067_3_lut (.I0(\state[0] ), .I1(n54244), .I2(\state[1] ), 
            .I3(GND_net), .O(n24110));   // verilog/tli4970.v(55[24:39])
    defparam i10067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10065_3_lut (.I0(\state[0] ), .I1(n54245), .I2(\state[1] ), 
            .I3(GND_net), .O(n24108));   // verilog/tli4970.v(55[24:39])
    defparam i10065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_951 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27294));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_951.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_952 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n27256));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_952.LUT_INIT = 16'hfffb;
    SB_LUT4 i15004_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29079));   // verilog/tli4970.v(55[24:39])
    defparam i15004_2_lut_2_lut.LUT_INIT = 16'h4444;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1) 
//

module \quadrature_decoder(1)  (encoder1_position, GND_net, VCC_net, b_prev, 
            a_new, position_31__N_4108, ENCODER1_B_N_keep, n2269, ENCODER1_A_N_keep, 
            n29392, n2274) /* synthesis lattice_noprune=1 */ ;
    output [31:0]encoder1_position;
    input GND_net;
    input VCC_net;
    output b_prev;
    output [1:0]a_new;
    output position_31__N_4108;
    input ENCODER1_B_N_keep;
    input n2269;
    input ENCODER1_A_N_keep;
    input n29392;
    output n2274;
    
    
    wire n44198, direction_N_4113, n44199;
    wire [31:0]n133;
    
    wire n44197, n44196, n44195, n44194, n44193, n44192, n44191, 
        n44190, n44189, n44188, n44187, n44186, n44185, n44184, 
        n44183, n44182, n44181, n44180, n44179, n44178, n44177, 
        n44176, n44175, n44174, n44173;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire position_31__N_4111, debounce_cnt, a_prev;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_4116, n29444, n29443, n44203, n44202, n44201, 
        n44200;
    
    SB_CARRY position_2293_add_4_28 (.CI(n44198), .I0(direction_N_4113), 
            .I1(encoder1_position[26]), .CO(n44199));
    SB_LUT4 position_2293_add_4_27_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[25]), .I3(n44197), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_27 (.CI(n44197), .I0(direction_N_4113), 
            .I1(encoder1_position[25]), .CO(n44198));
    SB_LUT4 position_2293_add_4_26_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[24]), .I3(n44196), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_26 (.CI(n44196), .I0(direction_N_4113), 
            .I1(encoder1_position[24]), .CO(n44197));
    SB_LUT4 position_2293_add_4_25_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[23]), .I3(n44195), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_25 (.CI(n44195), .I0(direction_N_4113), 
            .I1(encoder1_position[23]), .CO(n44196));
    SB_LUT4 position_2293_add_4_24_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[22]), .I3(n44194), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_24 (.CI(n44194), .I0(direction_N_4113), 
            .I1(encoder1_position[22]), .CO(n44195));
    SB_LUT4 position_2293_add_4_23_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[21]), .I3(n44193), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_23 (.CI(n44193), .I0(direction_N_4113), 
            .I1(encoder1_position[21]), .CO(n44194));
    SB_LUT4 position_2293_add_4_22_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[20]), .I3(n44192), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_22 (.CI(n44192), .I0(direction_N_4113), 
            .I1(encoder1_position[20]), .CO(n44193));
    SB_LUT4 position_2293_add_4_21_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[19]), .I3(n44191), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_21 (.CI(n44191), .I0(direction_N_4113), 
            .I1(encoder1_position[19]), .CO(n44192));
    SB_LUT4 position_2293_add_4_20_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[18]), .I3(n44190), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_20 (.CI(n44190), .I0(direction_N_4113), 
            .I1(encoder1_position[18]), .CO(n44191));
    SB_LUT4 position_2293_add_4_19_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[17]), .I3(n44189), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_19 (.CI(n44189), .I0(direction_N_4113), 
            .I1(encoder1_position[17]), .CO(n44190));
    SB_LUT4 position_2293_add_4_18_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[16]), .I3(n44188), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_18 (.CI(n44188), .I0(direction_N_4113), 
            .I1(encoder1_position[16]), .CO(n44189));
    SB_LUT4 position_2293_add_4_17_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[15]), .I3(n44187), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_17 (.CI(n44187), .I0(direction_N_4113), 
            .I1(encoder1_position[15]), .CO(n44188));
    SB_LUT4 position_2293_add_4_16_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[14]), .I3(n44186), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_16 (.CI(n44186), .I0(direction_N_4113), 
            .I1(encoder1_position[14]), .CO(n44187));
    SB_LUT4 position_2293_add_4_15_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[13]), .I3(n44185), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_15 (.CI(n44185), .I0(direction_N_4113), 
            .I1(encoder1_position[13]), .CO(n44186));
    SB_LUT4 position_2293_add_4_14_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[12]), .I3(n44184), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_14 (.CI(n44184), .I0(direction_N_4113), 
            .I1(encoder1_position[12]), .CO(n44185));
    SB_LUT4 position_2293_add_4_13_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[11]), .I3(n44183), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_13 (.CI(n44183), .I0(direction_N_4113), 
            .I1(encoder1_position[11]), .CO(n44184));
    SB_LUT4 position_2293_add_4_12_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[10]), .I3(n44182), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_12 (.CI(n44182), .I0(direction_N_4113), 
            .I1(encoder1_position[10]), .CO(n44183));
    SB_LUT4 position_2293_add_4_11_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[9]), .I3(n44181), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_11 (.CI(n44181), .I0(direction_N_4113), 
            .I1(encoder1_position[9]), .CO(n44182));
    SB_LUT4 position_2293_add_4_10_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[8]), .I3(n44180), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_10 (.CI(n44180), .I0(direction_N_4113), 
            .I1(encoder1_position[8]), .CO(n44181));
    SB_LUT4 position_2293_add_4_9_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[7]), .I3(n44179), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_9 (.CI(n44179), .I0(direction_N_4113), 
            .I1(encoder1_position[7]), .CO(n44180));
    SB_LUT4 position_2293_add_4_8_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[6]), .I3(n44178), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_8 (.CI(n44178), .I0(direction_N_4113), 
            .I1(encoder1_position[6]), .CO(n44179));
    SB_LUT4 position_2293_add_4_7_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[5]), .I3(n44177), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_7 (.CI(n44177), .I0(direction_N_4113), 
            .I1(encoder1_position[5]), .CO(n44178));
    SB_LUT4 position_2293_add_4_6_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[4]), .I3(n44176), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_6 (.CI(n44176), .I0(direction_N_4113), 
            .I1(encoder1_position[4]), .CO(n44177));
    SB_LUT4 position_2293_add_4_5_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[3]), .I3(n44175), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_5 (.CI(n44175), .I0(direction_N_4113), 
            .I1(encoder1_position[3]), .CO(n44176));
    SB_LUT4 position_2293_add_4_4_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[2]), .I3(n44174), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_4 (.CI(n44174), .I0(direction_N_4113), 
            .I1(encoder1_position[2]), .CO(n44175));
    SB_LUT4 position_2293_add_4_3_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[1]), .I3(n44173), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_3 (.CI(n44173), .I0(direction_N_4113), 
            .I1(encoder1_position[1]), .CO(n44174));
    SB_LUT4 position_2293_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n44173));
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_4111));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_4111), 
            .I3(a_new[1]), .O(position_31__N_4108));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 i39817_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_4116));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i39817_4_lut.LUT_INIT = 16'h8421;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n2269), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n2269), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n2269), .D(a_prev_N_4116));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n2274), .C(n2269), .D(n29392));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2293__i31 (.Q(encoder1_position[31]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i30 (.Q(encoder1_position[30]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i29 (.Q(encoder1_position[29]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i28 (.Q(encoder1_position[28]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i27 (.Q(encoder1_position[27]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i26 (.Q(encoder1_position[26]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i25 (.Q(encoder1_position[25]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i24 (.Q(encoder1_position[24]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i23 (.Q(encoder1_position[23]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i22 (.Q(encoder1_position[22]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i21 (.Q(encoder1_position[21]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i20 (.Q(encoder1_position[20]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i19 (.Q(encoder1_position[19]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i18 (.Q(encoder1_position[18]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i17 (.Q(encoder1_position[17]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i16 (.Q(encoder1_position[16]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i15 (.Q(encoder1_position[15]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i14 (.Q(encoder1_position[14]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i13 (.Q(encoder1_position[13]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i12 (.Q(encoder1_position[12]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i11 (.Q(encoder1_position[11]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i10 (.Q(encoder1_position[10]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i9 (.Q(encoder1_position[9]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i8 (.Q(encoder1_position[8]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i7 (.Q(encoder1_position[7]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i6 (.Q(encoder1_position[6]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i5 (.Q(encoder1_position[5]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i4 (.Q(encoder1_position[4]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i3 (.Q(encoder1_position[3]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i2 (.Q(encoder1_position[2]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i1 (.Q(encoder1_position[1]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2293__i0 (.Q(encoder1_position[0]), .C(n2269), .E(position_31__N_4108), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_4113));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n2269), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n2269), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i15368_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4116), .I2(a_new[1]), 
            .I3(a_prev), .O(n29444));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15368_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15367_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_4116), .I2(b_new[1]), 
            .I3(b_prev), .O(n29443));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 position_2293_add_4_33_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[31]), .I3(n44203), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2293_add_4_32_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[30]), .I3(n44202), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_32 (.CI(n44202), .I0(direction_N_4113), 
            .I1(encoder1_position[30]), .CO(n44203));
    SB_DFF a_prev_38 (.Q(a_prev), .C(n2269), .D(n29444));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n2269), .D(n29443));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2293_add_4_31_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[29]), .I3(n44201), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_31 (.CI(n44201), .I0(direction_N_4113), 
            .I1(encoder1_position[29]), .CO(n44202));
    SB_LUT4 position_2293_add_4_30_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[28]), .I3(n44200), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_30 (.CI(n44200), .I0(direction_N_4113), 
            .I1(encoder1_position[28]), .CO(n44201));
    SB_LUT4 position_2293_add_4_29_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[27]), .I3(n44199), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2293_add_4_29 (.CI(n44199), .I0(direction_N_4113), 
            .I1(encoder1_position[27]), .CO(n44200));
    SB_LUT4 position_2293_add_4_28_lut (.I0(GND_net), .I1(direction_N_4113), 
            .I2(encoder1_position[26]), .I3(n44198), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2293_add_4_28_lut.LUT_INIT = 16'hC33C;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (pwm_out, clk32MHz, GND_net, VCC_net, pwm_setpoint) /* synthesis syn_module_defined=1 */ ;
    output pwm_out;
    input clk32MHz;
    input GND_net;
    input VCC_net;
    input [23:0]pwm_setpoint;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire pwm_out_N_908;
    wire [23:0]n101;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire pwm_counter_23__N_906, n44078, n44077, n44076, n44075, n44074, 
        n44073, n44072, n44071, n44070, n44069, n44068, n44067, 
        n44066, n44065, n44064, n44063, n44062, n44061, n44060, 
        n44059, n44058, n44057, n44056, n8, n54642, n16, n10, 
        n54653, n12, n54676, n6, n39, n41, n45, n43, n37, 
        n29, n31, n23, n25, n35, n33, n11, n13, n15, n27, 
        n9, n17, n19, n21, n54666, n54660, n30, n55059, n55055, 
        n55452, n55233, n55498, n55324, n55325, n24, n54644, n55133, 
        n54810, n4, n55322, n55323, n54655, n55456, n54812, n55540, 
        n55541, n55529, n54646, n55388, n54818, n55478, n51181, 
        n22, n15_adj_4610, n20, n24_adj_4611, n19_adj_4612;
    
    SB_DFF pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .D(pwm_out_N_908));   // verilog/pwm.v(16[12] 26[6])
    SB_DFFSR pwm_counter_2282__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n101[23]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n101[22]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n101[21]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n101[20]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n101[19]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n101[18]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n101[17]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n101[16]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n101[15]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n101[14]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n101[13]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n101[12]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n101[11]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n101[10]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n101[9]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n101[8]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n101[7]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n101[6]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n101[5]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n101[4]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n101[3]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n101[2]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2282__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n101[1]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_2282_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n44078), .O(n101[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_2282_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n44077), .O(n101[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_24 (.CI(n44077), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n44078));
    SB_LUT4 pwm_counter_2282_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n44076), .O(n101[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_23 (.CI(n44076), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n44077));
    SB_LUT4 pwm_counter_2282_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n44075), .O(n101[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_22 (.CI(n44075), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n44076));
    SB_LUT4 pwm_counter_2282_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n44074), .O(n101[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_21 (.CI(n44074), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n44075));
    SB_LUT4 pwm_counter_2282_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n44073), .O(n101[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_20 (.CI(n44073), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n44074));
    SB_LUT4 pwm_counter_2282_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n44072), .O(n101[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_19 (.CI(n44072), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n44073));
    SB_LUT4 pwm_counter_2282_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n44071), .O(n101[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_18 (.CI(n44071), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n44072));
    SB_LUT4 pwm_counter_2282_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n44070), .O(n101[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_17 (.CI(n44070), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n44071));
    SB_LUT4 pwm_counter_2282_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n44069), .O(n101[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_16 (.CI(n44069), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n44070));
    SB_LUT4 pwm_counter_2282_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n44068), .O(n101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_15 (.CI(n44068), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n44069));
    SB_LUT4 pwm_counter_2282_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n44067), .O(n101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_14 (.CI(n44067), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n44068));
    SB_LUT4 pwm_counter_2282_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n44066), .O(n101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_13 (.CI(n44066), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n44067));
    SB_LUT4 pwm_counter_2282_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n44065), .O(n101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_12 (.CI(n44065), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n44066));
    SB_LUT4 pwm_counter_2282_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n44064), .O(n101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_11 (.CI(n44064), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n44065));
    SB_LUT4 pwm_counter_2282_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n44063), .O(n101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_10 (.CI(n44063), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n44064));
    SB_LUT4 pwm_counter_2282_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n44062), .O(n101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_9 (.CI(n44062), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n44063));
    SB_LUT4 pwm_counter_2282_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n44061), .O(n101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_8 (.CI(n44061), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n44062));
    SB_LUT4 pwm_counter_2282_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n44060), .O(n101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_7 (.CI(n44060), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n44061));
    SB_LUT4 pwm_counter_2282_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n44059), .O(n101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_6 (.CI(n44059), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n44060));
    SB_LUT4 pwm_counter_2282_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n44058), .O(n101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_5 (.CI(n44058), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n44059));
    SB_LUT4 pwm_counter_2282_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n44057), .O(n101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_4 (.CI(n44057), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n44058));
    SB_LUT4 pwm_counter_2282_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n44056), .O(n101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_3 (.CI(n44056), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n44057));
    SB_LUT4 pwm_counter_2282_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2282_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2282_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n44056));
    SB_DFFSR pwm_counter_2282__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n101[0]), 
            .R(pwm_counter_23__N_906));   // verilog/pwm.v(17[20:33])
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38849_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n54642));
    defparam i38849_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38860_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n54653));
    defparam i38860_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i38883_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n54676));   // verilog/pwm.v(21[8:24])
    defparam i38883_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38873_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n54666));
    defparam i38873_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i38867_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n54660));
    defparam i38867_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39266_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n54676), 
            .O(n55059));
    defparam i39266_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39262_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n55059), 
            .O(n55055));
    defparam i39262_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i39659_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n55055), 
            .O(n55452));
    defparam i39659_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39440_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n55452), 
            .O(n55233));
    defparam i39440_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i39705_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n55233), 
            .O(n55498));
    defparam i39705_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i39531_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n55324));   // verilog/pwm.v(21[8:24])
    defparam i39531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39532_3_lut (.I0(n55324), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n55325));   // verilog/pwm.v(21[8:24])
    defparam i39532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38851_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n54666), 
            .O(n54644));
    defparam i38851_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39340_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n54642), 
            .O(n55133));   // verilog/pwm.v(21[8:24])
    defparam i39340_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39017_3_lut (.I0(n55325), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n54810));   // verilog/pwm.v(21[8:24])
    defparam i39017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i39529_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n55322));   // verilog/pwm.v(21[8:24])
    defparam i39529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39530_3_lut (.I0(n55322), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n55323));   // verilog/pwm.v(21[8:24])
    defparam i39530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38862_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n54660), 
            .O(n54655));
    defparam i38862_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39663_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n54653), 
            .O(n55456));   // verilog/pwm.v(21[8:24])
    defparam i39663_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i39019_3_lut (.I0(n55323), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n54812));   // verilog/pwm.v(21[8:24])
    defparam i39019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39747_4_lut (.I0(n54812), .I1(n55456), .I2(n35), .I3(n54655), 
            .O(n55540));   // verilog/pwm.v(21[8:24])
    defparam i39747_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39748_3_lut (.I0(n55540), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n55541));   // verilog/pwm.v(21[8:24])
    defparam i39748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39736_3_lut (.I0(n55541), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n55529));   // verilog/pwm.v(21[8:24])
    defparam i39736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38853_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n55498), 
            .O(n54646));
    defparam i38853_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i39595_4_lut (.I0(n54810), .I1(n55133), .I2(n45), .I3(n54644), 
            .O(n55388));   // verilog/pwm.v(21[8:24])
    defparam i39595_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39025_3_lut (.I0(n55529), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n54818));   // verilog/pwm.v(21[8:24])
    defparam i39025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39685_4_lut (.I0(n54818), .I1(n55388), .I2(n45), .I3(n54646), 
            .O(n55478));   // verilog/pwm.v(21[8:24])
    defparam i39685_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39686_3_lut (.I0(n55478), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_908));   // verilog/pwm.v(21[8:24])
    defparam i39686_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n51181));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[16]), .I1(pwm_counter[14]), .I2(pwm_counter[19]), 
            .I3(pwm_counter[17]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n51181), .I1(pwm_counter[22]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15_adj_4610));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[13]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15_adj_4610), .I1(n22), .I2(pwm_counter[15]), 
            .I3(pwm_counter[18]), .O(n24_adj_4611));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[12]), .I1(pwm_counter[20]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4612));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i40493_4_lut (.I0(pwm_counter[23]), .I1(n19_adj_4612), .I2(n24_adj_4611), 
            .I3(n20), .O(pwm_counter_23__N_906));   // verilog/pwm.v(18[8:40])
    defparam i40493_4_lut.LUT_INIT = 16'h5554;
    
endmodule
