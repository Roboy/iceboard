-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Mar 24 2020 18:54:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : in std_logic;
    SPI_IO2 : in std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : in std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : out std_logic;
    PIN_19 : in std_logic;
    PIN_18 : out std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : inout std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : in std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \uart.n2132\ : std_logic;
signal \uart.n2133\ : std_logic;
signal \uart.n2134\ : std_logic;
signal \uart.n2135\ : std_logic;
signal \uart.n2136\ : std_logic;
signal \uart.n2137\ : std_logic;
signal \uart.n2138\ : std_logic;
signal \uart.n2139\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \uart.n2140\ : std_logic;
signal \uart.n2141\ : std_logic;
signal \uart.n2142\ : std_logic;
signal \uart.n2143\ : std_logic;
signal \uart.n2144\ : std_logic;
signal \uart.n2145\ : std_logic;
signal \uart.n2146\ : std_logic;
signal \uart.n2147\ : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal \uart.n2148\ : std_logic;
signal \uart.n2149\ : std_logic;
signal \uart.n2150\ : std_logic;
signal \uart.n2151\ : std_logic;
signal \uart.n2152\ : std_logic;
signal \uart.n2153\ : std_logic;
signal \uart.n2154\ : std_logic;
signal \uart.n2155\ : std_logic;
signal \bfn_1_21_0_\ : std_logic;
signal \uart.n2156\ : std_logic;
signal \uart.n2157\ : std_logic;
signal \uart.n2158\ : std_logic;
signal \uart.n2159\ : std_logic;
signal \uart.n2160\ : std_logic;
signal \uart.n2161\ : std_logic;
signal \uart.n2162\ : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal n2226 : std_logic;
signal n2227 : std_logic;
signal n2228 : std_logic;
signal n2229 : std_logic;
signal n2230 : std_logic;
signal n2231 : std_logic;
signal n2232 : std_logic;
signal n2233 : std_logic;
signal \bfn_1_23_0_\ : std_logic;
signal n2234 : std_logic;
signal n2235 : std_logic;
signal n2236 : std_logic;
signal n2237 : std_logic;
signal n2238 : std_logic;
signal n2239 : std_logic;
signal n2240 : std_logic;
signal n2241 : std_logic;
signal \bfn_1_24_0_\ : std_logic;
signal n2242 : std_logic;
signal n2243 : std_logic;
signal n2244 : std_logic;
signal n2245 : std_logic;
signal n2246 : std_logic;
signal n2247 : std_logic;
signal n2248 : std_logic;
signal n2249 : std_logic;
signal \bfn_1_25_0_\ : std_logic;
signal n2250 : std_logic;
signal n2251 : std_logic;
signal n2252 : std_logic;
signal n2253 : std_logic;
signal n2254 : std_logic;
signal n2255 : std_logic;
signal n2256 : std_logic;
signal \uart.r_Clock_Count_2\ : std_logic;
signal \uart.r_Clock_Count_0\ : std_logic;
signal \uart.r_Clock_Count_1\ : std_logic;
signal \uart.r_Clock_Count_3\ : std_logic;
signal \uart.r_Clock_Count_5\ : std_logic;
signal \uart.r_Clock_Count_4\ : std_logic;
signal \uart.n2006_cascade_\ : std_logic;
signal \uart.r_Clock_Count_6\ : std_logic;
signal \uart.r_Clock_Count_10\ : std_logic;
signal \uart.r_Clock_Count_22\ : std_logic;
signal \uart.r_Clock_Count_26\ : std_logic;
signal \uart.r_Clock_Count_13\ : std_logic;
signal \uart.r_Clock_Count_12\ : std_logic;
signal \uart.r_Clock_Count_29\ : std_logic;
signal \uart.n42_cascade_\ : std_logic;
signal \uart.r_Clock_Count_7\ : std_logic;
signal \uart.n45_cascade_\ : std_logic;
signal \uart.n2385\ : std_logic;
signal \r_SM_Main_2_N_233_1_cascade_\ : std_logic;
signal \uart.n1796\ : std_logic;
signal \uart.r_Clock_Count_8\ : std_logic;
signal \uart.r_Clock_Count_14\ : std_logic;
signal \uart.n34\ : std_logic;
signal \uart.r_Clock_Count_30\ : std_logic;
signal \uart.r_Clock_Count_28\ : std_logic;
signal \uart.r_Clock_Count_24\ : std_logic;
signal \uart.r_Clock_Count_23\ : std_logic;
signal \uart.n1\ : std_logic;
signal \uart.r_Clock_Count_11\ : std_logic;
signal \uart.r_Clock_Count_21\ : std_logic;
signal \uart.r_Clock_Count_17\ : std_logic;
signal \uart.r_Clock_Count_18\ : std_logic;
signal \uart.r_Clock_Count_20\ : std_logic;
signal \uart.r_Clock_Count_15\ : std_logic;
signal \uart.r_Clock_Count_25\ : std_logic;
signal \uart.r_Clock_Count_9\ : std_logic;
signal \uart.r_Clock_Count_27\ : std_logic;
signal \uart.r_Clock_Count_19\ : std_logic;
signal \uart.r_Clock_Count_16\ : std_logic;
signal \uart.r_Clock_Count_31\ : std_logic;
signal \uart.n39\ : std_logic;
signal \uart.n40\ : std_logic;
signal \uart.n37_cascade_\ : std_logic;
signal \uart.n38\ : std_logic;
signal \uart.n46\ : std_logic;
signal clk_divider_26 : std_logic;
signal clk_divider_9 : std_logic;
signal clk_divider_14 : std_logic;
signal clk_divider_17 : std_logic;
signal clk_divider_21 : std_logic;
signal clk_divider_22 : std_logic;
signal clk_divider_28 : std_logic;
signal clk_divider_6 : std_logic;
signal clk_divider_30 : std_logic;
signal clk_divider_27 : std_logic;
signal clk_divider_20 : std_logic;
signal clk_divider_19 : std_logic;
signal n44_adj_358 : std_logic;
signal \n42_adj_360_cascade_\ : std_logic;
signal n41_adj_361 : std_logic;
signal clk_divider_4 : std_logic;
signal clk_divider_0 : std_logic;
signal clk_divider_3 : std_logic;
signal \clk_divider_31__N_139\ : std_logic;
signal \uart.n3\ : std_logic;
signal clk_divider_1 : std_logic;
signal clk_divider_2 : std_logic;
signal n6_adj_324 : std_logic;
signal clk_divider_8 : std_logic;
signal clk_divider_15 : std_logic;
signal clk_divider_24 : std_logic;
signal clk_divider_11 : std_logic;
signal clk_divider_5 : std_logic;
signal clk_divider_10 : std_logic;
signal clk_divider_12 : std_logic;
signal clk_divider_18 : std_logic;
signal clk_divider_13 : std_logic;
signal clk_divider_29 : std_logic;
signal clk_divider_23 : std_logic;
signal clk_divider_16 : std_logic;
signal n43_adj_359 : std_logic;
signal clk_divider_31 : std_logic;
signal n50 : std_logic;
signal n10 : std_logic;
signal n26 : std_logic;
signal \bfn_2_23_0_\ : std_logic;
signal n25 : std_logic;
signal n2163 : std_logic;
signal n24 : std_logic;
signal n2164 : std_logic;
signal n23 : std_logic;
signal n2165 : std_logic;
signal n22 : std_logic;
signal n2166 : std_logic;
signal n21 : std_logic;
signal n2167 : std_logic;
signal n20 : std_logic;
signal n2168 : std_logic;
signal n19 : std_logic;
signal n2169 : std_logic;
signal n2170 : std_logic;
signal n18 : std_logic;
signal \bfn_2_24_0_\ : std_logic;
signal n17 : std_logic;
signal n2171 : std_logic;
signal n16 : std_logic;
signal n2172 : std_logic;
signal n15 : std_logic;
signal n2173 : std_logic;
signal n14 : std_logic;
signal n2174 : std_logic;
signal n13 : std_logic;
signal n2175 : std_logic;
signal n12 : std_logic;
signal n2176 : std_logic;
signal n11 : std_logic;
signal n2177 : std_logic;
signal n2178 : std_logic;
signal n10_adj_317 : std_logic;
signal \bfn_2_25_0_\ : std_logic;
signal n9 : std_logic;
signal n2179 : std_logic;
signal n8 : std_logic;
signal n2180 : std_logic;
signal n7 : std_logic;
signal n2181 : std_logic;
signal n6 : std_logic;
signal n2182 : std_logic;
signal n2183 : std_logic;
signal n2184 : std_logic;
signal n2185 : std_logic;
signal n2186 : std_logic;
signal \bfn_2_26_0_\ : std_logic;
signal n2187 : std_logic;
signal blink_counter_25 : std_logic;
signal \n2395_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal blink_counter_21 : std_logic;
signal blink_counter_24 : std_logic;
signal blink_counter_23 : std_logic;
signal blink_counter_22 : std_logic;
signal n2394 : std_logic;
signal \uart.n1711\ : std_logic;
signal \uart.o_Tx_Serial_N_312\ : std_logic;
signal clk_divider_7 : std_logic;
signal n40_adj_362 : std_logic;
signal clk_divider_25 : std_logic;
signal n45_adj_357 : std_logic;
signal n49 : std_logic;
signal counter_0 : std_logic;
signal \bfn_3_22_0_\ : std_logic;
signal counter_1 : std_logic;
signal n2195 : std_logic;
signal counter_2 : std_logic;
signal n2196 : std_logic;
signal counter_3 : std_logic;
signal n2197 : std_logic;
signal counter_4 : std_logic;
signal n2198 : std_logic;
signal counter_5 : std_logic;
signal n2199 : std_logic;
signal counter_6 : std_logic;
signal n2200 : std_logic;
signal counter_7 : std_logic;
signal n2201 : std_logic;
signal n2202 : std_logic;
signal \bfn_3_23_0_\ : std_logic;
signal n2203 : std_logic;
signal n2204 : std_logic;
signal n2205 : std_logic;
signal n2206 : std_logic;
signal n2207 : std_logic;
signal n2208 : std_logic;
signal n2209 : std_logic;
signal n2210 : std_logic;
signal \bfn_3_24_0_\ : std_logic;
signal n2211 : std_logic;
signal n2212 : std_logic;
signal n2213 : std_logic;
signal n2214 : std_logic;
signal n2215 : std_logic;
signal n2216 : std_logic;
signal n2217 : std_logic;
signal n2218 : std_logic;
signal \bfn_3_25_0_\ : std_logic;
signal n2219 : std_logic;
signal n2220 : std_logic;
signal n2221 : std_logic;
signal n2222 : std_logic;
signal n2223 : std_logic;
signal n2224 : std_logic;
signal n2225 : std_logic;
signal \uart.r_Bit_Index_2\ : std_logic;
signal \n2002_cascade_\ : std_logic;
signal \r_SM_Main_2_N_233_1\ : std_logic;
signal \n2308_cascade_\ : std_logic;
signal n2002 : std_logic;
signal \uart.n2428_cascade_\ : std_logic;
signal \uart.n2431\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \uart.n2422_cascade_\ : std_logic;
signal \uart.n2425\ : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal n1757 : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal data_out_5 : std_logic;
signal data_out_0 : std_logic;
signal data_out_3 : std_logic;
signal data_out_1 : std_logic;
signal data_out_2 : std_logic;
signal counter_13 : std_logic;
signal counter_23 : std_logic;
signal counter_11 : std_logic;
signal counter_14 : std_logic;
signal \n38_cascade_\ : std_logic;
signal \n44_cascade_\ : std_logic;
signal \counter_31__N_172_cascade_\ : std_logic;
signal data_out_4 : std_logic;
signal counter_31 : std_logic;
signal n44 : std_logic;
signal \r_SM_Main_2_N_236_0\ : std_logic;
signal data_out_6 : std_logic;
signal counter_22 : std_logic;
signal counter_30 : std_logic;
signal counter_19 : std_logic;
signal counter_26 : std_logic;
signal n36 : std_logic;
signal counter_12 : std_logic;
signal counter_8 : std_logic;
signal counter_15 : std_logic;
signal counter_25 : std_logic;
signal n40 : std_logic;
signal counter_17 : std_logic;
signal counter_24 : std_logic;
signal counter_21 : std_logic;
signal counter_16 : std_logic;
signal n39 : std_logic;
signal counter_20 : std_logic;
signal counter_10 : std_logic;
signal counter_29 : std_logic;
signal counter_28 : std_logic;
signal n37 : std_logic;
signal counter_18 : std_logic;
signal counter_27 : std_logic;
signal counter_9 : std_logic;
signal n35 : std_logic;
signal data_out_7 : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \uart.r_Bit_Index_1\ : std_logic;
signal \CLK_c\ : std_logic;
signal n2308 : std_logic;
signal \uart.n2310\ : std_logic;
signal diff_input : std_logic;
signal integrator_0 : std_logic;
signal \bfn_5_23_0_\ : std_logic;
signal integrator_1 : std_logic;
signal n2188 : std_logic;
signal integrator_2 : std_logic;
signal n2189 : std_logic;
signal integrator_3 : std_logic;
signal n2190 : std_logic;
signal integrator_4 : std_logic;
signal n2191 : std_logic;
signal integrator_5 : std_logic;
signal n2192 : std_logic;
signal integrator_6 : std_logic;
signal n2193 : std_logic;
signal n2194 : std_logic;
signal integrator_7 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_slow : std_logic;
signal \counter_31__N_172\ : std_logic;

signal \LED_wire\ : std_logic;
signal \PIN_18_wire\ : std_logic;
signal \PIN_2_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    PIN_18 <= \PIN_18_wire\;
    PIN_2 <= \PIN_2_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5970\,
            DIN => \N__5969\,
            DOUT => \N__5968\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5970\,
            PADOUT => \N__5969\,
            PADIN => \N__5968\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4358\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_18_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5961\,
            DIN => \N__5960\,
            DOUT => \N__5959\,
            PACKAGEPIN => \PIN_18_wire\
        );

    \PIN_18_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5961\,
            PADOUT => \N__5960\,
            PADIN => \N__5959\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5276\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__5825\,
            OUTPUTENABLE => '0'
        );

    \PIN_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5952\,
            DIN => \N__5951\,
            DOUT => \N__5950\,
            PACKAGEPIN => \PIN_2_wire\
        );

    \PIN_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5952\,
            PADOUT => \N__5951\,
            PADIN => \N__5950\,
            CLOCKENABLE => \N__3107\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3911\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__5399\,
            OUTPUTENABLE => '0'
        );

    \differential_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVDS_INPUT",
            PULLUP => '0'
        )
    port map (
            OE => \N__5943\,
            DIN => \N__5942\,
            DOUT => \N__5941\,
            PACKAGEPIN => PIN_13
        );

    \differential_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5943\,
            PADOUT => \N__5942\,
            PADIN => \N__5941\,
            CLOCKENABLE => 'H',
            DIN0 => diff_input,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5934\,
            DIN => \N__5933\,
            DOUT => \N__5932\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5934\,
            PADOUT => \N__5933\,
            PADIN => \N__5932\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__1307\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5911\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5908\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__5911\,
            I => integrator_2
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5908\,
            I => integrator_2
        );

    \I__1303\ : InMux
    port map (
            O => \N__5903\,
            I => n2189
        );

    \I__1302\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5896\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5899\,
            I => \N__5893\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5896\,
            I => integrator_3
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5893\,
            I => integrator_3
        );

    \I__1298\ : InMux
    port map (
            O => \N__5888\,
            I => n2190
        );

    \I__1297\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5881\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5878\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__5881\,
            I => integrator_4
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__5878\,
            I => integrator_4
        );

    \I__1293\ : InMux
    port map (
            O => \N__5873\,
            I => n2191
        );

    \I__1292\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5866\
        );

    \I__1291\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5863\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5866\,
            I => integrator_5
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5863\,
            I => integrator_5
        );

    \I__1288\ : InMux
    port map (
            O => \N__5858\,
            I => n2192
        );

    \I__1287\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5851\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5848\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5851\,
            I => integrator_6
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5848\,
            I => integrator_6
        );

    \I__1283\ : InMux
    port map (
            O => \N__5843\,
            I => n2193
        );

    \I__1282\ : InMux
    port map (
            O => \N__5840\,
            I => n2194
        );

    \I__1281\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5833\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5830\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5833\,
            I => integrator_7
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5830\,
            I => integrator_7
        );

    \I__1277\ : ClkMux
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5822\,
            I => \N__5819\
        );

    \I__1275\ : Span4Mux_s2_h
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__1274\ : Span4Mux_h
    port map (
            O => \N__5816\,
            I => \N__5809\
        );

    \I__1273\ : ClkMux
    port map (
            O => \N__5815\,
            I => \N__5806\
        );

    \I__1272\ : ClkMux
    port map (
            O => \N__5814\,
            I => \N__5801\
        );

    \I__1271\ : ClkMux
    port map (
            O => \N__5813\,
            I => \N__5798\
        );

    \I__1270\ : ClkMux
    port map (
            O => \N__5812\,
            I => \N__5795\
        );

    \I__1269\ : Sp12to4
    port map (
            O => \N__5809\,
            I => \N__5792\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__5806\,
            I => \N__5789\
        );

    \I__1267\ : ClkMux
    port map (
            O => \N__5805\,
            I => \N__5786\
        );

    \I__1266\ : ClkMux
    port map (
            O => \N__5804\,
            I => \N__5783\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5801\,
            I => \N__5780\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5798\,
            I => \N__5775\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5795\,
            I => \N__5775\
        );

    \I__1262\ : Span12Mux_v
    port map (
            O => \N__5792\,
            I => \N__5771\
        );

    \I__1261\ : Span4Mux_v
    port map (
            O => \N__5789\,
            I => \N__5766\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5786\,
            I => \N__5766\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5783\,
            I => \N__5763\
        );

    \I__1258\ : Span4Mux_v
    port map (
            O => \N__5780\,
            I => \N__5758\
        );

    \I__1257\ : Span4Mux_v
    port map (
            O => \N__5775\,
            I => \N__5758\
        );

    \I__1256\ : ClkMux
    port map (
            O => \N__5774\,
            I => \N__5755\
        );

    \I__1255\ : Span12Mux_h
    port map (
            O => \N__5771\,
            I => \N__5751\
        );

    \I__1254\ : Span4Mux_h
    port map (
            O => \N__5766\,
            I => \N__5748\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__5763\,
            I => \N__5745\
        );

    \I__1252\ : Span4Mux_s2_h
    port map (
            O => \N__5758\,
            I => \N__5740\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5755\,
            I => \N__5740\
        );

    \I__1250\ : ClkMux
    port map (
            O => \N__5754\,
            I => \N__5737\
        );

    \I__1249\ : Span12Mux_h
    port map (
            O => \N__5751\,
            I => \N__5734\
        );

    \I__1248\ : Span4Mux_v
    port map (
            O => \N__5748\,
            I => \N__5731\
        );

    \I__1247\ : Sp12to4
    port map (
            O => \N__5745\,
            I => \N__5724\
        );

    \I__1246\ : Sp12to4
    port map (
            O => \N__5740\,
            I => \N__5724\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5737\,
            I => \N__5724\
        );

    \I__1244\ : Odrv12
    port map (
            O => \N__5734\,
            I => clk_slow
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__5731\,
            I => clk_slow
        );

    \I__1242\ : Odrv12
    port map (
            O => \N__5724\,
            I => clk_slow
        );

    \I__1241\ : SRMux
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__1239\ : Span4Mux_s3_h
    port map (
            O => \N__5711\,
            I => \N__5697\
        );

    \I__1238\ : SRMux
    port map (
            O => \N__5710\,
            I => \N__5694\
        );

    \I__1237\ : SRMux
    port map (
            O => \N__5709\,
            I => \N__5691\
        );

    \I__1236\ : SRMux
    port map (
            O => \N__5708\,
            I => \N__5688\
        );

    \I__1235\ : SRMux
    port map (
            O => \N__5707\,
            I => \N__5685\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5682\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5675\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5704\,
            I => \N__5675\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5675\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5668\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5668\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5668\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__5697\,
            I => \counter_31__N_172\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5694\,
            I => \counter_31__N_172\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5691\,
            I => \counter_31__N_172\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5688\,
            I => \counter_31__N_172\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5685\,
            I => \counter_31__N_172\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5682\,
            I => \counter_31__N_172\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5675\,
            I => \counter_31__N_172\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5668\,
            I => \counter_31__N_172\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5647\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5644\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__5647\,
            I => counter_17
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5644\,
            I => counter_17
        );

    \I__1215\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5635\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5632\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5635\,
            I => counter_24
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5632\,
            I => counter_24
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__5627\,
            I => \N__5623\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5620\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5617\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5620\,
            I => counter_21
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__5617\,
            I => counter_21
        );

    \I__1206\ : InMux
    port map (
            O => \N__5612\,
            I => \N__5608\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5605\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5608\,
            I => counter_16
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5605\,
            I => counter_16
        );

    \I__1202\ : InMux
    port map (
            O => \N__5600\,
            I => \N__5594\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5594\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5594\,
            I => n39
        );

    \I__1199\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5587\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5584\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5587\,
            I => counter_20
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5584\,
            I => counter_20
        );

    \I__1195\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5575\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5572\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5575\,
            I => counter_10
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5572\,
            I => counter_10
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__5567\,
            I => \N__5563\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5560\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5557\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5560\,
            I => counter_29
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5557\,
            I => counter_29
        );

    \I__1186\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5548\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5545\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5548\,
            I => counter_28
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5545\,
            I => counter_28
        );

    \I__1182\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5537\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5537\,
            I => n37
        );

    \I__1180\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5530\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5527\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5530\,
            I => counter_18
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5527\,
            I => counter_18
        );

    \I__1176\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5518\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5515\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5518\,
            I => counter_27
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5515\,
            I => counter_27
        );

    \I__1172\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5506\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5503\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5506\,
            I => counter_9
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5503\,
            I => counter_9
        );

    \I__1168\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5495\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5495\,
            I => n35
        );

    \I__1166\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5489\,
            I => \N__5485\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5482\
        );

    \I__1163\ : Odrv12
    port map (
            O => \N__5485\,
            I => data_out_7
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__5482\,
            I => data_out_7
        );

    \I__1161\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5469\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5466\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5461\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5461\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5456\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5456\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__5469\,
            I => \r_Bit_Index_0\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5466\,
            I => \r_Bit_Index_0\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5461\,
            I => \r_Bit_Index_0\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5456\,
            I => \r_Bit_Index_0\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5444\,
            I => \N__5439\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__5443\,
            I => \N__5433\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__5442\,
            I => \N__5429\
        );

    \I__1147\ : Span4Mux_h
    port map (
            O => \N__5439\,
            I => \N__5426\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5423\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5437\,
            I => \N__5420\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5415\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5415\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5410\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5410\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__5426\,
            I => \uart.r_Bit_Index_1\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5423\,
            I => \uart.r_Bit_Index_1\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5420\,
            I => \uart.r_Bit_Index_1\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5415\,
            I => \uart.r_Bit_Index_1\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5410\,
            I => \uart.r_Bit_Index_1\
        );

    \I__1135\ : ClkMux
    port map (
            O => \N__5399\,
            I => \N__5336\
        );

    \I__1134\ : ClkMux
    port map (
            O => \N__5398\,
            I => \N__5336\
        );

    \I__1133\ : ClkMux
    port map (
            O => \N__5397\,
            I => \N__5336\
        );

    \I__1132\ : ClkMux
    port map (
            O => \N__5396\,
            I => \N__5336\
        );

    \I__1131\ : ClkMux
    port map (
            O => \N__5395\,
            I => \N__5336\
        );

    \I__1130\ : ClkMux
    port map (
            O => \N__5394\,
            I => \N__5336\
        );

    \I__1129\ : ClkMux
    port map (
            O => \N__5393\,
            I => \N__5336\
        );

    \I__1128\ : ClkMux
    port map (
            O => \N__5392\,
            I => \N__5336\
        );

    \I__1127\ : ClkMux
    port map (
            O => \N__5391\,
            I => \N__5336\
        );

    \I__1126\ : ClkMux
    port map (
            O => \N__5390\,
            I => \N__5336\
        );

    \I__1125\ : ClkMux
    port map (
            O => \N__5389\,
            I => \N__5336\
        );

    \I__1124\ : ClkMux
    port map (
            O => \N__5388\,
            I => \N__5336\
        );

    \I__1123\ : ClkMux
    port map (
            O => \N__5387\,
            I => \N__5336\
        );

    \I__1122\ : ClkMux
    port map (
            O => \N__5386\,
            I => \N__5336\
        );

    \I__1121\ : ClkMux
    port map (
            O => \N__5385\,
            I => \N__5336\
        );

    \I__1120\ : ClkMux
    port map (
            O => \N__5384\,
            I => \N__5336\
        );

    \I__1119\ : ClkMux
    port map (
            O => \N__5383\,
            I => \N__5336\
        );

    \I__1118\ : ClkMux
    port map (
            O => \N__5382\,
            I => \N__5336\
        );

    \I__1117\ : ClkMux
    port map (
            O => \N__5381\,
            I => \N__5336\
        );

    \I__1116\ : ClkMux
    port map (
            O => \N__5380\,
            I => \N__5336\
        );

    \I__1115\ : ClkMux
    port map (
            O => \N__5379\,
            I => \N__5336\
        );

    \I__1114\ : GlobalMux
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__1113\ : gio2CtrlBuf
    port map (
            O => \N__5333\,
            I => \CLK_c\
        );

    \I__1112\ : CEMux
    port map (
            O => \N__5330\,
            I => \N__5326\
        );

    \I__1111\ : CEMux
    port map (
            O => \N__5329\,
            I => \N__5323\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5326\,
            I => \N__5320\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__5323\,
            I => \N__5316\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__5320\,
            I => \N__5313\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5319\,
            I => \N__5310\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__5316\,
            I => n2308
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__5313\,
            I => n2308
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5310\,
            I => n2308
        );

    \I__1103\ : SRMux
    port map (
            O => \N__5303\,
            I => \N__5299\
        );

    \I__1102\ : SRMux
    port map (
            O => \N__5302\,
            I => \N__5296\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5299\,
            I => \N__5293\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5296\,
            I => \N__5290\
        );

    \I__1099\ : Span4Mux_h
    port map (
            O => \N__5293\,
            I => \N__5287\
        );

    \I__1098\ : Span4Mux_s3_h
    port map (
            O => \N__5290\,
            I => \N__5284\
        );

    \I__1097\ : Span4Mux_s1_h
    port map (
            O => \N__5287\,
            I => \N__5281\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__5284\,
            I => \uart.n2310\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__5281\,
            I => \uart.n2310\
        );

    \I__1094\ : IoInMux
    port map (
            O => \N__5276\,
            I => \N__5272\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__5275\,
            I => \N__5269\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5272\,
            I => \N__5266\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5263\
        );

    \I__1090\ : IoSpan4Mux
    port map (
            O => \N__5266\,
            I => \N__5260\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5263\,
            I => \N__5257\
        );

    \I__1088\ : Span4Mux_s2_v
    port map (
            O => \N__5260\,
            I => \N__5254\
        );

    \I__1087\ : Span4Mux_h
    port map (
            O => \N__5257\,
            I => \N__5251\
        );

    \I__1086\ : Sp12to4
    port map (
            O => \N__5254\,
            I => \N__5248\
        );

    \I__1085\ : Sp12to4
    port map (
            O => \N__5251\,
            I => \N__5245\
        );

    \I__1084\ : Span12Mux_h
    port map (
            O => \N__5248\,
            I => \N__5242\
        );

    \I__1083\ : Span12Mux_v
    port map (
            O => \N__5245\,
            I => \N__5239\
        );

    \I__1082\ : Span12Mux_h
    port map (
            O => \N__5242\,
            I => \N__5234\
        );

    \I__1081\ : Span12Mux_v
    port map (
            O => \N__5239\,
            I => \N__5234\
        );

    \I__1080\ : Odrv12
    port map (
            O => \N__5234\,
            I => diff_input
        );

    \I__1079\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5227\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5224\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5227\,
            I => integrator_0
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5224\,
            I => integrator_0
        );

    \I__1075\ : InMux
    port map (
            O => \N__5219\,
            I => \N__5215\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5218\,
            I => \N__5212\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5215\,
            I => integrator_1
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5212\,
            I => integrator_1
        );

    \I__1071\ : InMux
    port map (
            O => \N__5207\,
            I => n2188
        );

    \I__1070\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5200\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5197\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5200\,
            I => \N__5194\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5197\,
            I => counter_13
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__5194\,
            I => counter_13
        );

    \I__1065\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5185\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5182\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5185\,
            I => counter_23
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5182\,
            I => counter_23
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__5177\,
            I => \N__5173\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5170\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5173\,
            I => \N__5167\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5170\,
            I => counter_11
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5167\,
            I => counter_11
        );

    \I__1056\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5158\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5155\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5158\,
            I => counter_14
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5155\,
            I => counter_14
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__5150\,
            I => \n38_cascade_\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__5147\,
            I => \n44_cascade_\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__5144\,
            I => \counter_31__N_172_cascade_\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5138\,
            I => \N__5134\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5131\
        );

    \I__1046\ : Odrv12
    port map (
            O => \N__5134\,
            I => data_out_4
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5131\,
            I => data_out_4
        );

    \I__1044\ : InMux
    port map (
            O => \N__5126\,
            I => \N__5120\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5120\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5120\,
            I => \N__5116\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5113\
        );

    \I__1040\ : Span4Mux_h
    port map (
            O => \N__5116\,
            I => \N__5110\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5113\,
            I => counter_31
        );

    \I__1038\ : Odrv4
    port map (
            O => \N__5110\,
            I => counter_31
        );

    \I__1037\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5102\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5102\,
            I => n44
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__5099\,
            I => \N__5096\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5093\,
            I => \N__5089\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__5092\,
            I => \N__5086\
        );

    \I__1031\ : Span4Mux_s3_h
    port map (
            O => \N__5089\,
            I => \N__5083\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5080\
        );

    \I__1029\ : Sp12to4
    port map (
            O => \N__5083\,
            I => \N__5075\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__5080\,
            I => \N__5075\
        );

    \I__1027\ : Odrv12
    port map (
            O => \N__5075\,
            I => \r_SM_Main_2_N_236_0\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5069\,
            I => \N__5065\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5062\
        );

    \I__1023\ : Odrv12
    port map (
            O => \N__5065\,
            I => data_out_6
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__5062\,
            I => data_out_6
        );

    \I__1021\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5053\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5050\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5053\,
            I => counter_22
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5050\,
            I => counter_22
        );

    \I__1017\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5041\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5038\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5041\,
            I => counter_30
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5038\,
            I => counter_30
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__5033\,
            I => \N__5029\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5026\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5023\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5026\,
            I => counter_19
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5023\,
            I => counter_19
        );

    \I__1008\ : InMux
    port map (
            O => \N__5018\,
            I => \N__5014\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5011\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5014\,
            I => counter_26
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__5011\,
            I => counter_26
        );

    \I__1004\ : InMux
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5003\,
            I => n36
        );

    \I__1002\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4996\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4993\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4996\,
            I => counter_12
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4993\,
            I => counter_12
        );

    \I__998\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4984\
        );

    \I__997\ : InMux
    port map (
            O => \N__4987\,
            I => \N__4981\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4984\,
            I => counter_8
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4981\,
            I => counter_8
        );

    \I__994\ : CascadeMux
    port map (
            O => \N__4976\,
            I => \N__4972\
        );

    \I__993\ : InMux
    port map (
            O => \N__4975\,
            I => \N__4969\
        );

    \I__992\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4966\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4969\,
            I => counter_15
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4966\,
            I => counter_15
        );

    \I__989\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4957\
        );

    \I__988\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4954\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4957\,
            I => counter_25
        );

    \I__986\ : LocalMux
    port map (
            O => \N__4954\,
            I => counter_25
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__984\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4942\
        );

    \I__983\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4939\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4942\,
            I => \N__4934\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4939\,
            I => \N__4934\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__4934\,
            I => n40
        );

    \I__979\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4927\
        );

    \I__978\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4924\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4927\,
            I => \r_Tx_Data_3\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4924\,
            I => \r_Tx_Data_3\
        );

    \I__975\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4915\
        );

    \I__974\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4912\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4915\,
            I => \r_Tx_Data_7\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4912\,
            I => \r_Tx_Data_7\
        );

    \I__971\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4903\
        );

    \I__970\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4900\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4903\,
            I => \r_Tx_Data_0\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4900\,
            I => \r_Tx_Data_0\
        );

    \I__967\ : InMux
    port map (
            O => \N__4895\,
            I => \N__4877\
        );

    \I__966\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4877\
        );

    \I__965\ : InMux
    port map (
            O => \N__4893\,
            I => \N__4877\
        );

    \I__964\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4877\
        );

    \I__963\ : InMux
    port map (
            O => \N__4891\,
            I => \N__4877\
        );

    \I__962\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4870\
        );

    \I__961\ : InMux
    port map (
            O => \N__4889\,
            I => \N__4870\
        );

    \I__960\ : InMux
    port map (
            O => \N__4888\,
            I => \N__4870\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4877\,
            I => n1757
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4870\,
            I => n1757
        );

    \I__957\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4861\
        );

    \I__956\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4858\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4861\,
            I => \r_Tx_Data_2\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4858\,
            I => \r_Tx_Data_2\
        );

    \I__953\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4850\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4850\,
            I => \N__4846\
        );

    \I__951\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4843\
        );

    \I__950\ : Odrv12
    port map (
            O => \N__4846\,
            I => data_out_5
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4843\,
            I => data_out_5
        );

    \I__948\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4835\,
            I => \N__4831\
        );

    \I__946\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4828\
        );

    \I__945\ : Odrv4
    port map (
            O => \N__4831\,
            I => data_out_0
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4828\,
            I => data_out_0
        );

    \I__943\ : InMux
    port map (
            O => \N__4823\,
            I => \N__4819\
        );

    \I__942\ : InMux
    port map (
            O => \N__4822\,
            I => \N__4816\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4819\,
            I => data_out_3
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4816\,
            I => data_out_3
        );

    \I__939\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4808\,
            I => \N__4804\
        );

    \I__937\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4801\
        );

    \I__936\ : Odrv4
    port map (
            O => \N__4804\,
            I => data_out_1
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4801\,
            I => data_out_1
        );

    \I__934\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4793\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4793\,
            I => \N__4789\
        );

    \I__932\ : InMux
    port map (
            O => \N__4792\,
            I => \N__4786\
        );

    \I__931\ : Odrv12
    port map (
            O => \N__4789\,
            I => data_out_2
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4786\,
            I => data_out_2
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__4781\,
            I => \uart.n2428_cascade_\
        );

    \I__928\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4775\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4775\,
            I => \uart.n2431\
        );

    \I__926\ : InMux
    port map (
            O => \N__4772\,
            I => \N__4766\
        );

    \I__925\ : InMux
    port map (
            O => \N__4771\,
            I => \N__4766\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4766\,
            I => \r_Tx_Data_4\
        );

    \I__923\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4757\
        );

    \I__922\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4757\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4757\,
            I => \r_Tx_Data_5\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__4754\,
            I => \uart.n2422_cascade_\
        );

    \I__919\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4748\,
            I => \uart.n2425\
        );

    \I__917\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4739\
        );

    \I__916\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4739\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4739\,
            I => \r_Tx_Data_6\
        );

    \I__914\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4733\,
            I => \N__4726\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__4732\,
            I => \N__4722\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__4731\,
            I => \N__4716\
        );

    \I__910\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4713\
        );

    \I__909\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4710\
        );

    \I__908\ : Span4Mux_v
    port map (
            O => \N__4726\,
            I => \N__4707\
        );

    \I__907\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4704\
        );

    \I__906\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4697\
        );

    \I__905\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4697\
        );

    \I__904\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4697\
        );

    \I__903\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4692\
        );

    \I__902\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4692\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4713\,
            I => \r_SM_Main_1\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4710\,
            I => \r_SM_Main_1\
        );

    \I__899\ : Odrv4
    port map (
            O => \N__4707\,
            I => \r_SM_Main_1\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4704\,
            I => \r_SM_Main_1\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4697\,
            I => \r_SM_Main_1\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4692\,
            I => \r_SM_Main_1\
        );

    \I__895\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4674\
        );

    \I__894\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4667\
        );

    \I__893\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4667\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4674\,
            I => \N__4664\
        );

    \I__891\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4657\
        );

    \I__890\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4657\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4667\,
            I => \N__4652\
        );

    \I__888\ : Span4Mux_v
    port map (
            O => \N__4664\,
            I => \N__4652\
        );

    \I__887\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4649\
        );

    \I__886\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4646\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4657\,
            I => \r_SM_Main_0\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__4652\,
            I => \r_SM_Main_0\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4649\,
            I => \r_SM_Main_0\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4646\,
            I => \r_SM_Main_0\
        );

    \I__881\ : InMux
    port map (
            O => \N__4637\,
            I => \N__4633\
        );

    \I__880\ : SRMux
    port map (
            O => \N__4636\,
            I => \N__4626\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4633\,
            I => \N__4623\
        );

    \I__878\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4620\
        );

    \I__877\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4617\
        );

    \I__876\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4612\
        );

    \I__875\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4612\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4626\,
            I => \N__4605\
        );

    \I__873\ : Span4Mux_v
    port map (
            O => \N__4623\,
            I => \N__4605\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4620\,
            I => \N__4605\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4617\,
            I => \r_SM_Main_2\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4612\,
            I => \r_SM_Main_2\
        );

    \I__869\ : Odrv4
    port map (
            O => \N__4605\,
            I => \r_SM_Main_2\
        );

    \I__868\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4594\
        );

    \I__867\ : InMux
    port map (
            O => \N__4597\,
            I => \N__4591\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4594\,
            I => \r_Tx_Data_1\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4591\,
            I => \r_Tx_Data_1\
        );

    \I__864\ : InMux
    port map (
            O => \N__4586\,
            I => n2221
        );

    \I__863\ : InMux
    port map (
            O => \N__4583\,
            I => n2222
        );

    \I__862\ : InMux
    port map (
            O => \N__4580\,
            I => n2223
        );

    \I__861\ : InMux
    port map (
            O => \N__4577\,
            I => n2224
        );

    \I__860\ : InMux
    port map (
            O => \N__4574\,
            I => n2225
        );

    \I__859\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4566\
        );

    \I__858\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4563\
        );

    \I__857\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4560\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4566\,
            I => \uart.r_Bit_Index_2\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4563\,
            I => \uart.r_Bit_Index_2\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4560\,
            I => \uart.r_Bit_Index_2\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__4553\,
            I => \n2002_cascade_\
        );

    \I__852\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4543\
        );

    \I__851\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4538\
        );

    \I__850\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4538\
        );

    \I__849\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4533\
        );

    \I__848\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4533\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4543\,
            I => \N__4530\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4538\,
            I => \r_SM_Main_2_N_233_1\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4533\,
            I => \r_SM_Main_2_N_233_1\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__4530\,
            I => \r_SM_Main_2_N_233_1\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__4523\,
            I => \n2308_cascade_\
        );

    \I__842\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4516\
        );

    \I__841\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4513\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4516\,
            I => \N__4510\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4513\,
            I => n2002
        );

    \I__838\ : Odrv4
    port map (
            O => \N__4510\,
            I => n2002
        );

    \I__837\ : InMux
    port map (
            O => \N__4505\,
            I => n2211
        );

    \I__836\ : InMux
    port map (
            O => \N__4502\,
            I => n2212
        );

    \I__835\ : InMux
    port map (
            O => \N__4499\,
            I => n2213
        );

    \I__834\ : InMux
    port map (
            O => \N__4496\,
            I => n2214
        );

    \I__833\ : InMux
    port map (
            O => \N__4493\,
            I => n2215
        );

    \I__832\ : InMux
    port map (
            O => \N__4490\,
            I => n2216
        );

    \I__831\ : InMux
    port map (
            O => \N__4487\,
            I => n2217
        );

    \I__830\ : InMux
    port map (
            O => \N__4484\,
            I => \bfn_3_25_0_\
        );

    \I__829\ : InMux
    port map (
            O => \N__4481\,
            I => n2219
        );

    \I__828\ : InMux
    port map (
            O => \N__4478\,
            I => n2220
        );

    \I__827\ : InMux
    port map (
            O => \N__4475\,
            I => \bfn_3_23_0_\
        );

    \I__826\ : InMux
    port map (
            O => \N__4472\,
            I => n2203
        );

    \I__825\ : InMux
    port map (
            O => \N__4469\,
            I => n2204
        );

    \I__824\ : InMux
    port map (
            O => \N__4466\,
            I => n2205
        );

    \I__823\ : InMux
    port map (
            O => \N__4463\,
            I => n2206
        );

    \I__822\ : InMux
    port map (
            O => \N__4460\,
            I => n2207
        );

    \I__821\ : InMux
    port map (
            O => \N__4457\,
            I => n2208
        );

    \I__820\ : InMux
    port map (
            O => \N__4454\,
            I => n2209
        );

    \I__819\ : InMux
    port map (
            O => \N__4451\,
            I => \bfn_3_24_0_\
        );

    \I__818\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4445\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4445\,
            I => counter_0
        );

    \I__816\ : InMux
    port map (
            O => \N__4442\,
            I => \bfn_3_22_0_\
        );

    \I__815\ : InMux
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4436\,
            I => counter_1
        );

    \I__813\ : InMux
    port map (
            O => \N__4433\,
            I => n2195
        );

    \I__812\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4427\,
            I => counter_2
        );

    \I__810\ : InMux
    port map (
            O => \N__4424\,
            I => n2196
        );

    \I__809\ : InMux
    port map (
            O => \N__4421\,
            I => \N__4418\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4418\,
            I => counter_3
        );

    \I__807\ : InMux
    port map (
            O => \N__4415\,
            I => n2197
        );

    \I__806\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4409\,
            I => counter_4
        );

    \I__804\ : InMux
    port map (
            O => \N__4406\,
            I => n2198
        );

    \I__803\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__4400\,
            I => counter_5
        );

    \I__801\ : InMux
    port map (
            O => \N__4397\,
            I => n2199
        );

    \I__800\ : InMux
    port map (
            O => \N__4394\,
            I => \N__4391\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4391\,
            I => counter_6
        );

    \I__798\ : InMux
    port map (
            O => \N__4388\,
            I => n2200
        );

    \I__797\ : InMux
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4382\,
            I => counter_7
        );

    \I__795\ : InMux
    port map (
            O => \N__4379\,
            I => n2201
        );

    \I__794\ : InMux
    port map (
            O => \N__4376\,
            I => n2187
        );

    \I__793\ : InMux
    port map (
            O => \N__4373\,
            I => \N__4369\
        );

    \I__792\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4366\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4369\,
            I => blink_counter_25
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4366\,
            I => blink_counter_25
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__4361\,
            I => \n2395_cascade_\
        );

    \I__788\ : IoInMux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__786\ : Span4Mux_s1_v
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__785\ : Span4Mux_v
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__4346\,
            I => \LED_c\
        );

    \I__783\ : InMux
    port map (
            O => \N__4343\,
            I => \N__4337\
        );

    \I__782\ : InMux
    port map (
            O => \N__4342\,
            I => \N__4337\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4337\,
            I => \N__4333\
        );

    \I__780\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4330\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__4333\,
            I => blink_counter_21
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4330\,
            I => blink_counter_21
        );

    \I__777\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4318\
        );

    \I__776\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4318\
        );

    \I__775\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4315\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4318\,
            I => blink_counter_24
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4315\,
            I => blink_counter_24
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__4310\,
            I => \N__4306\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__4309\,
            I => \N__4303\
        );

    \I__770\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4298\
        );

    \I__769\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4298\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4298\,
            I => \N__4294\
        );

    \I__767\ : InMux
    port map (
            O => \N__4297\,
            I => \N__4291\
        );

    \I__766\ : Odrv4
    port map (
            O => \N__4294\,
            I => blink_counter_23
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4291\,
            I => blink_counter_23
        );

    \I__764\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4280\
        );

    \I__763\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4280\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4280\,
            I => \N__4276\
        );

    \I__761\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4273\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__4276\,
            I => blink_counter_22
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4273\,
            I => blink_counter_22
        );

    \I__758\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4265\,
            I => n2394
        );

    \I__756\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4259\,
            I => \uart.n1711\
        );

    \I__754\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4253\,
            I => \uart.o_Tx_Serial_N_312\
        );

    \I__752\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4247\,
            I => \N__4243\
        );

    \I__750\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4240\
        );

    \I__749\ : Span4Mux_h
    port map (
            O => \N__4243\,
            I => \N__4237\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4240\,
            I => clk_divider_7
        );

    \I__747\ : Odrv4
    port map (
            O => \N__4237\,
            I => clk_divider_7
        );

    \I__746\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4229\,
            I => n40_adj_362
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__4226\,
            I => \N__4223\
        );

    \I__743\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4220\,
            I => \N__4216\
        );

    \I__741\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4213\
        );

    \I__740\ : Span4Mux_h
    port map (
            O => \N__4216\,
            I => \N__4210\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4213\,
            I => clk_divider_25
        );

    \I__738\ : Odrv4
    port map (
            O => \N__4210\,
            I => clk_divider_25
        );

    \I__737\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4202\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4202\,
            I => n45_adj_357
        );

    \I__735\ : InMux
    port map (
            O => \N__4199\,
            I => \N__4193\
        );

    \I__734\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4193\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4193\,
            I => n49
        );

    \I__732\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4187\,
            I => n9
        );

    \I__730\ : InMux
    port map (
            O => \N__4184\,
            I => n2179
        );

    \I__729\ : InMux
    port map (
            O => \N__4181\,
            I => \N__4178\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4178\,
            I => n8
        );

    \I__727\ : InMux
    port map (
            O => \N__4175\,
            I => n2180
        );

    \I__726\ : InMux
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4169\,
            I => n7
        );

    \I__724\ : InMux
    port map (
            O => \N__4166\,
            I => n2181
        );

    \I__723\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4160\,
            I => n6
        );

    \I__721\ : InMux
    port map (
            O => \N__4157\,
            I => n2182
        );

    \I__720\ : InMux
    port map (
            O => \N__4154\,
            I => n2183
        );

    \I__719\ : InMux
    port map (
            O => \N__4151\,
            I => n2184
        );

    \I__718\ : InMux
    port map (
            O => \N__4148\,
            I => n2185
        );

    \I__717\ : InMux
    port map (
            O => \N__4145\,
            I => \bfn_2_26_0_\
        );

    \I__716\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4139\,
            I => n18
        );

    \I__714\ : InMux
    port map (
            O => \N__4136\,
            I => \bfn_2_24_0_\
        );

    \I__713\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4130\,
            I => n17
        );

    \I__711\ : InMux
    port map (
            O => \N__4127\,
            I => n2171
        );

    \I__710\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4121\,
            I => n16
        );

    \I__708\ : InMux
    port map (
            O => \N__4118\,
            I => n2172
        );

    \I__707\ : InMux
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4112\,
            I => n15
        );

    \I__705\ : InMux
    port map (
            O => \N__4109\,
            I => n2173
        );

    \I__704\ : InMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4103\,
            I => n14
        );

    \I__702\ : InMux
    port map (
            O => \N__4100\,
            I => n2174
        );

    \I__701\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4094\,
            I => n13
        );

    \I__699\ : InMux
    port map (
            O => \N__4091\,
            I => n2175
        );

    \I__698\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4085\,
            I => n12
        );

    \I__696\ : InMux
    port map (
            O => \N__4082\,
            I => n2176
        );

    \I__695\ : InMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4076\,
            I => n11
        );

    \I__693\ : InMux
    port map (
            O => \N__4073\,
            I => n2177
        );

    \I__692\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__4067\,
            I => n10_adj_317
        );

    \I__690\ : InMux
    port map (
            O => \N__4064\,
            I => \bfn_2_25_0_\
        );

    \I__689\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__4058\,
            I => n26
        );

    \I__687\ : InMux
    port map (
            O => \N__4055\,
            I => \bfn_2_23_0_\
        );

    \I__686\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4049\,
            I => n25
        );

    \I__684\ : InMux
    port map (
            O => \N__4046\,
            I => n2163
        );

    \I__683\ : InMux
    port map (
            O => \N__4043\,
            I => \N__4040\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4040\,
            I => n24
        );

    \I__681\ : InMux
    port map (
            O => \N__4037\,
            I => n2164
        );

    \I__680\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4031\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4031\,
            I => n23
        );

    \I__678\ : InMux
    port map (
            O => \N__4028\,
            I => n2165
        );

    \I__677\ : InMux
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4022\,
            I => n22
        );

    \I__675\ : InMux
    port map (
            O => \N__4019\,
            I => n2166
        );

    \I__674\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4013\,
            I => n21
        );

    \I__672\ : InMux
    port map (
            O => \N__4010\,
            I => n2167
        );

    \I__671\ : InMux
    port map (
            O => \N__4007\,
            I => \N__4004\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4004\,
            I => n20
        );

    \I__669\ : InMux
    port map (
            O => \N__4001\,
            I => n2168
        );

    \I__668\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3995\,
            I => n19
        );

    \I__666\ : InMux
    port map (
            O => \N__3992\,
            I => n2169
        );

    \I__665\ : InMux
    port map (
            O => \N__3989\,
            I => \N__3985\
        );

    \I__664\ : InMux
    port map (
            O => \N__3988\,
            I => \N__3982\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3985\,
            I => \N__3979\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3982\,
            I => clk_divider_4
        );

    \I__661\ : Odrv4
    port map (
            O => \N__3979\,
            I => clk_divider_4
        );

    \I__660\ : InMux
    port map (
            O => \N__3974\,
            I => \N__3970\
        );

    \I__659\ : InMux
    port map (
            O => \N__3973\,
            I => \N__3967\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3970\,
            I => clk_divider_0
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3967\,
            I => clk_divider_0
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__3962\,
            I => \N__3958\
        );

    \I__655\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3955\
        );

    \I__654\ : InMux
    port map (
            O => \N__3958\,
            I => \N__3952\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3955\,
            I => clk_divider_3
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3952\,
            I => clk_divider_3
        );

    \I__651\ : SRMux
    port map (
            O => \N__3947\,
            I => \N__3943\
        );

    \I__650\ : SRMux
    port map (
            O => \N__3946\,
            I => \N__3939\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3943\,
            I => \N__3935\
        );

    \I__648\ : SRMux
    port map (
            O => \N__3942\,
            I => \N__3932\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3939\,
            I => \N__3929\
        );

    \I__646\ : SRMux
    port map (
            O => \N__3938\,
            I => \N__3926\
        );

    \I__645\ : Span4Mux_v
    port map (
            O => \N__3935\,
            I => \N__3921\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3932\,
            I => \N__3921\
        );

    \I__643\ : Span4Mux_v
    port map (
            O => \N__3929\,
            I => \N__3916\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3926\,
            I => \N__3916\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__3921\,
            I => \clk_divider_31__N_139\
        );

    \I__640\ : Odrv4
    port map (
            O => \N__3916\,
            I => \clk_divider_31__N_139\
        );

    \I__639\ : IoInMux
    port map (
            O => \N__3911\,
            I => \N__3908\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3908\,
            I => \N__3905\
        );

    \I__637\ : Span12Mux_s1_v
    port map (
            O => \N__3905\,
            I => \N__3902\
        );

    \I__636\ : Odrv12
    port map (
            O => \N__3902\,
            I => \uart.n3\
        );

    \I__635\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3895\
        );

    \I__634\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3892\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3895\,
            I => clk_divider_1
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3892\,
            I => clk_divider_1
        );

    \I__631\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3883\
        );

    \I__630\ : InMux
    port map (
            O => \N__3886\,
            I => \N__3880\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3883\,
            I => clk_divider_2
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3880\,
            I => clk_divider_2
        );

    \I__627\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3872\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3872\,
            I => n6_adj_324
        );

    \I__625\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3865\
        );

    \I__624\ : InMux
    port map (
            O => \N__3868\,
            I => \N__3862\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3865\,
            I => clk_divider_8
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3862\,
            I => clk_divider_8
        );

    \I__621\ : InMux
    port map (
            O => \N__3857\,
            I => \N__3853\
        );

    \I__620\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3850\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3853\,
            I => clk_divider_15
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3850\,
            I => clk_divider_15
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__3845\,
            I => \N__3842\
        );

    \I__616\ : InMux
    port map (
            O => \N__3842\,
            I => \N__3838\
        );

    \I__615\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3835\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3838\,
            I => \N__3832\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3835\,
            I => clk_divider_24
        );

    \I__612\ : Odrv4
    port map (
            O => \N__3832\,
            I => clk_divider_24
        );

    \I__611\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3823\
        );

    \I__610\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3820\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3823\,
            I => clk_divider_11
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3820\,
            I => clk_divider_11
        );

    \I__607\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3811\
        );

    \I__606\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3808\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3811\,
            I => clk_divider_5
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3808\,
            I => clk_divider_5
        );

    \I__603\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3799\
        );

    \I__602\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3796\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3799\,
            I => clk_divider_10
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3796\,
            I => clk_divider_10
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__3791\,
            I => \N__3787\
        );

    \I__598\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3784\
        );

    \I__597\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3781\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3784\,
            I => clk_divider_12
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3781\,
            I => clk_divider_12
        );

    \I__594\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3772\
        );

    \I__593\ : InMux
    port map (
            O => \N__3775\,
            I => \N__3769\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3772\,
            I => \N__3766\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3769\,
            I => clk_divider_18
        );

    \I__590\ : Odrv4
    port map (
            O => \N__3766\,
            I => clk_divider_18
        );

    \I__589\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3757\
        );

    \I__588\ : InMux
    port map (
            O => \N__3760\,
            I => \N__3754\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3757\,
            I => clk_divider_13
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3754\,
            I => clk_divider_13
        );

    \I__585\ : InMux
    port map (
            O => \N__3749\,
            I => \N__3745\
        );

    \I__584\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3742\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3745\,
            I => \N__3739\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3742\,
            I => clk_divider_29
        );

    \I__581\ : Odrv4
    port map (
            O => \N__3739\,
            I => clk_divider_29
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__579\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3728\,
            I => \N__3724\
        );

    \I__577\ : InMux
    port map (
            O => \N__3727\,
            I => \N__3721\
        );

    \I__576\ : Span4Mux_h
    port map (
            O => \N__3724\,
            I => \N__3718\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3721\,
            I => clk_divider_23
        );

    \I__574\ : Odrv4
    port map (
            O => \N__3718\,
            I => clk_divider_23
        );

    \I__573\ : InMux
    port map (
            O => \N__3713\,
            I => \N__3709\
        );

    \I__572\ : InMux
    port map (
            O => \N__3712\,
            I => \N__3706\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3709\,
            I => \N__3703\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3706\,
            I => clk_divider_16
        );

    \I__569\ : Odrv4
    port map (
            O => \N__3703\,
            I => clk_divider_16
        );

    \I__568\ : InMux
    port map (
            O => \N__3698\,
            I => \N__3695\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3695\,
            I => n43_adj_359
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__3692\,
            I => \N__3688\
        );

    \I__565\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3683\
        );

    \I__564\ : InMux
    port map (
            O => \N__3688\,
            I => \N__3683\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3683\,
            I => \N__3679\
        );

    \I__562\ : InMux
    port map (
            O => \N__3682\,
            I => \N__3676\
        );

    \I__561\ : Span4Mux_h
    port map (
            O => \N__3679\,
            I => \N__3673\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3676\,
            I => clk_divider_31
        );

    \I__559\ : Odrv4
    port map (
            O => \N__3673\,
            I => clk_divider_31
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__557\ : InMux
    port map (
            O => \N__3665\,
            I => \N__3659\
        );

    \I__556\ : InMux
    port map (
            O => \N__3664\,
            I => \N__3659\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3659\,
            I => n50
        );

    \I__554\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3650\
        );

    \I__553\ : InMux
    port map (
            O => \N__3655\,
            I => \N__3650\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3650\,
            I => \N__3647\
        );

    \I__551\ : Odrv4
    port map (
            O => \N__3647\,
            I => n10
        );

    \I__550\ : InMux
    port map (
            O => \N__3644\,
            I => \N__3640\
        );

    \I__549\ : InMux
    port map (
            O => \N__3643\,
            I => \N__3637\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3640\,
            I => \uart.r_Clock_Count_20\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3637\,
            I => \uart.r_Clock_Count_20\
        );

    \I__546\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3628\
        );

    \I__545\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3625\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3628\,
            I => \uart.r_Clock_Count_15\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3625\,
            I => \uart.r_Clock_Count_15\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__3620\,
            I => \N__3616\
        );

    \I__541\ : InMux
    port map (
            O => \N__3619\,
            I => \N__3613\
        );

    \I__540\ : InMux
    port map (
            O => \N__3616\,
            I => \N__3610\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3613\,
            I => \uart.r_Clock_Count_25\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3610\,
            I => \uart.r_Clock_Count_25\
        );

    \I__537\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3601\
        );

    \I__536\ : InMux
    port map (
            O => \N__3604\,
            I => \N__3598\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3601\,
            I => \uart.r_Clock_Count_9\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3598\,
            I => \uart.r_Clock_Count_9\
        );

    \I__533\ : InMux
    port map (
            O => \N__3593\,
            I => \N__3589\
        );

    \I__532\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3586\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3589\,
            I => \N__3583\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3586\,
            I => \uart.r_Clock_Count_27\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__3583\,
            I => \uart.r_Clock_Count_27\
        );

    \I__528\ : InMux
    port map (
            O => \N__3578\,
            I => \N__3574\
        );

    \I__527\ : InMux
    port map (
            O => \N__3577\,
            I => \N__3571\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3574\,
            I => \uart.r_Clock_Count_19\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3571\,
            I => \uart.r_Clock_Count_19\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__3566\,
            I => \N__3562\
        );

    \I__523\ : InMux
    port map (
            O => \N__3565\,
            I => \N__3559\
        );

    \I__522\ : InMux
    port map (
            O => \N__3562\,
            I => \N__3556\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3559\,
            I => \uart.r_Clock_Count_16\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3556\,
            I => \uart.r_Clock_Count_16\
        );

    \I__519\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3547\
        );

    \I__518\ : InMux
    port map (
            O => \N__3550\,
            I => \N__3544\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3547\,
            I => \uart.r_Clock_Count_31\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3544\,
            I => \uart.r_Clock_Count_31\
        );

    \I__515\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3536\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3536\,
            I => \uart.n39\
        );

    \I__513\ : InMux
    port map (
            O => \N__3533\,
            I => \N__3530\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3530\,
            I => \uart.n40\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3527\,
            I => \uart.n37_cascade_\
        );

    \I__510\ : InMux
    port map (
            O => \N__3524\,
            I => \N__3521\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3521\,
            I => \uart.n38\
        );

    \I__508\ : InMux
    port map (
            O => \N__3518\,
            I => \N__3515\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3515\,
            I => \N__3512\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__3512\,
            I => \uart.n46\
        );

    \I__505\ : InMux
    port map (
            O => \N__3509\,
            I => \N__3506\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3506\,
            I => \N__3502\
        );

    \I__503\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3499\
        );

    \I__502\ : Span4Mux_h
    port map (
            O => \N__3502\,
            I => \N__3496\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3499\,
            I => clk_divider_26
        );

    \I__500\ : Odrv4
    port map (
            O => \N__3496\,
            I => clk_divider_26
        );

    \I__499\ : InMux
    port map (
            O => \N__3491\,
            I => \N__3487\
        );

    \I__498\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3484\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3487\,
            I => \N__3481\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3484\,
            I => clk_divider_9
        );

    \I__495\ : Odrv4
    port map (
            O => \N__3481\,
            I => clk_divider_9
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__3476\,
            I => \N__3473\
        );

    \I__493\ : InMux
    port map (
            O => \N__3473\,
            I => \N__3469\
        );

    \I__492\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3466\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3469\,
            I => \N__3463\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3466\,
            I => clk_divider_14
        );

    \I__489\ : Odrv4
    port map (
            O => \N__3463\,
            I => clk_divider_14
        );

    \I__488\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3455\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3451\
        );

    \I__486\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3448\
        );

    \I__485\ : Span4Mux_h
    port map (
            O => \N__3451\,
            I => \N__3445\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3448\,
            I => clk_divider_17
        );

    \I__483\ : Odrv4
    port map (
            O => \N__3445\,
            I => clk_divider_17
        );

    \I__482\ : InMux
    port map (
            O => \N__3440\,
            I => \N__3436\
        );

    \I__481\ : InMux
    port map (
            O => \N__3439\,
            I => \N__3433\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3436\,
            I => \N__3430\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3433\,
            I => clk_divider_21
        );

    \I__478\ : Odrv4
    port map (
            O => \N__3430\,
            I => clk_divider_21
        );

    \I__477\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3422\,
            I => \N__3418\
        );

    \I__475\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3415\
        );

    \I__474\ : Span4Mux_h
    port map (
            O => \N__3418\,
            I => \N__3412\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3415\,
            I => clk_divider_22
        );

    \I__472\ : Odrv4
    port map (
            O => \N__3412\,
            I => clk_divider_22
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__3407\,
            I => \N__3404\
        );

    \I__470\ : InMux
    port map (
            O => \N__3404\,
            I => \N__3401\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3401\,
            I => \N__3397\
        );

    \I__468\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3394\
        );

    \I__467\ : Span4Mux_h
    port map (
            O => \N__3397\,
            I => \N__3391\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3394\,
            I => clk_divider_28
        );

    \I__465\ : Odrv4
    port map (
            O => \N__3391\,
            I => clk_divider_28
        );

    \I__464\ : InMux
    port map (
            O => \N__3386\,
            I => \N__3382\
        );

    \I__463\ : InMux
    port map (
            O => \N__3385\,
            I => \N__3379\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3382\,
            I => clk_divider_6
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3379\,
            I => clk_divider_6
        );

    \I__460\ : InMux
    port map (
            O => \N__3374\,
            I => \N__3371\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3371\,
            I => \N__3367\
        );

    \I__458\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3364\
        );

    \I__457\ : Span4Mux_v
    port map (
            O => \N__3367\,
            I => \N__3361\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3364\,
            I => clk_divider_30
        );

    \I__455\ : Odrv4
    port map (
            O => \N__3361\,
            I => clk_divider_30
        );

    \I__454\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3353\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3353\,
            I => \N__3349\
        );

    \I__452\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3346\
        );

    \I__451\ : Span4Mux_h
    port map (
            O => \N__3349\,
            I => \N__3343\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3346\,
            I => clk_divider_27
        );

    \I__449\ : Odrv4
    port map (
            O => \N__3343\,
            I => clk_divider_27
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__3338\,
            I => \N__3335\
        );

    \I__447\ : InMux
    port map (
            O => \N__3335\,
            I => \N__3331\
        );

    \I__446\ : InMux
    port map (
            O => \N__3334\,
            I => \N__3328\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3331\,
            I => \N__3325\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3328\,
            I => clk_divider_20
        );

    \I__443\ : Odrv4
    port map (
            O => \N__3325\,
            I => clk_divider_20
        );

    \I__442\ : InMux
    port map (
            O => \N__3320\,
            I => \N__3316\
        );

    \I__441\ : InMux
    port map (
            O => \N__3319\,
            I => \N__3313\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3316\,
            I => \N__3310\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3313\,
            I => clk_divider_19
        );

    \I__438\ : Odrv4
    port map (
            O => \N__3310\,
            I => clk_divider_19
        );

    \I__437\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3302\,
            I => n44_adj_358
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__3299\,
            I => \n42_adj_360_cascade_\
        );

    \I__434\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3293\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3293\,
            I => n41_adj_361
        );

    \I__432\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3286\
        );

    \I__431\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3283\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3286\,
            I => \uart.r_Clock_Count_13\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3283\,
            I => \uart.r_Clock_Count_13\
        );

    \I__428\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3274\
        );

    \I__427\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3271\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3274\,
            I => \uart.r_Clock_Count_12\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3271\,
            I => \uart.r_Clock_Count_12\
        );

    \I__424\ : InMux
    port map (
            O => \N__3266\,
            I => \N__3262\
        );

    \I__423\ : InMux
    port map (
            O => \N__3265\,
            I => \N__3259\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3262\,
            I => \N__3256\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3259\,
            I => \uart.r_Clock_Count_29\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__3256\,
            I => \uart.r_Clock_Count_29\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__3251\,
            I => \uart.n42_cascade_\
        );

    \I__418\ : InMux
    port map (
            O => \N__3248\,
            I => \N__3244\
        );

    \I__417\ : InMux
    port map (
            O => \N__3247\,
            I => \N__3241\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3244\,
            I => \uart.r_Clock_Count_7\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3241\,
            I => \uart.r_Clock_Count_7\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__3236\,
            I => \uart.n45_cascade_\
        );

    \I__413\ : InMux
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__3230\,
            I => \uart.n2385\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__3227\,
            I => \r_SM_Main_2_N_233_1_cascade_\
        );

    \I__410\ : SRMux
    port map (
            O => \N__3224\,
            I => \N__3221\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3221\,
            I => \N__3218\
        );

    \I__408\ : Span4Mux_s1_h
    port map (
            O => \N__3218\,
            I => \N__3212\
        );

    \I__407\ : SRMux
    port map (
            O => \N__3217\,
            I => \N__3209\
        );

    \I__406\ : SRMux
    port map (
            O => \N__3216\,
            I => \N__3206\
        );

    \I__405\ : SRMux
    port map (
            O => \N__3215\,
            I => \N__3203\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__3212\,
            I => \uart.n1796\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3209\,
            I => \uart.n1796\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3206\,
            I => \uart.n1796\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3203\,
            I => \uart.n1796\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__3194\,
            I => \N__3190\
        );

    \I__399\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3187\
        );

    \I__398\ : InMux
    port map (
            O => \N__3190\,
            I => \N__3184\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3187\,
            I => \uart.r_Clock_Count_8\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3184\,
            I => \uart.r_Clock_Count_8\
        );

    \I__395\ : InMux
    port map (
            O => \N__3179\,
            I => \N__3175\
        );

    \I__394\ : InMux
    port map (
            O => \N__3178\,
            I => \N__3172\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3175\,
            I => \uart.r_Clock_Count_14\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3172\,
            I => \uart.r_Clock_Count_14\
        );

    \I__391\ : InMux
    port map (
            O => \N__3167\,
            I => \N__3164\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3164\,
            I => \uart.n34\
        );

    \I__389\ : InMux
    port map (
            O => \N__3161\,
            I => \N__3157\
        );

    \I__388\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3154\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3157\,
            I => \uart.r_Clock_Count_30\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3154\,
            I => \uart.r_Clock_Count_30\
        );

    \I__385\ : InMux
    port map (
            O => \N__3149\,
            I => \N__3145\
        );

    \I__384\ : InMux
    port map (
            O => \N__3148\,
            I => \N__3142\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3145\,
            I => \uart.r_Clock_Count_28\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3142\,
            I => \uart.r_Clock_Count_28\
        );

    \I__381\ : CascadeMux
    port map (
            O => \N__3137\,
            I => \N__3134\
        );

    \I__380\ : InMux
    port map (
            O => \N__3134\,
            I => \N__3130\
        );

    \I__379\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3127\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3130\,
            I => \N__3124\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3127\,
            I => \uart.r_Clock_Count_24\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__3124\,
            I => \uart.r_Clock_Count_24\
        );

    \I__375\ : InMux
    port map (
            O => \N__3119\,
            I => \N__3115\
        );

    \I__374\ : InMux
    port map (
            O => \N__3118\,
            I => \N__3112\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3115\,
            I => \uart.r_Clock_Count_23\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3112\,
            I => \uart.r_Clock_Count_23\
        );

    \I__371\ : CEMux
    port map (
            O => \N__3107\,
            I => \N__3103\
        );

    \I__370\ : CEMux
    port map (
            O => \N__3106\,
            I => \N__3100\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3103\,
            I => \N__3097\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3100\,
            I => \N__3091\
        );

    \I__367\ : Span4Mux_s2_v
    port map (
            O => \N__3097\,
            I => \N__3088\
        );

    \I__366\ : CEMux
    port map (
            O => \N__3096\,
            I => \N__3085\
        );

    \I__365\ : CEMux
    port map (
            O => \N__3095\,
            I => \N__3082\
        );

    \I__364\ : CEMux
    port map (
            O => \N__3094\,
            I => \N__3079\
        );

    \I__363\ : Sp12to4
    port map (
            O => \N__3091\,
            I => \N__3074\
        );

    \I__362\ : Sp12to4
    port map (
            O => \N__3088\,
            I => \N__3074\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3085\,
            I => \uart.n1\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3082\,
            I => \uart.n1\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__3079\,
            I => \uart.n1\
        );

    \I__358\ : Odrv12
    port map (
            O => \N__3074\,
            I => \uart.n1\
        );

    \I__357\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3061\
        );

    \I__356\ : InMux
    port map (
            O => \N__3064\,
            I => \N__3058\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3061\,
            I => \uart.r_Clock_Count_11\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3058\,
            I => \uart.r_Clock_Count_11\
        );

    \I__353\ : InMux
    port map (
            O => \N__3053\,
            I => \N__3049\
        );

    \I__352\ : InMux
    port map (
            O => \N__3052\,
            I => \N__3046\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3049\,
            I => \uart.r_Clock_Count_21\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3046\,
            I => \uart.r_Clock_Count_21\
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__3041\,
            I => \N__3037\
        );

    \I__348\ : InMux
    port map (
            O => \N__3040\,
            I => \N__3034\
        );

    \I__347\ : InMux
    port map (
            O => \N__3037\,
            I => \N__3031\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3034\,
            I => \uart.r_Clock_Count_17\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__3031\,
            I => \uart.r_Clock_Count_17\
        );

    \I__344\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3022\
        );

    \I__343\ : InMux
    port map (
            O => \N__3025\,
            I => \N__3019\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3022\,
            I => \uart.r_Clock_Count_18\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3019\,
            I => \uart.r_Clock_Count_18\
        );

    \I__340\ : InMux
    port map (
            O => \N__3014\,
            I => n2252
        );

    \I__339\ : InMux
    port map (
            O => \N__3011\,
            I => n2253
        );

    \I__338\ : InMux
    port map (
            O => \N__3008\,
            I => n2254
        );

    \I__337\ : InMux
    port map (
            O => \N__3005\,
            I => n2255
        );

    \I__336\ : InMux
    port map (
            O => \N__3002\,
            I => n2256
        );

    \I__335\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2995\
        );

    \I__334\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2992\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2995\,
            I => \uart.r_Clock_Count_2\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2992\,
            I => \uart.r_Clock_Count_2\
        );

    \I__331\ : InMux
    port map (
            O => \N__2987\,
            I => \N__2983\
        );

    \I__330\ : InMux
    port map (
            O => \N__2986\,
            I => \N__2980\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2983\,
            I => \uart.r_Clock_Count_0\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2980\,
            I => \uart.r_Clock_Count_0\
        );

    \I__327\ : CascadeMux
    port map (
            O => \N__2975\,
            I => \N__2971\
        );

    \I__326\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2968\
        );

    \I__325\ : InMux
    port map (
            O => \N__2971\,
            I => \N__2965\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2968\,
            I => \uart.r_Clock_Count_1\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2965\,
            I => \uart.r_Clock_Count_1\
        );

    \I__322\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2956\
        );

    \I__321\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2953\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2956\,
            I => \uart.r_Clock_Count_3\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2953\,
            I => \uart.r_Clock_Count_3\
        );

    \I__318\ : InMux
    port map (
            O => \N__2948\,
            I => \N__2944\
        );

    \I__317\ : InMux
    port map (
            O => \N__2947\,
            I => \N__2941\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2944\,
            I => \uart.r_Clock_Count_5\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2941\,
            I => \uart.r_Clock_Count_5\
        );

    \I__314\ : InMux
    port map (
            O => \N__2936\,
            I => \N__2932\
        );

    \I__313\ : InMux
    port map (
            O => \N__2935\,
            I => \N__2929\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2932\,
            I => \uart.r_Clock_Count_4\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2929\,
            I => \uart.r_Clock_Count_4\
        );

    \I__310\ : CascadeMux
    port map (
            O => \N__2924\,
            I => \uart.n2006_cascade_\
        );

    \I__309\ : InMux
    port map (
            O => \N__2921\,
            I => \N__2917\
        );

    \I__308\ : InMux
    port map (
            O => \N__2920\,
            I => \N__2914\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2917\,
            I => \uart.r_Clock_Count_6\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2914\,
            I => \uart.r_Clock_Count_6\
        );

    \I__305\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2905\
        );

    \I__304\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2902\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2905\,
            I => \uart.r_Clock_Count_10\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2902\,
            I => \uart.r_Clock_Count_10\
        );

    \I__301\ : InMux
    port map (
            O => \N__2897\,
            I => \N__2893\
        );

    \I__300\ : InMux
    port map (
            O => \N__2896\,
            I => \N__2890\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2893\,
            I => \uart.r_Clock_Count_22\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2890\,
            I => \uart.r_Clock_Count_22\
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__296\ : InMux
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2879\,
            I => \N__2875\
        );

    \I__294\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2872\
        );

    \I__293\ : Span4Mux_v
    port map (
            O => \N__2875\,
            I => \N__2869\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2872\,
            I => \uart.r_Clock_Count_26\
        );

    \I__291\ : Odrv4
    port map (
            O => \N__2869\,
            I => \uart.r_Clock_Count_26\
        );

    \I__290\ : InMux
    port map (
            O => \N__2864\,
            I => n2243
        );

    \I__289\ : InMux
    port map (
            O => \N__2861\,
            I => n2244
        );

    \I__288\ : InMux
    port map (
            O => \N__2858\,
            I => n2245
        );

    \I__287\ : InMux
    port map (
            O => \N__2855\,
            I => n2246
        );

    \I__286\ : InMux
    port map (
            O => \N__2852\,
            I => n2247
        );

    \I__285\ : InMux
    port map (
            O => \N__2849\,
            I => n2248
        );

    \I__284\ : InMux
    port map (
            O => \N__2846\,
            I => \bfn_1_25_0_\
        );

    \I__283\ : InMux
    port map (
            O => \N__2843\,
            I => n2250
        );

    \I__282\ : InMux
    port map (
            O => \N__2840\,
            I => n2251
        );

    \I__281\ : InMux
    port map (
            O => \N__2837\,
            I => n2234
        );

    \I__280\ : InMux
    port map (
            O => \N__2834\,
            I => n2235
        );

    \I__279\ : InMux
    port map (
            O => \N__2831\,
            I => n2236
        );

    \I__278\ : InMux
    port map (
            O => \N__2828\,
            I => n2237
        );

    \I__277\ : InMux
    port map (
            O => \N__2825\,
            I => n2238
        );

    \I__276\ : InMux
    port map (
            O => \N__2822\,
            I => n2239
        );

    \I__275\ : InMux
    port map (
            O => \N__2819\,
            I => n2240
        );

    \I__274\ : InMux
    port map (
            O => \N__2816\,
            I => \bfn_1_24_0_\
        );

    \I__273\ : InMux
    port map (
            O => \N__2813\,
            I => n2242
        );

    \I__272\ : InMux
    port map (
            O => \N__2810\,
            I => \bfn_1_22_0_\
        );

    \I__271\ : InMux
    port map (
            O => \N__2807\,
            I => n2226
        );

    \I__270\ : InMux
    port map (
            O => \N__2804\,
            I => n2227
        );

    \I__269\ : InMux
    port map (
            O => \N__2801\,
            I => n2228
        );

    \I__268\ : InMux
    port map (
            O => \N__2798\,
            I => n2229
        );

    \I__267\ : InMux
    port map (
            O => \N__2795\,
            I => n2230
        );

    \I__266\ : InMux
    port map (
            O => \N__2792\,
            I => n2231
        );

    \I__265\ : InMux
    port map (
            O => \N__2789\,
            I => n2232
        );

    \I__264\ : InMux
    port map (
            O => \N__2786\,
            I => \bfn_1_23_0_\
        );

    \I__263\ : InMux
    port map (
            O => \N__2783\,
            I => \uart.n2154\
        );

    \I__262\ : InMux
    port map (
            O => \N__2780\,
            I => \bfn_1_21_0_\
        );

    \I__261\ : InMux
    port map (
            O => \N__2777\,
            I => \uart.n2156\
        );

    \I__260\ : InMux
    port map (
            O => \N__2774\,
            I => \uart.n2157\
        );

    \I__259\ : InMux
    port map (
            O => \N__2771\,
            I => \uart.n2158\
        );

    \I__258\ : InMux
    port map (
            O => \N__2768\,
            I => \uart.n2159\
        );

    \I__257\ : InMux
    port map (
            O => \N__2765\,
            I => \uart.n2160\
        );

    \I__256\ : InMux
    port map (
            O => \N__2762\,
            I => \uart.n2161\
        );

    \I__255\ : InMux
    port map (
            O => \N__2759\,
            I => \uart.n2162\
        );

    \I__254\ : InMux
    port map (
            O => \N__2756\,
            I => \uart.n2145\
        );

    \I__253\ : InMux
    port map (
            O => \N__2753\,
            I => \uart.n2146\
        );

    \I__252\ : InMux
    port map (
            O => \N__2750\,
            I => \bfn_1_20_0_\
        );

    \I__251\ : InMux
    port map (
            O => \N__2747\,
            I => \uart.n2148\
        );

    \I__250\ : InMux
    port map (
            O => \N__2744\,
            I => \uart.n2149\
        );

    \I__249\ : InMux
    port map (
            O => \N__2741\,
            I => \uart.n2150\
        );

    \I__248\ : InMux
    port map (
            O => \N__2738\,
            I => \uart.n2151\
        );

    \I__247\ : InMux
    port map (
            O => \N__2735\,
            I => \uart.n2152\
        );

    \I__246\ : InMux
    port map (
            O => \N__2732\,
            I => \uart.n2153\
        );

    \I__245\ : InMux
    port map (
            O => \N__2729\,
            I => \uart.n2135\
        );

    \I__244\ : InMux
    port map (
            O => \N__2726\,
            I => \uart.n2136\
        );

    \I__243\ : InMux
    port map (
            O => \N__2723\,
            I => \uart.n2137\
        );

    \I__242\ : InMux
    port map (
            O => \N__2720\,
            I => \uart.n2138\
        );

    \I__241\ : InMux
    port map (
            O => \N__2717\,
            I => \bfn_1_19_0_\
        );

    \I__240\ : InMux
    port map (
            O => \N__2714\,
            I => \uart.n2140\
        );

    \I__239\ : InMux
    port map (
            O => \N__2711\,
            I => \uart.n2141\
        );

    \I__238\ : InMux
    port map (
            O => \N__2708\,
            I => \uart.n2142\
        );

    \I__237\ : InMux
    port map (
            O => \N__2705\,
            I => \uart.n2143\
        );

    \I__236\ : InMux
    port map (
            O => \N__2702\,
            I => \uart.n2144\
        );

    \I__235\ : IoInMux
    port map (
            O => \N__2699\,
            I => \N__2696\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2696\,
            I => \N__2693\
        );

    \I__233\ : IoSpan4Mux
    port map (
            O => \N__2693\,
            I => \N__2690\
        );

    \I__232\ : IoSpan4Mux
    port map (
            O => \N__2690\,
            I => \N__2687\
        );

    \I__231\ : IoSpan4Mux
    port map (
            O => \N__2687\,
            I => \N__2684\
        );

    \I__230\ : Odrv4
    port map (
            O => \N__2684\,
            I => \CLK_pad_gb_input\
        );

    \I__229\ : InMux
    port map (
            O => \N__2681\,
            I => \bfn_1_18_0_\
        );

    \I__228\ : InMux
    port map (
            O => \N__2678\,
            I => \uart.n2132\
        );

    \I__227\ : InMux
    port map (
            O => \N__2675\,
            I => \uart.n2133\
        );

    \I__226\ : InMux
    port map (
            O => \N__2672\,
            I => \uart.n2134\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart.n2139\,
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart.n2147\,
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_1_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart.n2155\,
            carryinitout => \bfn_1_21_0_\
        );

    \IN_MUX_bfv_5_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_23_0_\
        );

    \IN_MUX_bfv_3_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_22_0_\
        );

    \IN_MUX_bfv_3_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2202,
            carryinitout => \bfn_3_23_0_\
        );

    \IN_MUX_bfv_3_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2210,
            carryinitout => \bfn_3_24_0_\
        );

    \IN_MUX_bfv_3_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2218,
            carryinitout => \bfn_3_25_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_1_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2233,
            carryinitout => \bfn_1_23_0_\
        );

    \IN_MUX_bfv_1_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2241,
            carryinitout => \bfn_1_24_0_\
        );

    \IN_MUX_bfv_1_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2249,
            carryinitout => \bfn_1_25_0_\
        );

    \IN_MUX_bfv_2_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_23_0_\
        );

    \IN_MUX_bfv_2_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2170,
            carryinitout => \bfn_2_24_0_\
        );

    \IN_MUX_bfv_2_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2178,
            carryinitout => \bfn_2_25_0_\
        );

    \IN_MUX_bfv_2_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2186,
            carryinitout => \bfn_2_26_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2699\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uart.r_Clock_Count_121__i0_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2986\,
            in2 => \_gnd_net_\,
            in3 => \N__2681\,
            lcout => \uart.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \uart.n2132\,
            clk => \N__5379\,
            ce => \N__3106\,
            sr => \N__3216\
        );

    \uart.r_Clock_Count_121__i1_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2974\,
            in2 => \_gnd_net_\,
            in3 => \N__2678\,
            lcout => \uart.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \uart.n2132\,
            carryout => \uart.n2133\,
            clk => \N__5379\,
            ce => \N__3106\,
            sr => \N__3216\
        );

    \uart.r_Clock_Count_121__i2_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2998\,
            in2 => \_gnd_net_\,
            in3 => \N__2675\,
            lcout => \uart.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \uart.n2133\,
            carryout => \uart.n2134\,
            clk => \N__5379\,
            ce => \N__3106\,
            sr => \N__3216\
        );

    \uart.r_Clock_Count_121__i3_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2960\,
            in2 => \_gnd_net_\,
            in3 => \N__2672\,
            lcout => \uart.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \uart.n2134\,
            carryout => \uart.n2135\,
            clk => \N__5379\,
            ce => \N__3106\,
            sr => \N__3216\
        );

    \uart.r_Clock_Count_121__i4_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2936\,
            in2 => \_gnd_net_\,
            in3 => \N__2729\,
            lcout => \uart.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \uart.n2135\,
            carryout => \uart.n2136\,
            clk => \N__5379\,
            ce => \N__3106\,
            sr => \N__3216\
        );

    \uart.r_Clock_Count_121__i5_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2948\,
            in2 => \_gnd_net_\,
            in3 => \N__2726\,
            lcout => \uart.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \uart.n2136\,
            carryout => \uart.n2137\,
            clk => \N__5379\,
            ce => \N__3106\,
            sr => \N__3216\
        );

    \uart.r_Clock_Count_121__i6_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2921\,
            in2 => \_gnd_net_\,
            in3 => \N__2723\,
            lcout => \uart.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \uart.n2137\,
            carryout => \uart.n2138\,
            clk => \N__5379\,
            ce => \N__3106\,
            sr => \N__3216\
        );

    \uart.r_Clock_Count_121__i7_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3248\,
            in2 => \_gnd_net_\,
            in3 => \N__2720\,
            lcout => \uart.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \uart.n2138\,
            carryout => \uart.n2139\,
            clk => \N__5379\,
            ce => \N__3106\,
            sr => \N__3216\
        );

    \uart.r_Clock_Count_121__i8_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3193\,
            in2 => \_gnd_net_\,
            in3 => \N__2717\,
            lcout => \uart.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \uart.n2140\,
            clk => \N__5380\,
            ce => \N__3095\,
            sr => \N__3215\
        );

    \uart.r_Clock_Count_121__i9_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3605\,
            in2 => \_gnd_net_\,
            in3 => \N__2714\,
            lcout => \uart.r_Clock_Count_9\,
            ltout => OPEN,
            carryin => \uart.n2140\,
            carryout => \uart.n2141\,
            clk => \N__5380\,
            ce => \N__3095\,
            sr => \N__3215\
        );

    \uart.r_Clock_Count_121__i10_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2909\,
            in2 => \_gnd_net_\,
            in3 => \N__2711\,
            lcout => \uart.r_Clock_Count_10\,
            ltout => OPEN,
            carryin => \uart.n2141\,
            carryout => \uart.n2142\,
            clk => \N__5380\,
            ce => \N__3095\,
            sr => \N__3215\
        );

    \uart.r_Clock_Count_121__i11_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3065\,
            in2 => \_gnd_net_\,
            in3 => \N__2708\,
            lcout => \uart.r_Clock_Count_11\,
            ltout => OPEN,
            carryin => \uart.n2142\,
            carryout => \uart.n2143\,
            clk => \N__5380\,
            ce => \N__3095\,
            sr => \N__3215\
        );

    \uart.r_Clock_Count_121__i12_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3278\,
            in2 => \_gnd_net_\,
            in3 => \N__2705\,
            lcout => \uart.r_Clock_Count_12\,
            ltout => OPEN,
            carryin => \uart.n2143\,
            carryout => \uart.n2144\,
            clk => \N__5380\,
            ce => \N__3095\,
            sr => \N__3215\
        );

    \uart.r_Clock_Count_121__i13_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3290\,
            in2 => \_gnd_net_\,
            in3 => \N__2702\,
            lcout => \uart.r_Clock_Count_13\,
            ltout => OPEN,
            carryin => \uart.n2144\,
            carryout => \uart.n2145\,
            clk => \N__5380\,
            ce => \N__3095\,
            sr => \N__3215\
        );

    \uart.r_Clock_Count_121__i14_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3179\,
            in2 => \_gnd_net_\,
            in3 => \N__2756\,
            lcout => \uart.r_Clock_Count_14\,
            ltout => OPEN,
            carryin => \uart.n2145\,
            carryout => \uart.n2146\,
            clk => \N__5380\,
            ce => \N__3095\,
            sr => \N__3215\
        );

    \uart.r_Clock_Count_121__i15_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3632\,
            in2 => \_gnd_net_\,
            in3 => \N__2753\,
            lcout => \uart.r_Clock_Count_15\,
            ltout => OPEN,
            carryin => \uart.n2146\,
            carryout => \uart.n2147\,
            clk => \N__5380\,
            ce => \N__3095\,
            sr => \N__3215\
        );

    \uart.r_Clock_Count_121__i16_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3565\,
            in2 => \_gnd_net_\,
            in3 => \N__2750\,
            lcout => \uart.r_Clock_Count_16\,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => \uart.n2148\,
            clk => \N__5381\,
            ce => \N__3094\,
            sr => \N__3217\
        );

    \uart.r_Clock_Count_121__i17_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3040\,
            in2 => \_gnd_net_\,
            in3 => \N__2747\,
            lcout => \uart.r_Clock_Count_17\,
            ltout => OPEN,
            carryin => \uart.n2148\,
            carryout => \uart.n2149\,
            clk => \N__5381\,
            ce => \N__3094\,
            sr => \N__3217\
        );

    \uart.r_Clock_Count_121__i18_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3026\,
            in2 => \_gnd_net_\,
            in3 => \N__2744\,
            lcout => \uart.r_Clock_Count_18\,
            ltout => OPEN,
            carryin => \uart.n2149\,
            carryout => \uart.n2150\,
            clk => \N__5381\,
            ce => \N__3094\,
            sr => \N__3217\
        );

    \uart.r_Clock_Count_121__i19_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3578\,
            in2 => \_gnd_net_\,
            in3 => \N__2741\,
            lcout => \uart.r_Clock_Count_19\,
            ltout => OPEN,
            carryin => \uart.n2150\,
            carryout => \uart.n2151\,
            clk => \N__5381\,
            ce => \N__3094\,
            sr => \N__3217\
        );

    \uart.r_Clock_Count_121__i20_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3644\,
            in2 => \_gnd_net_\,
            in3 => \N__2738\,
            lcout => \uart.r_Clock_Count_20\,
            ltout => OPEN,
            carryin => \uart.n2151\,
            carryout => \uart.n2152\,
            clk => \N__5381\,
            ce => \N__3094\,
            sr => \N__3217\
        );

    \uart.r_Clock_Count_121__i21_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3053\,
            in2 => \_gnd_net_\,
            in3 => \N__2735\,
            lcout => \uart.r_Clock_Count_21\,
            ltout => OPEN,
            carryin => \uart.n2152\,
            carryout => \uart.n2153\,
            clk => \N__5381\,
            ce => \N__3094\,
            sr => \N__3217\
        );

    \uart.r_Clock_Count_121__i22_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2897\,
            in2 => \_gnd_net_\,
            in3 => \N__2732\,
            lcout => \uart.r_Clock_Count_22\,
            ltout => OPEN,
            carryin => \uart.n2153\,
            carryout => \uart.n2154\,
            clk => \N__5381\,
            ce => \N__3094\,
            sr => \N__3217\
        );

    \uart.r_Clock_Count_121__i23_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3119\,
            in2 => \_gnd_net_\,
            in3 => \N__2783\,
            lcout => \uart.r_Clock_Count_23\,
            ltout => OPEN,
            carryin => \uart.n2154\,
            carryout => \uart.n2155\,
            clk => \N__5381\,
            ce => \N__3094\,
            sr => \N__3217\
        );

    \uart.r_Clock_Count_121__i24_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3133\,
            in2 => \_gnd_net_\,
            in3 => \N__2780\,
            lcout => \uart.r_Clock_Count_24\,
            ltout => OPEN,
            carryin => \bfn_1_21_0_\,
            carryout => \uart.n2156\,
            clk => \N__5383\,
            ce => \N__3096\,
            sr => \N__3224\
        );

    \uart.r_Clock_Count_121__i25_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3619\,
            in2 => \_gnd_net_\,
            in3 => \N__2777\,
            lcout => \uart.r_Clock_Count_25\,
            ltout => OPEN,
            carryin => \uart.n2156\,
            carryout => \uart.n2157\,
            clk => \N__5383\,
            ce => \N__3096\,
            sr => \N__3224\
        );

    \uart.r_Clock_Count_121__i26_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2878\,
            in2 => \_gnd_net_\,
            in3 => \N__2774\,
            lcout => \uart.r_Clock_Count_26\,
            ltout => OPEN,
            carryin => \uart.n2157\,
            carryout => \uart.n2158\,
            clk => \N__5383\,
            ce => \N__3096\,
            sr => \N__3224\
        );

    \uart.r_Clock_Count_121__i27_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3592\,
            in2 => \_gnd_net_\,
            in3 => \N__2771\,
            lcout => \uart.r_Clock_Count_27\,
            ltout => OPEN,
            carryin => \uart.n2158\,
            carryout => \uart.n2159\,
            clk => \N__5383\,
            ce => \N__3096\,
            sr => \N__3224\
        );

    \uart.r_Clock_Count_121__i28_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3149\,
            in2 => \_gnd_net_\,
            in3 => \N__2768\,
            lcout => \uart.r_Clock_Count_28\,
            ltout => OPEN,
            carryin => \uart.n2159\,
            carryout => \uart.n2160\,
            clk => \N__5383\,
            ce => \N__3096\,
            sr => \N__3224\
        );

    \uart.r_Clock_Count_121__i29_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3265\,
            in2 => \_gnd_net_\,
            in3 => \N__2765\,
            lcout => \uart.r_Clock_Count_29\,
            ltout => OPEN,
            carryin => \uart.n2160\,
            carryout => \uart.n2161\,
            clk => \N__5383\,
            ce => \N__3096\,
            sr => \N__3224\
        );

    \uart.r_Clock_Count_121__i30_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3161\,
            in2 => \_gnd_net_\,
            in3 => \N__2762\,
            lcout => \uart.r_Clock_Count_30\,
            ltout => OPEN,
            carryin => \uart.n2161\,
            carryout => \uart.n2162\,
            clk => \N__5383\,
            ce => \N__3096\,
            sr => \N__3224\
        );

    \uart.r_Clock_Count_121__i31_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3551\,
            in2 => \_gnd_net_\,
            in3 => \N__2759\,
            lcout => \uart.r_Clock_Count_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5383\,
            ce => \N__3096\,
            sr => \N__3224\
        );

    \clk_divider_116__i0_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3974\,
            in2 => \_gnd_net_\,
            in3 => \N__2810\,
            lcout => clk_divider_0,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => n2226,
            clk => \N__5385\,
            ce => 'H',
            sr => \N__3938\
        );

    \clk_divider_116__i1_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3899\,
            in2 => \_gnd_net_\,
            in3 => \N__2807\,
            lcout => clk_divider_1,
            ltout => OPEN,
            carryin => n2226,
            carryout => n2227,
            clk => \N__5385\,
            ce => 'H',
            sr => \N__3938\
        );

    \clk_divider_116__i2_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3887\,
            in2 => \_gnd_net_\,
            in3 => \N__2804\,
            lcout => clk_divider_2,
            ltout => OPEN,
            carryin => n2227,
            carryout => n2228,
            clk => \N__5385\,
            ce => 'H',
            sr => \N__3938\
        );

    \clk_divider_116__i3_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3961\,
            in2 => \_gnd_net_\,
            in3 => \N__2801\,
            lcout => clk_divider_3,
            ltout => OPEN,
            carryin => n2228,
            carryout => n2229,
            clk => \N__5385\,
            ce => 'H',
            sr => \N__3938\
        );

    \clk_divider_116__i4_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3988\,
            in2 => \_gnd_net_\,
            in3 => \N__2798\,
            lcout => clk_divider_4,
            ltout => OPEN,
            carryin => n2229,
            carryout => n2230,
            clk => \N__5385\,
            ce => 'H',
            sr => \N__3938\
        );

    \clk_divider_116__i5_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3815\,
            in2 => \_gnd_net_\,
            in3 => \N__2795\,
            lcout => clk_divider_5,
            ltout => OPEN,
            carryin => n2230,
            carryout => n2231,
            clk => \N__5385\,
            ce => 'H',
            sr => \N__3938\
        );

    \clk_divider_116__i6_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3386\,
            in2 => \_gnd_net_\,
            in3 => \N__2792\,
            lcout => clk_divider_6,
            ltout => OPEN,
            carryin => n2231,
            carryout => n2232,
            clk => \N__5385\,
            ce => 'H',
            sr => \N__3938\
        );

    \clk_divider_116__i7_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4246\,
            in2 => \_gnd_net_\,
            in3 => \N__2789\,
            lcout => clk_divider_7,
            ltout => OPEN,
            carryin => n2232,
            carryout => n2233,
            clk => \N__5385\,
            ce => 'H',
            sr => \N__3938\
        );

    \clk_divider_116__i8_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3869\,
            in2 => \_gnd_net_\,
            in3 => \N__2786\,
            lcout => clk_divider_8,
            ltout => OPEN,
            carryin => \bfn_1_23_0_\,
            carryout => n2234,
            clk => \N__5388\,
            ce => 'H',
            sr => \N__3942\
        );

    \clk_divider_116__i9_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3490\,
            in2 => \_gnd_net_\,
            in3 => \N__2837\,
            lcout => clk_divider_9,
            ltout => OPEN,
            carryin => n2234,
            carryout => n2235,
            clk => \N__5388\,
            ce => 'H',
            sr => \N__3942\
        );

    \clk_divider_116__i10_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3803\,
            in2 => \_gnd_net_\,
            in3 => \N__2834\,
            lcout => clk_divider_10,
            ltout => OPEN,
            carryin => n2235,
            carryout => n2236,
            clk => \N__5388\,
            ce => 'H',
            sr => \N__3942\
        );

    \clk_divider_116__i11_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3827\,
            in2 => \_gnd_net_\,
            in3 => \N__2831\,
            lcout => clk_divider_11,
            ltout => OPEN,
            carryin => n2236,
            carryout => n2237,
            clk => \N__5388\,
            ce => 'H',
            sr => \N__3942\
        );

    \clk_divider_116__i12_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3790\,
            in2 => \_gnd_net_\,
            in3 => \N__2828\,
            lcout => clk_divider_12,
            ltout => OPEN,
            carryin => n2237,
            carryout => n2238,
            clk => \N__5388\,
            ce => 'H',
            sr => \N__3942\
        );

    \clk_divider_116__i13_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3761\,
            in2 => \_gnd_net_\,
            in3 => \N__2825\,
            lcout => clk_divider_13,
            ltout => OPEN,
            carryin => n2238,
            carryout => n2239,
            clk => \N__5388\,
            ce => 'H',
            sr => \N__3942\
        );

    \clk_divider_116__i14_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3472\,
            in2 => \_gnd_net_\,
            in3 => \N__2822\,
            lcout => clk_divider_14,
            ltout => OPEN,
            carryin => n2239,
            carryout => n2240,
            clk => \N__5388\,
            ce => 'H',
            sr => \N__3942\
        );

    \clk_divider_116__i15_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3857\,
            in2 => \_gnd_net_\,
            in3 => \N__2819\,
            lcout => clk_divider_15,
            ltout => OPEN,
            carryin => n2240,
            carryout => n2241,
            clk => \N__5388\,
            ce => 'H',
            sr => \N__3942\
        );

    \clk_divider_116__i16_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3712\,
            in2 => \_gnd_net_\,
            in3 => \N__2816\,
            lcout => clk_divider_16,
            ltout => OPEN,
            carryin => \bfn_1_24_0_\,
            carryout => n2242,
            clk => \N__5392\,
            ce => 'H',
            sr => \N__3946\
        );

    \clk_divider_116__i17_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3454\,
            in2 => \_gnd_net_\,
            in3 => \N__2813\,
            lcout => clk_divider_17,
            ltout => OPEN,
            carryin => n2242,
            carryout => n2243,
            clk => \N__5392\,
            ce => 'H',
            sr => \N__3946\
        );

    \clk_divider_116__i18_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3775\,
            in2 => \_gnd_net_\,
            in3 => \N__2864\,
            lcout => clk_divider_18,
            ltout => OPEN,
            carryin => n2243,
            carryout => n2244,
            clk => \N__5392\,
            ce => 'H',
            sr => \N__3946\
        );

    \clk_divider_116__i19_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3319\,
            in2 => \_gnd_net_\,
            in3 => \N__2861\,
            lcout => clk_divider_19,
            ltout => OPEN,
            carryin => n2244,
            carryout => n2245,
            clk => \N__5392\,
            ce => 'H',
            sr => \N__3946\
        );

    \clk_divider_116__i20_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3334\,
            in2 => \_gnd_net_\,
            in3 => \N__2858\,
            lcout => clk_divider_20,
            ltout => OPEN,
            carryin => n2245,
            carryout => n2246,
            clk => \N__5392\,
            ce => 'H',
            sr => \N__3946\
        );

    \clk_divider_116__i21_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3439\,
            in2 => \_gnd_net_\,
            in3 => \N__2855\,
            lcout => clk_divider_21,
            ltout => OPEN,
            carryin => n2246,
            carryout => n2247,
            clk => \N__5392\,
            ce => 'H',
            sr => \N__3946\
        );

    \clk_divider_116__i22_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3421\,
            in2 => \_gnd_net_\,
            in3 => \N__2852\,
            lcout => clk_divider_22,
            ltout => OPEN,
            carryin => n2247,
            carryout => n2248,
            clk => \N__5392\,
            ce => 'H',
            sr => \N__3946\
        );

    \clk_divider_116__i23_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3727\,
            in2 => \_gnd_net_\,
            in3 => \N__2849\,
            lcout => clk_divider_23,
            ltout => OPEN,
            carryin => n2248,
            carryout => n2249,
            clk => \N__5392\,
            ce => 'H',
            sr => \N__3946\
        );

    \clk_divider_116__i24_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3841\,
            in2 => \_gnd_net_\,
            in3 => \N__2846\,
            lcout => clk_divider_24,
            ltout => OPEN,
            carryin => \bfn_1_25_0_\,
            carryout => n2250,
            clk => \N__5395\,
            ce => 'H',
            sr => \N__3947\
        );

    \clk_divider_116__i25_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4219\,
            in2 => \_gnd_net_\,
            in3 => \N__2843\,
            lcout => clk_divider_25,
            ltout => OPEN,
            carryin => n2250,
            carryout => n2251,
            clk => \N__5395\,
            ce => 'H',
            sr => \N__3947\
        );

    \clk_divider_116__i26_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3505\,
            in2 => \_gnd_net_\,
            in3 => \N__2840\,
            lcout => clk_divider_26,
            ltout => OPEN,
            carryin => n2251,
            carryout => n2252,
            clk => \N__5395\,
            ce => 'H',
            sr => \N__3947\
        );

    \clk_divider_116__i27_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3352\,
            in2 => \_gnd_net_\,
            in3 => \N__3014\,
            lcout => clk_divider_27,
            ltout => OPEN,
            carryin => n2252,
            carryout => n2253,
            clk => \N__5395\,
            ce => 'H',
            sr => \N__3947\
        );

    \clk_divider_116__i28_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3400\,
            in2 => \_gnd_net_\,
            in3 => \N__3011\,
            lcout => clk_divider_28,
            ltout => OPEN,
            carryin => n2253,
            carryout => n2254,
            clk => \N__5395\,
            ce => 'H',
            sr => \N__3947\
        );

    \clk_divider_116__i29_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3748\,
            in2 => \_gnd_net_\,
            in3 => \N__3008\,
            lcout => clk_divider_29,
            ltout => OPEN,
            carryin => n2254,
            carryout => n2255,
            clk => \N__5395\,
            ce => 'H',
            sr => \N__3947\
        );

    \clk_divider_116__i30_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3370\,
            in2 => \_gnd_net_\,
            in3 => \N__3005\,
            lcout => clk_divider_30,
            ltout => OPEN,
            carryin => n2255,
            carryout => n2256,
            clk => \N__5395\,
            ce => 'H',
            sr => \N__3947\
        );

    \clk_divider_116__i31_LC_1_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3682\,
            in2 => \_gnd_net_\,
            in3 => \N__3002\,
            lcout => clk_divider_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5395\,
            ce => 'H',
            sr => \N__3947\
        );

    \uart.i806_4_lut_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__2999\,
            in1 => \N__2987\,
            in2 => \N__2975\,
            in3 => \N__2959\,
            lcout => OPEN,
            ltout => \uart.n2006_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i3_4_lut_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2947\,
            in1 => \N__2935\,
            in2 => \N__2924\,
            in3 => \N__2920\,
            lcout => \uart.n2385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_SM_Main_i2_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4547\,
            in1 => \N__4678\,
            in2 => \N__4732\,
            in3 => \N__4630\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i18_4_lut_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2908\,
            in1 => \N__2896\,
            in2 => \N__2885\,
            in3 => \N__3289\,
            lcout => OPEN,
            ltout => \uart.n42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i21_4_lut_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3277\,
            in1 => \N__3266\,
            in2 => \N__3251\,
            in3 => \N__3167\,
            lcout => OPEN,
            ltout => \uart.n45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i1_4_lut_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__3518\,
            in1 => \N__3247\,
            in2 => \N__3236\,
            in3 => \N__3233\,
            lcout => \r_SM_Main_2_N_233_1\,
            ltout => \r_SM_Main_2_N_233_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i1088_4_lut_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110001"
        )
    port map (
            in0 => \N__4721\,
            in1 => \N__4677\,
            in2 => \N__3227\,
            in3 => \N__4629\,
            lcout => \uart.n1796\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i10_2_lut_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3194\,
            in3 => \N__3178\,
            lcout => \uart.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i515_4_lut_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__4520\,
            in1 => \N__4720\,
            in2 => \N__5099\,
            in3 => \N__4546\,
            lcout => \uart.n1711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i15_4_lut_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3160\,
            in1 => \N__3148\,
            in2 => \N__3137\,
            in3 => \N__3118\,
            lcout => \uart.n39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i1_1_lut_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4631\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i16_4_lut_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3064\,
            in1 => \N__3052\,
            in2 => \N__3041\,
            in3 => \N__3025\,
            lcout => \uart.n40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i14_4_lut_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3643\,
            in1 => \N__3631\,
            in2 => \N__3620\,
            in3 => \N__3604\,
            lcout => \uart.n38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i13_4_lut_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3593\,
            in1 => \N__3577\,
            in2 => \N__3566\,
            in3 => \N__3550\,
            lcout => OPEN,
            ltout => \uart.n37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i22_4_lut_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3539\,
            in1 => \N__3533\,
            in2 => \N__3527\,
            in3 => \N__3524\,
            lcout => \uart.n46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18_4_lut_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3509\,
            in1 => \N__3491\,
            in2 => \N__3476\,
            in3 => \N__3458\,
            lcout => n44_adj_358,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_1_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3440\,
            in1 => \N__3425\,
            in2 => \N__3407\,
            in3 => \N__3385\,
            lcout => n41_adj_361,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16_4_lut_adj_2_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3374\,
            in1 => \N__3356\,
            in2 => \N__3338\,
            in3 => \N__3320\,
            lcout => OPEN,
            ltout => \n42_adj_360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3305\,
            in1 => \N__3698\,
            in2 => \N__3299\,
            in3 => \N__3296\,
            lcout => n50,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i291_4_lut_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__3989\,
            in1 => \N__3973\,
            in2 => \N__3962\,
            in3 => \N__3875\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i708_4_lut_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__3655\,
            in1 => \N__3664\,
            in2 => \N__3692\,
            in3 => \N__4198\,
            lcout => \clk_divider_31__N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_SM_Main_2__I_0_62_i3_3_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011101"
        )
    port map (
            in0 => \N__4736\,
            in1 => \N__4256\,
            in2 => \_gnd_net_\,
            in3 => \N__4679\,
            lcout => \uart.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3898\,
            in2 => \_gnd_net_\,
            in3 => \N__3886\,
            lcout => n6_adj_324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_adj_4_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3868\,
            in1 => \N__3856\,
            in2 => \N__3845\,
            in3 => \N__3826\,
            lcout => n40_adj_362,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3814\,
            in1 => \N__3802\,
            in2 => \N__3791\,
            in3 => \N__3776\,
            lcout => n45_adj_357,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i17_4_lut_adj_3_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3760\,
            in1 => \N__3749\,
            in2 => \N__3734\,
            in3 => \N__3713\,
            lcout => n43_adj_359,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_slow_25_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__4199\,
            in1 => \N__3691\,
            in2 => \N__3668\,
            in3 => \N__3656\,
            lcout => clk_slow,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i0_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4061\,
            in2 => \_gnd_net_\,
            in3 => \N__4055\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_2_23_0_\,
            carryout => n2163,
            clk => \N__5393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i1_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4052\,
            in2 => \_gnd_net_\,
            in3 => \N__4046\,
            lcout => n25,
            ltout => OPEN,
            carryin => n2163,
            carryout => n2164,
            clk => \N__5393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i2_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4043\,
            in2 => \_gnd_net_\,
            in3 => \N__4037\,
            lcout => n24,
            ltout => OPEN,
            carryin => n2164,
            carryout => n2165,
            clk => \N__5393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i3_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4034\,
            in2 => \_gnd_net_\,
            in3 => \N__4028\,
            lcout => n23,
            ltout => OPEN,
            carryin => n2165,
            carryout => n2166,
            clk => \N__5393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i4_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4025\,
            in2 => \_gnd_net_\,
            in3 => \N__4019\,
            lcout => n22,
            ltout => OPEN,
            carryin => n2166,
            carryout => n2167,
            clk => \N__5393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i5_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4016\,
            in2 => \_gnd_net_\,
            in3 => \N__4010\,
            lcout => n21,
            ltout => OPEN,
            carryin => n2167,
            carryout => n2168,
            clk => \N__5393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i6_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4007\,
            in2 => \_gnd_net_\,
            in3 => \N__4001\,
            lcout => n20,
            ltout => OPEN,
            carryin => n2168,
            carryout => n2169,
            clk => \N__5393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i7_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3998\,
            in2 => \_gnd_net_\,
            in3 => \N__3992\,
            lcout => n19,
            ltout => OPEN,
            carryin => n2169,
            carryout => n2170,
            clk => \N__5393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i8_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4142\,
            in2 => \_gnd_net_\,
            in3 => \N__4136\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_2_24_0_\,
            carryout => n2171,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i9_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4133\,
            in2 => \_gnd_net_\,
            in3 => \N__4127\,
            lcout => n17,
            ltout => OPEN,
            carryin => n2171,
            carryout => n2172,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i10_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4124\,
            in2 => \_gnd_net_\,
            in3 => \N__4118\,
            lcout => n16,
            ltout => OPEN,
            carryin => n2172,
            carryout => n2173,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i11_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4115\,
            in2 => \_gnd_net_\,
            in3 => \N__4109\,
            lcout => n15,
            ltout => OPEN,
            carryin => n2173,
            carryout => n2174,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i12_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4106\,
            in2 => \_gnd_net_\,
            in3 => \N__4100\,
            lcout => n14,
            ltout => OPEN,
            carryin => n2174,
            carryout => n2175,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i13_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4097\,
            in2 => \_gnd_net_\,
            in3 => \N__4091\,
            lcout => n13,
            ltout => OPEN,
            carryin => n2175,
            carryout => n2176,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i14_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4088\,
            in2 => \_gnd_net_\,
            in3 => \N__4082\,
            lcout => n12,
            ltout => OPEN,
            carryin => n2176,
            carryout => n2177,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i15_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4079\,
            in2 => \_gnd_net_\,
            in3 => \N__4073\,
            lcout => n11,
            ltout => OPEN,
            carryin => n2177,
            carryout => n2178,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i16_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4070\,
            in2 => \_gnd_net_\,
            in3 => \N__4064\,
            lcout => n10_adj_317,
            ltout => OPEN,
            carryin => \bfn_2_25_0_\,
            carryout => n2179,
            clk => \N__5397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i17_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4190\,
            in2 => \_gnd_net_\,
            in3 => \N__4184\,
            lcout => n9,
            ltout => OPEN,
            carryin => n2179,
            carryout => n2180,
            clk => \N__5397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i18_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4181\,
            in2 => \_gnd_net_\,
            in3 => \N__4175\,
            lcout => n8,
            ltout => OPEN,
            carryin => n2180,
            carryout => n2181,
            clk => \N__5397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i19_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4172\,
            in2 => \_gnd_net_\,
            in3 => \N__4166\,
            lcout => n7,
            ltout => OPEN,
            carryin => n2181,
            carryout => n2182,
            clk => \N__5397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i20_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4163\,
            in2 => \_gnd_net_\,
            in3 => \N__4157\,
            lcout => n6,
            ltout => OPEN,
            carryin => n2182,
            carryout => n2183,
            clk => \N__5397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i21_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4336\,
            in2 => \_gnd_net_\,
            in3 => \N__4154\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n2183,
            carryout => n2184,
            clk => \N__5397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i22_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4279\,
            in2 => \_gnd_net_\,
            in3 => \N__4151\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n2184,
            carryout => n2185,
            clk => \N__5397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i23_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4297\,
            in2 => \_gnd_net_\,
            in3 => \N__4148\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n2185,
            carryout => n2186,
            clk => \N__5397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i24_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4323\,
            in2 => \_gnd_net_\,
            in3 => \N__4145\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_2_26_0_\,
            carryout => n2187,
            clk => \N__5398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_119__i25_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4372\,
            in2 => \_gnd_net_\,
            in3 => \N__4376\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1070_4_lut_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111000"
        )
    port map (
            in0 => \N__4343\,
            in1 => \N__4325\,
            in2 => \N__4310\,
            in3 => \N__4286\,
            lcout => OPEN,
            ltout => \n2395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1071_3_lut_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__4373\,
            in1 => \_gnd_net_\,
            in2 => \N__4361\,
            in3 => \N__4268\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1069_4_lut_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000100010"
        )
    port map (
            in0 => \N__4342\,
            in1 => \N__4324\,
            in2 => \N__4309\,
            in3 => \N__4285\,
            lcout => n2394,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_SM_Main_i0_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__4549\,
            in1 => \N__4672\,
            in2 => \_gnd_net_\,
            in3 => \N__4262\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5384\,
            ce => 'H',
            sr => \N__4636\
        );

    \uart.r_SM_Main_i1_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4673\,
            in1 => \N__4729\,
            in2 => \_gnd_net_\,
            in3 => \N__4548\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5384\,
            ce => 'H',
            sr => \N__4636\
        );

    \uart.r_Bit_Index_i2_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__4571\,
            in1 => \N__5447\,
            in2 => \_gnd_net_\,
            in3 => \N__5477\,
            lcout => \uart.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5386\,
            ce => \N__5329\,
            sr => \N__5302\
        );

    \uart.i8225_i1_3_lut_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4570\,
            in1 => \N__4751\,
            in2 => \_gnd_net_\,
            in3 => \N__4778\,
            lcout => \uart.o_Tx_Serial_N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i23_4_lut_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4250\,
            in1 => \N__4232\,
            in2 => \N__4226\,
            in3 => \N__4205\,
            lcout => n49,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_117__i0_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4448\,
            in2 => \_gnd_net_\,
            in3 => \N__4442\,
            lcout => counter_0,
            ltout => OPEN,
            carryin => \bfn_3_22_0_\,
            carryout => n2195,
            clk => \N__5754\,
            ce => 'H',
            sr => \N__5709\
        );

    \counter_117__i1_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4439\,
            in2 => \_gnd_net_\,
            in3 => \N__4433\,
            lcout => counter_1,
            ltout => OPEN,
            carryin => n2195,
            carryout => n2196,
            clk => \N__5754\,
            ce => 'H',
            sr => \N__5709\
        );

    \counter_117__i2_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4430\,
            in2 => \_gnd_net_\,
            in3 => \N__4424\,
            lcout => counter_2,
            ltout => OPEN,
            carryin => n2196,
            carryout => n2197,
            clk => \N__5754\,
            ce => 'H',
            sr => \N__5709\
        );

    \counter_117__i3_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4421\,
            in2 => \_gnd_net_\,
            in3 => \N__4415\,
            lcout => counter_3,
            ltout => OPEN,
            carryin => n2197,
            carryout => n2198,
            clk => \N__5754\,
            ce => 'H',
            sr => \N__5709\
        );

    \counter_117__i4_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4412\,
            in2 => \_gnd_net_\,
            in3 => \N__4406\,
            lcout => counter_4,
            ltout => OPEN,
            carryin => n2198,
            carryout => n2199,
            clk => \N__5754\,
            ce => 'H',
            sr => \N__5709\
        );

    \counter_117__i5_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4403\,
            in2 => \_gnd_net_\,
            in3 => \N__4397\,
            lcout => counter_5,
            ltout => OPEN,
            carryin => n2199,
            carryout => n2200,
            clk => \N__5754\,
            ce => 'H',
            sr => \N__5709\
        );

    \counter_117__i6_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4394\,
            in2 => \_gnd_net_\,
            in3 => \N__4388\,
            lcout => counter_6,
            ltout => OPEN,
            carryin => n2200,
            carryout => n2201,
            clk => \N__5754\,
            ce => 'H',
            sr => \N__5709\
        );

    \counter_117__i7_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4385\,
            in2 => \_gnd_net_\,
            in3 => \N__4379\,
            lcout => counter_7,
            ltout => OPEN,
            carryin => n2201,
            carryout => n2202,
            clk => \N__5754\,
            ce => 'H',
            sr => \N__5709\
        );

    \counter_117__i8_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4988\,
            in2 => \_gnd_net_\,
            in3 => \N__4475\,
            lcout => counter_8,
            ltout => OPEN,
            carryin => \bfn_3_23_0_\,
            carryout => n2203,
            clk => \N__5812\,
            ce => 'H',
            sr => \N__5707\
        );

    \counter_117__i9_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5510\,
            in2 => \_gnd_net_\,
            in3 => \N__4472\,
            lcout => counter_9,
            ltout => OPEN,
            carryin => n2203,
            carryout => n2204,
            clk => \N__5812\,
            ce => 'H',
            sr => \N__5707\
        );

    \counter_117__i10_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5579\,
            in2 => \_gnd_net_\,
            in3 => \N__4469\,
            lcout => counter_10,
            ltout => OPEN,
            carryin => n2204,
            carryout => n2205,
            clk => \N__5812\,
            ce => 'H',
            sr => \N__5707\
        );

    \counter_117__i11_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5176\,
            in2 => \_gnd_net_\,
            in3 => \N__4466\,
            lcout => counter_11,
            ltout => OPEN,
            carryin => n2205,
            carryout => n2206,
            clk => \N__5812\,
            ce => 'H',
            sr => \N__5707\
        );

    \counter_117__i12_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5000\,
            in2 => \_gnd_net_\,
            in3 => \N__4463\,
            lcout => counter_12,
            ltout => OPEN,
            carryin => n2206,
            carryout => n2207,
            clk => \N__5812\,
            ce => 'H',
            sr => \N__5707\
        );

    \counter_117__i13_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5203\,
            in2 => \_gnd_net_\,
            in3 => \N__4460\,
            lcout => counter_13,
            ltout => OPEN,
            carryin => n2207,
            carryout => n2208,
            clk => \N__5812\,
            ce => 'H',
            sr => \N__5707\
        );

    \counter_117__i14_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5162\,
            in2 => \_gnd_net_\,
            in3 => \N__4457\,
            lcout => counter_14,
            ltout => OPEN,
            carryin => n2208,
            carryout => n2209,
            clk => \N__5812\,
            ce => 'H',
            sr => \N__5707\
        );

    \counter_117__i15_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4975\,
            in2 => \_gnd_net_\,
            in3 => \N__4454\,
            lcout => counter_15,
            ltout => OPEN,
            carryin => n2209,
            carryout => n2210,
            clk => \N__5812\,
            ce => 'H',
            sr => \N__5707\
        );

    \counter_117__i16_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5612\,
            in2 => \_gnd_net_\,
            in3 => \N__4451\,
            lcout => counter_16,
            ltout => OPEN,
            carryin => \bfn_3_24_0_\,
            carryout => n2211,
            clk => \N__5814\,
            ce => 'H',
            sr => \N__5710\
        );

    \counter_117__i17_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5651\,
            in2 => \_gnd_net_\,
            in3 => \N__4505\,
            lcout => counter_17,
            ltout => OPEN,
            carryin => n2211,
            carryout => n2212,
            clk => \N__5814\,
            ce => 'H',
            sr => \N__5710\
        );

    \counter_117__i18_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5534\,
            in2 => \_gnd_net_\,
            in3 => \N__4502\,
            lcout => counter_18,
            ltout => OPEN,
            carryin => n2212,
            carryout => n2213,
            clk => \N__5814\,
            ce => 'H',
            sr => \N__5710\
        );

    \counter_117__i19_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5032\,
            in2 => \_gnd_net_\,
            in3 => \N__4499\,
            lcout => counter_19,
            ltout => OPEN,
            carryin => n2213,
            carryout => n2214,
            clk => \N__5814\,
            ce => 'H',
            sr => \N__5710\
        );

    \counter_117__i20_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5591\,
            in2 => \_gnd_net_\,
            in3 => \N__4496\,
            lcout => counter_20,
            ltout => OPEN,
            carryin => n2214,
            carryout => n2215,
            clk => \N__5814\,
            ce => 'H',
            sr => \N__5710\
        );

    \counter_117__i21_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5626\,
            in2 => \_gnd_net_\,
            in3 => \N__4493\,
            lcout => counter_21,
            ltout => OPEN,
            carryin => n2215,
            carryout => n2216,
            clk => \N__5814\,
            ce => 'H',
            sr => \N__5710\
        );

    \counter_117__i22_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5057\,
            in2 => \_gnd_net_\,
            in3 => \N__4490\,
            lcout => counter_22,
            ltout => OPEN,
            carryin => n2216,
            carryout => n2217,
            clk => \N__5814\,
            ce => 'H',
            sr => \N__5710\
        );

    \counter_117__i23_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5189\,
            in2 => \_gnd_net_\,
            in3 => \N__4487\,
            lcout => counter_23,
            ltout => OPEN,
            carryin => n2217,
            carryout => n2218,
            clk => \N__5814\,
            ce => 'H',
            sr => \N__5710\
        );

    \counter_117__i24_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5639\,
            in2 => \_gnd_net_\,
            in3 => \N__4484\,
            lcout => counter_24,
            ltout => OPEN,
            carryin => \bfn_3_25_0_\,
            carryout => n2219,
            clk => \N__5813\,
            ce => 'H',
            sr => \N__5717\
        );

    \counter_117__i25_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4961\,
            in2 => \_gnd_net_\,
            in3 => \N__4481\,
            lcout => counter_25,
            ltout => OPEN,
            carryin => n2219,
            carryout => n2220,
            clk => \N__5813\,
            ce => 'H',
            sr => \N__5717\
        );

    \counter_117__i26_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5018\,
            in2 => \_gnd_net_\,
            in3 => \N__4478\,
            lcout => counter_26,
            ltout => OPEN,
            carryin => n2220,
            carryout => n2221,
            clk => \N__5813\,
            ce => 'H',
            sr => \N__5717\
        );

    \counter_117__i27_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5522\,
            in2 => \_gnd_net_\,
            in3 => \N__4586\,
            lcout => counter_27,
            ltout => OPEN,
            carryin => n2221,
            carryout => n2222,
            clk => \N__5813\,
            ce => 'H',
            sr => \N__5717\
        );

    \counter_117__i28_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5552\,
            in2 => \_gnd_net_\,
            in3 => \N__4583\,
            lcout => counter_28,
            ltout => OPEN,
            carryin => n2222,
            carryout => n2223,
            clk => \N__5813\,
            ce => 'H',
            sr => \N__5717\
        );

    \counter_117__i29_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5566\,
            in2 => \_gnd_net_\,
            in3 => \N__4580\,
            lcout => counter_29,
            ltout => OPEN,
            carryin => n2223,
            carryout => n2224,
            clk => \N__5813\,
            ce => 'H',
            sr => \N__5717\
        );

    \counter_117__i30_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5045\,
            in2 => \_gnd_net_\,
            in3 => \N__4577\,
            lcout => counter_30,
            ltout => OPEN,
            carryin => n2224,
            carryout => n2225,
            clk => \N__5813\,
            ce => 'H',
            sr => \N__5717\
        );

    \counter_117__i31_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5119\,
            in2 => \_gnd_net_\,
            in3 => \N__4574\,
            lcout => counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5813\,
            ce => 'H',
            sr => \N__5717\
        );

    \uart.i2_3_lut_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4569\,
            in1 => \N__5437\,
            in2 => \_gnd_net_\,
            in3 => \N__5474\,
            lcout => n2002,
            ltout => \n2002_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Bit_Index_i0_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010010101010"
        )
    port map (
            in0 => \N__5475\,
            in1 => \N__4730\,
            in2 => \N__4553\,
            in3 => \N__5319\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i1095_3_lut_4_lut_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__4662\,
            in1 => \N__4632\,
            in2 => \N__4731\,
            in3 => \N__4550\,
            lcout => n2308,
            ltout => \n2308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i1091_2_lut_3_lut_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4719\,
            in2 => \N__4523\,
            in3 => \N__4519\,
            lcout => \uart.n2310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Tx_Data_i4_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5141\,
            in1 => \N__4888\,
            in2 => \_gnd_net_\,
            in3 => \N__4772\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Bit_Index_0__bdd_4_lut_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__4930\,
            in1 => \N__4864\,
            in2 => \N__5442\,
            in3 => \N__5472\,
            lcout => OPEN,
            ltout => \uart.n2428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.n2428_bdd_4_lut_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__4906\,
            in1 => \N__5432\,
            in2 => \N__4781\,
            in3 => \N__4597\,
            lcout => \uart.n2431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Tx_Data_i5_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4889\,
            in1 => \N__4853\,
            in2 => \_gnd_net_\,
            in3 => \N__4763\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Bit_Index_0__bdd_4_lut_1104_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__5473\,
            in1 => \N__4918\,
            in2 => \N__5443\,
            in3 => \N__4744\,
            lcout => OPEN,
            ltout => \uart.n2422_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.n2422_bdd_4_lut_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__4771\,
            in1 => \N__4762\,
            in2 => \N__4754\,
            in3 => \N__5436\,
            lcout => \uart.n2425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Tx_Data_i6_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5072\,
            in1 => \N__4890\,
            in2 => \_gnd_net_\,
            in3 => \N__4745\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.i2_3_lut_4_lut_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4725\,
            in1 => \N__4663\,
            in2 => \N__5092\,
            in3 => \N__4637\,
            lcout => n1757,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Tx_Data_i1_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4811\,
            in1 => \N__4892\,
            in2 => \_gnd_net_\,
            in3 => \N__4598\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Tx_Data_i3_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4894\,
            in1 => \N__4823\,
            in2 => \_gnd_net_\,
            in3 => \N__4931\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Tx_Data_i7_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4895\,
            in1 => \N__5492\,
            in2 => \_gnd_net_\,
            in3 => \N__4919\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Tx_Data_i0_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4838\,
            in1 => \N__4891\,
            in2 => \_gnd_net_\,
            in3 => \N__4907\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Tx_Data_i2_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4893\,
            in1 => \N__4796\,
            in2 => \_gnd_net_\,
            in3 => \N__4865\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_out_i0_i5_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__5705\,
            in1 => \N__4849\,
            in2 => \_gnd_net_\,
            in3 => \N__5870\,
            lcout => data_out_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_out_i0_i0_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4834\,
            in1 => \N__5231\,
            in2 => \_gnd_net_\,
            in3 => \N__5703\,
            lcout => data_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_out_i0_i3_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__5704\,
            in1 => \N__4822\,
            in2 => \_gnd_net_\,
            in3 => \N__5900\,
            lcout => data_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_out_i0_i1_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4807\,
            in1 => \N__5219\,
            in2 => \_gnd_net_\,
            in3 => \N__5700\,
            lcout => data_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_out_i0_i2_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__5701\,
            in1 => \N__4792\,
            in2 => \_gnd_net_\,
            in3 => \N__5915\,
            lcout => data_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5204\,
            in1 => \N__5188\,
            in2 => \N__5177\,
            in3 => \N__5161\,
            lcout => OPEN,
            ltout => \n38_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i21_4_lut_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5006\,
            in1 => \N__5540\,
            in2 => \N__5150\,
            in3 => \N__5498\,
            lcout => n44,
            ltout => \n44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i710_4_lut_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__5599\,
            in1 => \N__5125\,
            in2 => \N__5147\,
            in3 => \N__4945\,
            lcout => \counter_31__N_172\,
            ltout => \counter_31__N_172_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_out_i0_i4_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5137\,
            in2 => \N__5144\,
            in3 => \N__5885\,
            lcout => data_out_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \send_29_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__5600\,
            in1 => \N__5126\,
            in2 => \N__4949\,
            in3 => \N__5105\,
            lcout => \r_SM_Main_2_N_236_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_out_i0_i6_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__5702\,
            in1 => \N__5068\,
            in2 => \_gnd_net_\,
            in3 => \N__5855\,
            lcout => data_out_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5056\,
            in1 => \N__5044\,
            in2 => \N__5033\,
            in3 => \N__5017\,
            lcout => n36,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i17_4_lut_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4999\,
            in1 => \N__4987\,
            in2 => \N__4976\,
            in3 => \N__4960\,
            lcout => n40,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16_4_lut_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5650\,
            in1 => \N__5638\,
            in2 => \N__5627\,
            in3 => \N__5611\,
            lcout => n39,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5590\,
            in1 => \N__5578\,
            in2 => \N__5567\,
            in3 => \N__5551\,
            lcout => n37,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_3_lut_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5533\,
            in1 => \N__5521\,
            in2 => \_gnd_net_\,
            in3 => \N__5509\,
            lcout => n35,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_out_i0_i7_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5836\,
            in1 => \N__5488\,
            in2 => \_gnd_net_\,
            in3 => \N__5706\,
            lcout => data_out_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.r_Bit_Index_i1_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5438\,
            in2 => \_gnd_net_\,
            in3 => \N__5476\,
            lcout => \uart.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5391\,
            ce => \N__5330\,
            sr => \N__5303\
        );

    \integrator_118__i0_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5230\,
            in2 => \N__5275\,
            in3 => \_gnd_net_\,
            lcout => integrator_0,
            ltout => OPEN,
            carryin => \bfn_5_23_0_\,
            carryout => n2188,
            clk => \N__5815\,
            ce => 'H',
            sr => \N__5708\
        );

    \integrator_118__i1_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5218\,
            in2 => \_gnd_net_\,
            in3 => \N__5207\,
            lcout => integrator_1,
            ltout => OPEN,
            carryin => n2188,
            carryout => n2189,
            clk => \N__5815\,
            ce => 'H',
            sr => \N__5708\
        );

    \integrator_118__i2_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5914\,
            in2 => \_gnd_net_\,
            in3 => \N__5903\,
            lcout => integrator_2,
            ltout => OPEN,
            carryin => n2189,
            carryout => n2190,
            clk => \N__5815\,
            ce => 'H',
            sr => \N__5708\
        );

    \integrator_118__i3_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5899\,
            in2 => \_gnd_net_\,
            in3 => \N__5888\,
            lcout => integrator_3,
            ltout => OPEN,
            carryin => n2190,
            carryout => n2191,
            clk => \N__5815\,
            ce => 'H',
            sr => \N__5708\
        );

    \integrator_118__i4_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5884\,
            in2 => \_gnd_net_\,
            in3 => \N__5873\,
            lcout => integrator_4,
            ltout => OPEN,
            carryin => n2191,
            carryout => n2192,
            clk => \N__5815\,
            ce => 'H',
            sr => \N__5708\
        );

    \integrator_118__i5_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5869\,
            in2 => \_gnd_net_\,
            in3 => \N__5858\,
            lcout => integrator_5,
            ltout => OPEN,
            carryin => n2192,
            carryout => n2193,
            clk => \N__5815\,
            ce => 'H',
            sr => \N__5708\
        );

    \integrator_118__i6_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5854\,
            in2 => \_gnd_net_\,
            in3 => \N__5843\,
            lcout => integrator_6,
            ltout => OPEN,
            carryin => n2193,
            carryout => n2194,
            clk => \N__5815\,
            ce => 'H',
            sr => \N__5708\
        );

    \integrator_118__i7_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5837\,
            in2 => \_gnd_net_\,
            in3 => \N__5840\,
            lcout => integrator_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5815\,
            ce => 'H',
            sr => \N__5708\
        );
end \INTERFACE\;
