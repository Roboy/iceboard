// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Sun Sep 22 19:35:58 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    output PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    output PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    output PIN_3 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    output PIN_4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    output PIN_5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    output PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    input PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    input PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    input PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    inout PIN_13 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    inout PIN_14 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    inout PIN_15 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    inout PIN_16 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    input PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    input PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    input PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    input PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    input PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    input PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire GND_net, VCC_net, CLK_c, LED_c, PIN_1_c_5, PIN_2_c_4, PIN_3_c_3, 
        PIN_4_c_2, PIN_5_c_1, PIN_6_c_0, PIN_8_c_1, PIN_9_c_0, PIN_23_c_0, 
        PIN_24_c_1, tx_o, tx_enable, rx_i;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(75[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(76[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(77[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(78[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(79[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(80[22:24])
    
    wire n47641;
    wire [23:0]Kd;   // verilog/TinyFPGA_B.v(81[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(82[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(83[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(84[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(85[22:30])
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(86[22:34])
    
    wire hall1, hall2, hall3;
    wire [23:0]pwm;   // verilog/TinyFPGA_B.v(94[10:13])
    wire [31:0]motor_state;   // verilog/TinyFPGA_B.v(143[22:33])
    wire [31:0]motor_state_23__N_25;
    wire [24:0]displacement_23__N_91;
    wire [23:0]displacement_23__N_1;
    
    wire rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(88[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(92[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(92[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(92[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(92[12:19])
    
    wire n37403;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(94[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(94[12:26])
    
    wire n20156;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(94[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(99[12:33])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(109[11:16])
    
    wire n37402, n249, n248, n37401, n37400, n37399, n37398, n37397, 
        n122, n37396, n47595;
    wire [31:0]\FRAME_MATCHER.state_31__N_1860 ;
    
    wire n37395, n37394, n47576, n47574, n37393, n47566, n47564, 
        n48543, n47554, n47552, n48631, n47548, n47226, n47546, 
        n47542, n47540, n2299, n37392, n2298, n2297, n47532, n37391, 
        n37390, n47530, n37389, n37388, n37387, n37386, n37385, 
        n47524, n48150, n47521, n37384, n37383, n47512, n37382, 
        n37381, n37380, n37379, n37378, n37377, n37376, n47492, 
        n47214, n36941, n37375, n36940, n37374, n37373, n37372, 
        n37371, n737, n37370, n47483, n37369, n47212, n36939, 
        n37368, n37367, n36938, n37366, n37365, n37364, n37363, 
        n37362, n37361, n37360, n37359, n48305, n36937, n36936, 
        n24414, n24413, n24412, n6933, n47203, n37358, n42006, 
        n37357, n37356, n37355, n37354, n22624, n37353, n22621, 
        n47199, n37352, n37351, n37350, n37349, n37348, n37347, 
        n37346, n37345, n37344, n37343, n37342, n36693, n36692, 
        n36691, n36690, n36689, n36688, n36687, n36686, n36685, 
        n36684, n36683, n36682, n36681, n36680, n36679, n22618, 
        n6, n4, n36678, n2, n36677, n36676, n36675, n36674, 
        n22615, n36673, n36672, n22612, n36671, n22609, n22606, 
        n48147, n22603, n22600, n22597, n4_adj_3953, n2243, n2119, 
        n2296, n2295, n2294, n2293, n2266, n2265, n2264, n2263, 
        n2241, n37341, n37340, n2854, n37339, n48489, n37338, 
        n22594, n22591, n22588, n2_adj_3954, n48156, n37337, n22585, 
        n24320, n47323, n47181, n37336, n22582, n22579, n24405, 
        n3758, n37335, n2_adj_3955, n47285, n29023, n47281, n47275, 
        n22576, n47171, n37334, n37333, n37332, n37331, n37330, 
        n37329, n37328, n47167, n37327, n37326, n37325, n37324, 
        n37323, n37322, n37321, n37320, n37319, n37318, n37317, 
        n37316, n37315, n37314, n37313, n37312, n28694, n37311, 
        n37310, n37309, n48505, n37308, n48639, n37307, n37306, 
        n47161, n37305, n37304, n37303, n37302, n37301, n47157, 
        n37300, n37299, n37298, n37297, n37296, n37295, n37294, 
        n37293, n37292, n37291, n37290, n37289, n24319, n37288, 
        n37287, n37286, n37285, n37284, n37283, n37282, n37281, 
        n37280, n37279, n37278, n37277, n37276, n37275, n37274, 
        n37273, n24318, n37272, n37271, n37270, n37269, n37268, 
        n37267, n37266, n37265, n24317, n24316, n24306, n37264, 
        n37263, n47135, n37262, n24158, n224, n6838, n47123, n99, 
        n98, n97, n96, n95, n94, n93, n92, n91, n90, n89, 
        n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, 
        n78, n77, n75, n74, n73, n72, n71, n70, n69, n68, 
        n67, n66, n65, n64, n63, n62, n61, n60, n59, n58, 
        n57, n56, n55, n54, n53, n25, n24, n23, n22, n21, 
        n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, 
        n10, n9, n8, n7, n6_adj_3956, n5, n4_adj_3957, n3, n37261, 
        n37260, n47119, n37259, n37258, n37257, n37256, n28517, 
        n48195, n24407, n37255, n47115, n24403, n37254, n24307, 
        n37253, n47111, n37252, n24404, n37251, n7027, n47939, 
        n7002, n6978, n6955, n37250, n3823, n3822, n3821, n3820, 
        n3819, n3818, n3817, n3816, n3815, n3814, n3813, n3812, 
        n3811, n3810, n3809, n3808, n3807, n3806, n3805, n3804, 
        n3803, n3802, n3801, n3800, n37249, n37248, n37247, n37246, 
        n37245, n37244, n48126, n15_adj_3958, n28989, n15_adj_3959, 
        n37243, n2262, n2261, n2260, n2259, n4016, n2258, n37242, 
        n2257, n47089;
    wire [31:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(23[23:26])
    wire [31:0]\PID_CONTROLLER.err_prev ;   // verilog/motorControl.v(24[23:31])
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(25[23:29])
    wire [8:0]pwm_count;   // verilog/motorControl.v(55[13:22])
    
    wire n48536, n48125, n24315, n25_adj_3960, n24_adj_3961, n23_adj_3962, 
        n22_adj_3963, n21_adj_3964, n20_adj_3965, n19_adj_3966, n18_adj_3967, 
        n17_adj_3968, n16_adj_3969, n15_adj_3970, n14_adj_3971, n13_adj_3972, 
        n12_adj_3973, n11_adj_3974, n10_adj_3975, n9_adj_3976, n8_adj_3977, 
        n7_adj_3978, n6_adj_3979;
    wire [31:0]pwm_23__N_2951;
    
    wire pwm_23__N_2948, n387, n37241, n3840, n413, n415, n416, 
        n421, n37240, n47081, n455, n456, n457, n458, n459, 
        n460, n461, n462, n463, n465, n468, n469, n470, n471, 
        n37239, n4_adj_3980, n48114, n4_adj_3981, n47077, n2256, 
        n37238, n2255, n2254, n2253, n2252, n37237, n2251, n2250, 
        n2249, n37236, n2244, n2245, n37235, n37234, n37233, n24391, 
        n24411, n37232, n37231, n868, n869, n870, n871, n872, 
        n873, n874, n875, n37230, n24408, n37229, n24401, n24402, 
        n37228, n37227, n48637, n2248, quadA_debounced, quadB_debounced, 
        count_enable, n37226, n37225, n37224, n47071, n37223, n37222, 
        n47069, quadA_debounced_adj_3982, quadB_debounced_adj_3983, count_enable_adj_3984, 
        n37221, n37220, n37219, n37218, n46682, n2316, n2315, 
        n2314, n2313, n37217, n4038, n37216, n15_adj_3985, n48199, 
        r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n4_adj_3986, n37215, n37214, n2247, n37213, n24314, n24313, 
        n24312, n37212, n37211, n37210, n2246;
    wire [2:0]r_Bit_Index_adj_4404;   // verilog/uart_tx.v(33[16:27])
    
    wire n37209, n24311, n24310, n24309, n2312, n37208, n2311, 
        n2310, n2309, n37207, n37206, n2308, n2307, n2306, n2305, 
        n2304, n2303, n2302, n37205, n2301, n37204;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    wire [1:0]reg_B_adj_4411;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n37203, n2300, n37202, n37201, n37200, n6912, n37199, 
        n48259, n37198, n37197, n3362, n24406, n37196, n37195, 
        n37194, n37193, n48324, n3_adj_3992, n48545, n369, n370, 
        n371, n372, n373, n374, n375, n376, n377, n378, n379, 
        n380, n381, n382, n383, n384, n385, n386, n387_adj_3993, 
        n388, n389, n390, n391, n392, n393, n47026, n47993, 
        n510, n533, n534, n558, n47013, n648, n649, n671, n672, 
        n47995, n6855, n783, n784, n785, n806, n807, n914, n915, 
        n916, n917, n918, n938, n939, n1043, n1044, n1045, n1046, 
        n1047, n1048, n1067, n1068, n23785, n23783, n1169, n1170, 
        n1171, n1172, n1173, n1174, n1175, n48635, n1193, n1194, 
        n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
        n1316, n1317, n43447, n6873, n1412, n1413, n1414, n1415, 
        n1416, n1417, n1418, n1419, n1420, n1436, n1437, n24308, 
        n46968, n46964, n1529, n1530, n1531, n1532, n1533, n1534, 
        n1535, n1536, n1537, n1538, n1553, n1554, n6743, n6744, 
        n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, 
        n6753, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
        n1650, n1651, n1652, n1653, n1667, n1668, n48271, n1754, 
        n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
        n1763, n1764, n1765, n1778, n1779, n1862, n1863, n1864, 
        n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
        n1873, n1874, n1886, n1887, n46943, n6841, n6842, n6843, 
        n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, 
        n6852, n6853, n6854, n1967, n1968, n1969, n1970, n1971, 
        n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
        n1980, n1991, n1992, n6858, n6859, n6860, n6861, n6862, 
        n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, 
        n6871, n6872, n2069, n2070, n2071, n2072, n2073, n2074, 
        n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
        n2083, n2093, n2094, n46937, n6876, n6877, n6878, n6879, 
        n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, 
        n6888, n6889, n6890, n6891, n2168, n2169, n2170, n2171, 
        n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
        n2180, n2181, n2182, n2183, n5826, n2192, n2193, n6895, 
        n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, 
        n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, 
        n48015, n2264_adj_3994, n2265_adj_3995, n2266_adj_3996, n2267, 
        n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, 
        n2276, n2277, n2278, n2279, n2280, n2288, n2289, n6915, 
        n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
        n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, 
        n6932, n6218, n46927, n2357, n2358, n2359, n2360, n2361, 
        n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
        n2370, n2371, n2372, n2373, n2374, n2381, n2382, n6936, 
        n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, 
        n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, 
        n6953, n6954, n2447, n2448, n2449, n2450, n2451, n2452, 
        n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
        n2461, n2462, n2463, n2464, n2465, n2471, n2472, n48017, 
        n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, 
        n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, 
        n6974, n6975, n6976, n6977, n6579, n2534, n2535, n2536, 
        n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
        n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
        n2553, n43773, n2558, n2559, n43351, n6981, n6982, n6983, 
        n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, 
        n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, 
        n7000, n7001, n5827, n2618, n2619, n2620, n2621, n2622, 
        n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
        n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
        n2642, n2643, n7005, n7006, n7007, n7008, n7009, n7010, 
        n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, 
        n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, 
        n43349, n2699, n2700, n2701, n2702, n2703, n2704, n2705, 
        n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
        n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2723, 
        n2724, n8_adj_3997, n49493, n2777, n2798, n2799, n2801, 
        n2802, n22534, n28227, n23966, n23965, n23964, n23963, 
        n28170, n23962, n23961, n23960, n23959, n6219, n23958, 
        n6580, n48541, n6650, n48640, n5828, n46891, n63_adj_3998, 
        n46887, n46881, n6220, n5_adj_3999, n6581, n6690, n22573, 
        n6651, n5829, n46873, n22513, n6221, n48281, n6582, n6730, 
        n6691, n6652, n5830, n46836, n48389, n47463, n48332, n9_adj_4000, 
        n15_adj_4001, n9_adj_4002, n11_adj_4003, n15_adj_4004, n1, 
        n9_adj_4005, n11_adj_4006, n15_adj_4007, n46829, n9_adj_4008, 
        n11_adj_4009, n15_adj_4010, n44475, n6837, n22525, n22512, 
        n4_adj_4011, n6_adj_4012, n8_adj_4013, n9_adj_4014, n11_adj_4015, 
        n13_adj_4016, n15_adj_4017, n23957, n23956, n23955, n23954, 
        n23953, n23952, n23951, n23950, n39599, n23949, n23948, 
        n23947, n23946, n23945, n23944, n23943, n23941, n23940, 
        n23939, n23938, n23937, n23936, n23935, n23934, n23933, 
        n23932, n23931, n23930, n23929, n23928, n23927, n23926, 
        n23925, n23924, n23923, n23922, n23921, n23920, n23919, 
        n23918, n23915, n23914, n23913, n23909, n23907, n23906, 
        n23904, n23903, n23901, n23900, n23898, n23897, n23895, 
        n23894, n23892, n23891, n23889, n23888, n23887, n23886, 
        n23885, n23884, n23883, n23882, n23881, n23878, n23875, 
        n23872, n23868, n23866, n23865, n23863, n23862, n23860, 
        n23859, n23857, n23856, n37162, n23854, n23853, n23851, 
        n23850, n37161, n23848, n23847, n6892, n46820, n37160, 
        n37159, n37158, n37157, n46808, n37156, n5025, n6222, 
        n48039, n6583, n6784, n6731, n6692, n6653, n5831, n46796, 
        n6223, n22528, n48041, n6584, n6825, n6785, n6732, n46793, 
        n6693, n6654, n6224, n4_adj_4018, n6_adj_4019, n8_adj_4020, 
        n9_adj_4021, n11_adj_4022, n13_adj_4023, n15_adj_4024, n5023, 
        n36777, n36776, n6796, n46787, n6836, n36775, n23845, 
        n36774, n36773, n6585, n6826, n6786, n6733, n6694, n6655, 
        n2_adj_4025, n3_adj_4026, n4_adj_4027, n5_adj_4028, n6_adj_4029, 
        n7_adj_4030, n8_adj_4031, n9_adj_4032, n10_adj_4033, n11_adj_4034, 
        n12_adj_4035, n13_adj_4036, n14_adj_4037, n15_adj_4038, n16_adj_4039, 
        n17_adj_4040, n18_adj_4041, n19_adj_4042, n20_adj_4043, n21_adj_4044, 
        n22_adj_4045, n23_adj_4046, n24_adj_4047, n25_adj_4048, n2_adj_4049, 
        n3_adj_4050, n4_adj_4051, n5_adj_4052, n6_adj_4053, n7_adj_4054, 
        n8_adj_4055, n9_adj_4056, n10_adj_4057, n11_adj_4058, n12_adj_4059, 
        n13_adj_4060, n14_adj_4061, n15_adj_4062, n16_adj_4063, n17_adj_4064, 
        n18_adj_4065, n19_adj_4066, n20_adj_4067, n21_adj_4068, n22_adj_4069, 
        n23_adj_4070, n24_adj_4071, n25_adj_4072, n6586, n6827, n6787, 
        n6734, n6695, n46783, n6656, n8_adj_4073, n6_adj_4074, n46777, 
        n46775, n46773, n4_adj_4075, n6828, n46769, n6788, n6735, 
        n6696, n6657, n46, n46767, n6829, n48289, n6789, n6736, 
        n44, n6697, n46765, n6658, n24482, n24478, n42, n48347, 
        n24477, n24476, n24475, n24474, n24473, n24472, n24471, 
        n24470, n24469, n24468, n24467, n24466, n24465, n24464, 
        n24463, n24462, n24461, n24460, n6830, n6790, n6737, n6698, 
        n24459, n40, n42_adj_4076, n44_adj_4077, n45, n24458, n24457, 
        n24456, n24454, n24453, n24452, n24451, n24450, n24449, 
        n24448, n24447, n24444, n24443, n24442, n38, n40_adj_4078, 
        n42_adj_4079, n43, n47945, n48345, n24441, n24440, n24439, 
        n24438, n24437, n24436, n24434, n24431, n24430, n24426, 
        n2_adj_4080, n6831, n6791, n6738, n6699, n24423, n36, 
        n38_adj_4081, n40_adj_4082, n41, n48393, n24422, n24421, 
        n24420, n24419, n24418, n24417, n24416, n24415, n24304, 
        n23828, n24305, n24303, n46751, n24302, n34, n36_adj_4083, 
        n38_adj_4084, n39, n41_adj_4085, n43_adj_4086, n44_adj_4087, 
        n45_adj_4088, n47947, n24301, n24300, n24298, n23821, n24299, 
        n24297, n24296, n23817, n24295, n6832, n6792, n6739, n23816, 
        n32, n34_adj_4089, n37, n39_adj_4090, n41_adj_4091, n48339, 
        n43_adj_4092, n47949, n48214, n24294, n23815, n24293, n23655, 
        n24292, n24291, n23649, n24290, n30, n31, n32_adj_4093, 
        n33, n34_adj_4094, n35, n37_adj_4095, n39_adj_4096, n48337, 
        n41_adj_4097, n42_adj_4098, n43_adj_4099, n45_adj_4100, n48538, 
        n24289, n23814, n6833, n6793, n28, n29, n30_adj_4101, 
        n31_adj_4102, n32_adj_4103, n33_adj_4104, n35_adj_4105, n37_adj_4106, 
        n48335, n39_adj_4107, n40_adj_4108, n41_adj_4109, n43_adj_4110, 
        n47955, n48333, n48515, n23812, n6740, n26, n27, n28_adj_4111, 
        n29_adj_4112, n30_adj_4113, n31_adj_4114, n33_adj_4115, n35_adj_4116, 
        n48331, n37_adj_4117, n38_adj_4118, n39_adj_4119, n41_adj_4120, 
        n48540, n23616, n24288, n24287, n24_adj_4121, n25_adj_4122, 
        n26_adj_4123, n27_adj_4124, n28_adj_4125, n29_adj_4126, n30_adj_4127, 
        n31_adj_4128, n32_adj_4129, n33_adj_4130, n35_adj_4131, n36_adj_4132, 
        n37_adj_4133, n39_adj_4134, n41_adj_4135, n43_adj_4136, n44_adj_4137, 
        n45_adj_4138, n47957, n22_adj_4139, n23_adj_4140, n24_adj_4141, 
        n25_adj_4142, n26_adj_4143, n27_adj_4144, n28_adj_4145, n29_adj_4146, 
        n30_adj_4147, n31_adj_4148, n33_adj_4149, n34_adj_4150, n35_adj_4151, 
        n37_adj_4152, n39_adj_4153, n41_adj_4154, n42_adj_4155, n43_adj_4156, 
        n48109, n48105, n48323, n6834, n6794, n24284, n23808, 
        n20_adj_4157, n21_adj_4158, n22_adj_4159, n23_adj_4160, n24_adj_4161, 
        n25_adj_4162, n26_adj_4163, n27_adj_4164, n28_adj_4165, n29_adj_4166, 
        n31_adj_4167, n32_adj_4168, n33_adj_4169, n35_adj_4170, n37_adj_4171, 
        n39_adj_4172, n48546, n41_adj_4173, n47965, n48548, n18_adj_4174, 
        n19_adj_4175, n20_adj_4176, n21_adj_4177, n22_adj_4178, n23_adj_4179, 
        n24_adj_4180, n25_adj_4181, n26_adj_4182, n27_adj_4183, n29_adj_4184, 
        n30_adj_4185, n31_adj_4186, n33_adj_4187, n35_adj_4188, n48235, 
        n37_adj_4189, n48638, n39_adj_4190, n41_adj_4191, n47525, 
        n43_adj_4192, n45_adj_4193, n48237, n48517, n16_adj_4194, 
        n17_adj_4195, n18_adj_4196, n19_adj_4197, n20_adj_4198, n21_adj_4199, 
        n22_adj_4200, n23_adj_4201, n25_adj_4202, n27_adj_4203, n28_adj_4204, 
        n29_adj_4205, n31_adj_4206, n33_adj_4207, n35_adj_4208, n37_adj_4209, 
        n39_adj_4210, n41_adj_4211, n43_adj_4212, n48608, n48055, 
        n14_adj_4213, n16_adj_4214, n17_adj_4215, n18_adj_4216, n19_adj_4217, 
        n20_adj_4218, n21_adj_4219, n22_adj_4220, n23_adj_4221, n25_adj_4222, 
        n26_adj_4223, n27_adj_4224, n29_adj_4225, n31_adj_4226, n33_adj_4227, 
        n35_adj_4228, n37_adj_4229, n39_adj_4230, n40_adj_4231, n41_adj_4232, 
        n43_adj_4233, n45_adj_4234, n48519, n12_adj_4235, n14_adj_4236, 
        n15_adj_4237, n16_adj_4238, n17_adj_4239, n18_adj_4240, n19_adj_4241, 
        n20_adj_4242, n21_adj_4243, n23_adj_4244, n24_adj_4245, n25_adj_4246, 
        n27_adj_4247, n29_adj_4248, n48493, n31_adj_4249, n33_adj_4250, 
        n35_adj_4251, n37_adj_4252, n38_adj_4253, n39_adj_4254, n41_adj_4255, 
        n43_adj_4256, n48471, n48641, n6835, n6795, n10_adj_4257, 
        n12_adj_4258, n13_adj_4259, n14_adj_4260, n15_adj_4261, n16_adj_4262, 
        n17_adj_4263, n18_adj_4264, n19_adj_4265, n21_adj_4266, n22_adj_4267, 
        n23_adj_4268, n25_adj_4269, n27_adj_4270, n29_adj_4271, n48129, 
        n31_adj_4272, n33_adj_4273, n35_adj_4274, n36_adj_4275, n37_adj_4276, 
        n39_adj_4277, n41_adj_4278, n48636, n6754, n8_adj_4279, n10_adj_4280, 
        n11_adj_4281, n12_adj_4282, n13_adj_4283, n14_adj_4284, n15_adj_4285, 
        n16_adj_4286, n17_adj_4287, n19_adj_4288, n20_adj_4289, n21_adj_4290, 
        n23_adj_4291, n25_adj_4292, n48120, n27_adj_4293, n29_adj_4294, 
        n31_adj_4295, n33_adj_4296, n34_adj_4297, n35_adj_4298, n37_adj_4299, 
        n39_adj_4300, n48117, n47967, n48633, n6_adj_4301, n8_adj_4302, 
        n9_adj_4303, n10_adj_4304, n11_adj_4305, n12_adj_4306, n13_adj_4307, 
        n14_adj_4308, n15_adj_4309, n17_adj_4310, n19_adj_4311, n21_adj_4312, 
        n23_adj_4313, n48111, n25_adj_4314, n47969, n27_adj_4315, 
        n29_adj_4316, n31_adj_4317, n32_adj_4318, n33_adj_4319, n35_adj_4320, 
        n37_adj_4321, n48313, n48469, n4_adj_4322, n6_adj_4323, n7_adj_4324, 
        n8_adj_4325, n9_adj_4326, n10_adj_4327, n11_adj_4328, n12_adj_4329, 
        n13_adj_4330, n15_adj_4331, n16_adj_4332, n17_adj_4333, n19_adj_4334, 
        n21_adj_4335, n48311, n23_adj_4336, n24_adj_4337, n25_adj_4338, 
        n27_adj_4339, n48309, n29_adj_4340, n30_adj_4341, n31_adj_4342, 
        n33_adj_4343, n35_adj_4344, n37_adj_4345, n48415, n39_adj_4346, 
        n40_adj_4347, n41_adj_4348, n43_adj_4349, n48130, n45_adj_4350, 
        n48417, n48059, n46736, n46730, n48295, n46710, n46706, 
        n37553, n46702, n37552, n37551, n48075, n37550, n46700, 
        n37549, n37548, n37547, n37546, n48079, n37545, n46684, 
        n37544, n37543, n46675, n37542, n46673, n37541, n37540, 
        n37539, n37538, n37537, n37536, n37535, n37534, n37533, 
        n44107, n37532, n37531, n50013, n46661, n46659, n37530, 
        n46657, n37529, n37528, n46655, n37527, n37526, n37525, 
        n37524, n48312, n48316, n37523, n37522, n37521, n37520, 
        n37519, n46641, n37518, n37517, n46639, n37516, n37515, 
        n46637, n37514, n37513, n37512, n22531, n37511, n37510, 
        n37509, n37508, n48310, n46635, n22511, n22633, n22630, 
        n22627, n43347, n22498, n22539, n37441, n37440, n46604, 
        n37439, n37438, n37437, n37436, n37435, n1_adj_4351, n37434, 
        n37433, n24410, n37432, n24409, n37431, n37430, n37429, 
        n37428, n37427, n37426, n48119, n37425, n37424, n37423, 
        n37422, n37421, n37420, n37419, n46996, n37418, n44592, 
        n37417, n37416, n37415, n37414, n37413, n37412, n37411, 
        n37410, n37409, n37408, n24388, n37407, n48121, n37406, 
        n37405, n37404, n46591, n46590, n30_adj_4352, n29_adj_4353, 
        n24_adj_4354, n23_adj_4355, n22_adj_4356, n21_adj_4357, n20_adj_4358, 
        n19_adj_4359, n48131, n18_adj_4360, n17_adj_4361, n46573, 
        n46571, n46569, n46567, n46565, n48143, n48141, n10_adj_4362, 
        n48148, n5_adj_4363, n41480, n48149, n49328, n44154, n48155, 
        n46540, n46539, n48537, n41946, n3_adj_4364, n5_adj_4365, 
        n6_adj_4366, n44066, n48193, n47933, n48629, n48196, n48627, 
        n48625, n48624, n48597, n48626, n48593, n48628, n48594, 
        n48572, n48571, n48606, n48558, n48557, n48610, n48551, 
        n48549, n48547, n48496, n48494, n48492, n48490, n48486, 
        n48482, n48480, n48395, n48478, n48476, n48474, n48470, 
        n47268, n47587, n48427, n48408, n48404, n48544, n48542, 
        n48394, n48118, n48374, n48491, n48371, n48368, n48366, 
        n48495, n48362, n48497, n48499, n48113, n48501, n48348, 
        n48346, n48342, n48340, n48338, n48336, n48250, n48248, 
        n48239, n48220, n48216, n48210, n48341, n48110, n48144, 
        n48136, n48135, n47865, n47841, n47837, n47825, n47789, 
        n47747, n47701, n47687, n44557, n47657;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n2292({n2293, n2294, n2295, 
            n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, 
            n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, 
            n2312, n2313, n2314, n2315, n2316}), .encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .data_o({quadA_debounced, quadB_debounced}), 
            .clk32MHz(clk32MHz), .n23941(n23941), .n23940(n23940), .n23939(n23939), 
            .n23938(n23938), .n23937(n23937), .n23936(n23936), .n23935(n23935), 
            .n23934(n23934), .n23933(n23933), .n23932(n23932), .n23931(n23931), 
            .n23930(n23930), .n23929(n23929), .n23928(n23928), .n23927(n23927), 
            .n23926(n23926), .n23925(n23925), .n23924(n23924), .n23923(n23923), 
            .n23922(n23922), .n23921(n23921), .n23920(n23920), .n23919(n23919), 
            .n23814(n23814), .count_enable(count_enable), .n24423(n24423), 
            .PIN_8_c_1(PIN_8_c_1), .reg_B({reg_B}), .PIN_9_c_0(PIN_9_c_0), 
            .n23816(n23816), .n44475(n44475)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(175[15] 180[4])
    SB_IO rx_input (.PACKAGE_PIN(PIN_13), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), .D_OUT_1(GND_net), 
          .D_OUT_0(GND_net), .D_IN_0(rx_i)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam rx_input.PIN_TYPE = 6'b000001;
    defparam rx_input.PULLUP = 1'b1;
    defparam rx_input.NEG_TRIGGER = 1'b0;
    defparam rx_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(PIN_16), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall2_input (.PACKAGE_PIN(PIN_15), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_14), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    motorControl control (.GND_net(GND_net), .VCC_net(VCC_net), .\PID_CONTROLLER.err[31] (\PID_CONTROLLER.err [31]), 
            .\Kd[1] (Kd[1]), .\Kd[0] (Kd[0]), .\Kd[2] (Kd[2]), .\Kd[3] (Kd[3]), 
            .\deadband[3] (deadband[3]), .\Kd[4] (Kd[4]), .\Kd[5] (Kd[5]), 
            .\Kd[6] (Kd[6]), .\motor_state[23] (motor_state[23]), .\deadband[4] (deadband[4]), 
            .\Kd[7] (Kd[7]), .\motor_state[22] (motor_state[22]), .setpoint({setpoint}), 
            .\motor_state[21] (motor_state[21]), .\motor_state[20] (motor_state[20]), 
            .\Kp[1] (Kp[1]), .\PID_CONTROLLER.err[23] (\PID_CONTROLLER.err [23]), 
            .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), .\motor_state[19] (motor_state[19]), 
            .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\motor_state[18] (motor_state[18]), 
            .\Kp[5] (Kp[5]), .n24454(n24454), .pwm({pwm}), .clk32MHz(clk32MHz), 
            .n24451(n24451), .n24450(n24450), .n24449(n24449), .n24448(n24448), 
            .n24447(n24447), .n41480(n41480), .n24444(n24444), .n24443(n24443), 
            .n24442(n24442), .n24441(n24441), .n24440(n24440), .n24439(n24439), 
            .n24438(n24438), .n24437(n24437), .n24436(n24436), .n24434(n24434), 
            .n24431(n24431), .n24430(n24430), .n24426(n24426), .\Kp[6] (Kp[6]), 
            .\Kp[7] (Kp[7]), .\PID_CONTROLLER.err[14] (\PID_CONTROLLER.err [14]), 
            .\PID_CONTROLLER.err[15] (\PID_CONTROLLER.err [15]), .\deadband[5] (deadband[5]), 
            .\PID_CONTROLLER.err[21] (\PID_CONTROLLER.err [21]), .\PID_CONTROLLER.err[22] (\PID_CONTROLLER.err [22]), 
            .\motor_state[17] (motor_state[17]), .\motor_state[16] (motor_state[16]), 
            .\motor_state[15] (motor_state[15]), .\motor_state[14] (motor_state[14]), 
            .\motor_state[13] (motor_state[13]), .\Ki[1] (Ki[1]), .\PID_CONTROLLER.err[0] (\PID_CONTROLLER.err [0]), 
            .\motor_state[12] (motor_state[12]), .\Ki[0] (Ki[0]), .\motor_state[11] (motor_state[11]), 
            .\motor_state[10] (motor_state[10]), .\Ki[2] (Ki[2]), .\motor_state[9] (motor_state[9]), 
            .\Ki[3] (Ki[3]), .\motor_state[8] (motor_state[8]), .\Ki[4] (Ki[4]), 
            .\motor_state[7] (motor_state[7]), .\PWMLimit[2] (PWMLimit[2]), 
            .\motor_state[6] (motor_state[6]), .\motor_state[5] (motor_state[5]), 
            .\motor_state[4] (motor_state[4]), .\Ki[5] (Ki[5]), .\motor_state[3] (motor_state[3]), 
            .\pwm_23__N_2951[7] (pwm_23__N_2951[7]), .\Ki[6] (Ki[6]), .\motor_state[2] (motor_state[2]), 
            .\motor_state[1] (motor_state[1]), .\Ki[7] (Ki[7]), .\pwm_23__N_2951[5] (pwm_23__N_2951[5]), 
            .\motor_state[0] (motor_state[0]), .\pwm_23__N_2951[4] (pwm_23__N_2951[4]), 
            .\deadband[6] (deadband[6]), .\PID_CONTROLLER.err_prev[31] (\PID_CONTROLLER.err_prev [31]), 
            .\deadband[7] (deadband[7]), .\PID_CONTROLLER.err_prev[23] (\PID_CONTROLLER.err_prev [23]), 
            .\PID_CONTROLLER.err_prev[22] (\PID_CONTROLLER.err_prev [22]), 
            .\PID_CONTROLLER.err_prev[21] (\PID_CONTROLLER.err_prev [21]), 
            .\PID_CONTROLLER.err_prev[20] (\PID_CONTROLLER.err_prev [20]), 
            .\PWMLimit[3] (PWMLimit[3]), .\deadband[8] (deadband[8]), .\PID_CONTROLLER.err_prev[19] (\PID_CONTROLLER.err_prev [19]), 
            .\PID_CONTROLLER.err_prev[18] (\PID_CONTROLLER.err_prev [18]), 
            .\PID_CONTROLLER.err_prev[17] (\PID_CONTROLLER.err_prev [17]), 
            .\PID_CONTROLLER.err_prev[16] (\PID_CONTROLLER.err_prev [16]), 
            .\PID_CONTROLLER.err_prev[15] (\PID_CONTROLLER.err_prev [15]), 
            .\PID_CONTROLLER.err_prev[14] (\PID_CONTROLLER.err_prev [14]), 
            .\PID_CONTROLLER.err_prev[13] (\PID_CONTROLLER.err_prev [13]), 
            .\PID_CONTROLLER.err_prev[12] (\PID_CONTROLLER.err_prev [12]), 
            .\PID_CONTROLLER.err_prev[11] (\PID_CONTROLLER.err_prev [11]), 
            .\PID_CONTROLLER.err_prev[10] (\PID_CONTROLLER.err_prev [10]), 
            .\PID_CONTROLLER.err_prev[9] (\PID_CONTROLLER.err_prev [9]), .\deadband[9] (deadband[9]), 
            .\PID_CONTROLLER.err_prev[8] (\PID_CONTROLLER.err_prev [8]), .\PID_CONTROLLER.err_prev[7] (\PID_CONTROLLER.err_prev [7]), 
            .\PID_CONTROLLER.err_prev[6] (\PID_CONTROLLER.err_prev [6]), .\PID_CONTROLLER.err_prev[5] (\PID_CONTROLLER.err_prev [5]), 
            .\PID_CONTROLLER.err_prev[4] (\PID_CONTROLLER.err_prev [4]), .\PID_CONTROLLER.err_prev[3] (\PID_CONTROLLER.err_prev [3]), 
            .\PID_CONTROLLER.err_prev[2] (\PID_CONTROLLER.err_prev [2]), .\PID_CONTROLLER.err_prev[1] (\PID_CONTROLLER.err_prev [1]), 
            .\PID_CONTROLLER.err_prev[0] (\PID_CONTROLLER.err_prev [0]), .n22(n22_adj_4356), 
            .n21(n21_adj_4357), .n24(n24_adj_4354), .n20(n20_adj_4358), 
            .n23(n23_adj_4355), .n19(n19_adj_4359), .\PID_CONTROLLER.err[10] (\PID_CONTROLLER.err [10]), 
            .\PID_CONTROLLER.err[11] (\PID_CONTROLLER.err [11]), .IntegralLimit({IntegralLimit}), 
            .n17(n17_adj_4361), .n48196(n48196), .n18(n18_adj_4360), .n868(n868), 
            .n869(n869), .n870(n870), .n871(n871), .n872(n872), .n873(n873), 
            .n874(n874), .n875(n875), .n46539(n46539), .\PID_CONTROLLER.err[9] (\PID_CONTROLLER.err [9]), 
            .\PID_CONTROLLER.err[8] (\PID_CONTROLLER.err [8]), .\PID_CONTROLLER.err[7] (\PID_CONTROLLER.err [7]), 
            .\PID_CONTROLLER.err[6] (\PID_CONTROLLER.err [6]), .\PID_CONTROLLER.err[5] (\PID_CONTROLLER.err [5]), 
            .\PID_CONTROLLER.err[4] (\PID_CONTROLLER.err [4]), .\PID_CONTROLLER.err[3] (\PID_CONTROLLER.err [3]), 
            .\PID_CONTROLLER.err[2] (\PID_CONTROLLER.err [2]), .\PID_CONTROLLER.err[1] (\PID_CONTROLLER.err [1]), 
            .\pwm_count[8] (pwm_count[8]), .\pwm_count[7] (pwm_count[7]), 
            .\pwm_count[6] (pwm_count[6]), .\pwm_count[5] (pwm_count[5]), 
            .\pwm_count[4] (pwm_count[4]), .\pwm_count[3] (pwm_count[3]), 
            .\pwm_count[2] (pwm_count[2]), .\pwm_count[1] (pwm_count[1]), 
            .n23966(n23966), .n23965(n23965), .n23964(n23964), .n23963(n23963), 
            .n23962(n23962), .n23961(n23961), .n23960(n23960), .n23959(n23959), 
            .n23958(n23958), .n23957(n23957), .n23956(n23956), .n23955(n23955), 
            .n23954(n23954), .n23953(n23953), .n23952(n23952), .n23951(n23951), 
            .n23950(n23950), .n23949(n23949), .n23948(n23948), .n23947(n23947), 
            .n23946(n23946), .n23945(n23945), .n23944(n23944), .n23943(n23943), 
            .\PID_CONTROLLER.result[4] (\PID_CONTROLLER.result [4]), .\PID_CONTROLLER.result[5] (\PID_CONTROLLER.result [5]), 
            .\PID_CONTROLLER.result[7] (\PID_CONTROLLER.result [7]), .PIN_6_c_0(PIN_6_c_0), 
            .PIN_5_c_1(PIN_5_c_1), .PIN_4_c_2(PIN_4_c_2), .PIN_3_c_3(PIN_3_c_3), 
            .PIN_2_c_4(PIN_2_c_4), .\PID_CONTROLLER.err[12] (\PID_CONTROLLER.err [12]), 
            .\PID_CONTROLLER.err[13] (\PID_CONTROLLER.err [13]), .\PID_CONTROLLER.err[16] (\PID_CONTROLLER.err [16]), 
            .\PID_CONTROLLER.err[17] (\PID_CONTROLLER.err [17]), .\PID_CONTROLLER.err[18] (\PID_CONTROLLER.err [18]), 
            .\PID_CONTROLLER.err[19] (\PID_CONTROLLER.err [19]), .\PID_CONTROLLER.err[20] (\PID_CONTROLLER.err [20]), 
            .hall3(hall3), .PIN_1_c_5(PIN_1_c_5), .n413(n413), .n415(n415), 
            .n23812(n23812), .n416(n416), .n421(n421), .n470(n470), 
            .n469(n469), .n468(n468), .pwm_23__N_2948(pwm_23__N_2948), 
            .n28170(n28170), .\PWMLimit[4] (PWMLimit[4]), .n387(n387), 
            .n28227(n28227), .\PWMLimit[5] (PWMLimit[5]), .n465(n465), 
            .n1(n1), .\PWMLimit[7] (PWMLimit[7]), .n463(n463), .n462(n462), 
            .n461(n461), .n460(n460), .n459(n459), .n458(n458), .n457(n457), 
            .n456(n456), .n455(n455), .\PWMLimit[9] (PWMLimit[9]), .n9(n9_adj_4000), 
            .n15(n15_adj_4001), .\deadband[2] (deadband[2]), .\deadband[0] (deadband[0]), 
            .\deadband[1] (deadband[1]), .\PWMLimit[6] (PWMLimit[6]), .n11(n11_adj_4006), 
            .n9_adj_10(n9_adj_4005), .n15_adj_11(n15_adj_4007), .\PWMLimit[8] (PWMLimit[8]), 
            .n11_adj_12(n11_adj_4003), .n9_adj_13(n9_adj_4002), .n15_adj_14(n15_adj_4004), 
            .n11_adj_15(n11_adj_4009), .n9_adj_16(n9_adj_4008), .n15_adj_17(n15_adj_4010), 
            .n471(n471), .\PWMLimit[0] (PWMLimit[0]), .\PWMLimit[1] (PWMLimit[1]), 
            .hall2(hall2), .hall1(hall1), .n29(n29_adj_4353), .n30(n30_adj_4352), 
            .n48193(n48193), .n46604(n46604), .n46565(n46565), .n46567(n46567), 
            .n46573(n46573), .n46571(n46571), .n46569(n46569), .n44066(n44066), 
            .n4(n4_adj_4011)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(152[16] 168[4])
    SB_IO PIN_5_pad (.PACKAGE_PIN(PIN_5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_5_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_5_pad.PIN_TYPE = 6'b011001;
    defparam PIN_5_pad.PULLUP = 1'b0;
    defparam PIN_5_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n36690), .I0(displacement_23__N_91[20]), 
            .I1(n3_adj_3992), .CO(n36691));
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_91[19]), 
            .I2(n6_adj_3979), .I3(n36689), .O(displacement_23__N_1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3033_25_lut (.I0(n249), .I1(n49328), .I2(n248), .I3(n37441), 
            .O(displacement_23__N_91[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3033_24_lut (.I0(n393), .I1(n49328), .I2(n392), .I3(n37440), 
            .O(displacement_23__N_91[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n36689), .I0(displacement_23__N_91[19]), 
            .I1(n6_adj_3979), .CO(n36690));
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_91[18]), 
            .I2(n7_adj_3978), .I3(n36688), .O(displacement_23__N_1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n36688), .I0(displacement_23__N_91[18]), 
            .I1(n7_adj_3978), .CO(n36689));
    SB_CARRY add_3033_24 (.CI(n37440), .I0(n49328), .I1(n392), .CO(n37441));
    SB_LUT4 add_3033_23_lut (.I0(n534), .I1(n49328), .I2(n533), .I3(n37439), 
            .O(displacement_23__N_91[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_91[17]), 
            .I2(n8_adj_3977), .I3(n36687), .O(displacement_23__N_1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3033_23 (.CI(n37439), .I0(n49328), .I1(n533), .CO(n37440));
    SB_LUT4 add_3033_22_lut (.I0(n672), .I1(n49328), .I2(n671), .I3(n37438), 
            .O(displacement_23__N_91[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n36687), .I0(displacement_23__N_91[17]), 
            .I1(n8_adj_3977), .CO(n36688));
    SB_CARRY add_3033_22 (.CI(n37438), .I0(n49328), .I1(n671), .CO(n37439));
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_91[16]), 
            .I2(n9_adj_3976), .I3(n36686), .O(displacement_23__N_1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n36686), .I0(displacement_23__N_91[16]), 
            .I1(n9_adj_3976), .CO(n36687));
    SB_LUT4 add_3033_21_lut (.I0(n807), .I1(n49328), .I2(n806), .I3(n37437), 
            .O(displacement_23__N_91[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_91[15]), 
            .I2(n10_adj_3975), .I3(n36685), .O(displacement_23__N_1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n36685), .I0(displacement_23__N_91[15]), 
            .I1(n10_adj_3975), .CO(n36686));
    SB_CARRY add_3033_21 (.CI(n37437), .I0(n49328), .I1(n806), .CO(n37438));
    SB_LUT4 add_3033_20_lut (.I0(n939), .I1(n49328), .I2(n938), .I3(n37436), 
            .O(displacement_23__N_91[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_20 (.CI(n37436), .I0(n49328), .I1(n938), .CO(n37437));
    SB_LUT4 add_3033_19_lut (.I0(n1068), .I1(n49328), .I2(n1067), .I3(n37435), 
            .O(displacement_23__N_91[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_91[14]), 
            .I2(n11_adj_3974), .I3(n36684), .O(displacement_23__N_1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3033_19 (.CI(n37435), .I0(n49328), .I1(n1067), .CO(n37436));
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n36684), .I0(displacement_23__N_91[14]), 
            .I1(n11_adj_3974), .CO(n36685));
    SB_LUT4 add_3033_18_lut (.I0(n1194), .I1(n49328), .I2(n1193), .I3(n37434), 
            .O(displacement_23__N_91[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_91[13]), 
            .I2(n12_adj_3973), .I3(n36683), .O(displacement_23__N_1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n36683), .I0(displacement_23__N_91[13]), 
            .I1(n12_adj_3973), .CO(n36684));
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_91[12]), 
            .I2(n13_adj_3972), .I3(n36682), .O(displacement_23__N_1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4298));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3033_18 (.CI(n37434), .I0(n49328), .I1(n1193), .CO(n37435));
    SB_LUT4 add_3033_17_lut (.I0(n1317), .I1(n49328), .I2(n1316), .I3(n37433), 
            .O(displacement_23__N_91[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n36682), .I0(displacement_23__N_91[12]), 
            .I1(n13_adj_3972), .CO(n36683));
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_91[11]), 
            .I2(n14_adj_3971), .I3(n36681), .O(displacement_23__N_1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3033_17 (.CI(n37433), .I0(n49328), .I1(n1316), .CO(n37434));
    SB_LUT4 add_3033_16_lut (.I0(n1437), .I1(n49328), .I2(n1436), .I3(n37432), 
            .O(displacement_23__N_91[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n36681), .I0(displacement_23__N_91[11]), 
            .I1(n14_adj_3971), .CO(n36682));
    SB_CARRY add_3033_16 (.CI(n37432), .I0(n49328), .I1(n1436), .CO(n37433));
    SB_LUT4 add_3033_15_lut (.I0(n1554), .I1(n49328), .I2(n1553), .I3(n37431), 
            .O(displacement_23__N_91[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_15 (.CI(n37431), .I0(n49328), .I1(n1553), .CO(n37432));
    SB_LUT4 add_3033_14_lut (.I0(n1668), .I1(n49328), .I2(n1667), .I3(n37430), 
            .O(displacement_23__N_91[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_14 (.CI(n37430), .I0(n49328), .I1(n1667), .CO(n37431));
    SB_LUT4 add_3033_13_lut (.I0(n1779), .I1(n49328), .I2(n1778), .I3(n37429), 
            .O(displacement_23__N_91[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_13 (.CI(n37429), .I0(n49328), .I1(n1778), .CO(n37430));
    SB_LUT4 add_3033_12_lut (.I0(n1887), .I1(n49328), .I2(n1886), .I3(n37428), 
            .O(displacement_23__N_91[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_12 (.CI(n37428), .I0(n49328), .I1(n1886), .CO(n37429));
    SB_LUT4 add_3033_11_lut (.I0(n1992), .I1(n49328), .I2(n1991), .I3(n37427), 
            .O(displacement_23__N_91[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_11 (.CI(n37427), .I0(n49328), .I1(n1991), .CO(n37428));
    SB_LUT4 div_12_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4300));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3033_10_lut (.I0(n2094), .I1(n49328), .I2(n2093), .I3(n37426), 
            .O(displacement_23__N_91[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_10 (.CI(n37426), .I0(n49328), .I1(n2093), .CO(n37427));
    SB_LUT4 add_3033_9_lut (.I0(n2193), .I1(n49328), .I2(n2192), .I3(n37425), 
            .O(displacement_23__N_91[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_9 (.CI(n37425), .I0(n49328), .I1(n2192), .CO(n37426));
    SB_LUT4 add_3033_8_lut (.I0(n2289), .I1(n49328), .I2(n2288), .I3(n37424), 
            .O(displacement_23__N_91[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_8 (.CI(n37424), .I0(n49328), .I1(n2288), .CO(n37425));
    SB_LUT4 add_3033_7_lut (.I0(n2382), .I1(n49328), .I2(n2381), .I3(n37423), 
            .O(displacement_23__N_91[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_7 (.CI(n37423), .I0(n49328), .I1(n2381), .CO(n37424));
    SB_LUT4 div_12_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4296));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3033_6_lut (.I0(n2472), .I1(n49328), .I2(n2471), .I3(n37422), 
            .O(displacement_23__N_91[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_6 (.CI(n37422), .I0(n49328), .I1(n2471), .CO(n37423));
    SB_LUT4 add_3033_5_lut (.I0(n2559), .I1(n49328), .I2(n2558), .I3(n37421), 
            .O(displacement_23__N_91[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_5 (.CI(n37421), .I0(n49328), .I1(n2558), .CO(n37422));
    SB_LUT4 add_3033_4_lut (.I0(n2643), .I1(n49328), .I2(n2642), .I3(n37420), 
            .O(displacement_23__N_91[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_4 (.CI(n37420), .I0(n49328), .I1(n2642), .CO(n37421));
    SB_LUT4 add_3033_3_lut (.I0(n2724), .I1(n49328), .I2(n2723), .I3(n37419), 
            .O(displacement_23__N_91[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_3 (.CI(n37419), .I0(n49328), .I1(n2723), .CO(n37420));
    SB_LUT4 add_3033_2_lut (.I0(n2802), .I1(n49328), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_91[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_2 (.CI(VCC_net), .I0(n49328), .I1(n2801), .CO(n37419));
    SB_LUT4 add_3032_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n37418), 
            .O(n7005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n37417), 
            .O(n7006)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_91[10]), 
            .I2(n15_adj_3970), .I3(n36680), .O(displacement_23__N_1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_24 (.CI(n37417), .I0(n2700), .I1(n79), .CO(n37418));
    SB_LUT4 add_3032_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n37416), 
            .O(n7007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_23 (.CI(n37416), .I0(n2701), .I1(n80), .CO(n37417));
    SB_LUT4 add_3032_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n37415), 
            .O(n7008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_22 (.CI(n37415), .I0(n2702), .I1(n81), .CO(n37416));
    SB_LUT4 add_3032_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n37414), 
            .O(n7009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_21 (.CI(n37414), .I0(n2703), .I1(n82), .CO(n37415));
    SB_LUT4 add_3032_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n37413), 
            .O(n7010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_20 (.CI(n37413), .I0(n2704), .I1(n83), .CO(n37414));
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n36680), .I0(displacement_23__N_91[10]), 
            .I1(n15_adj_3970), .CO(n36681));
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_91[9]), 
            .I2(n16_adj_3969), .I3(n36679), .O(displacement_23__N_1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n37412), 
            .O(n7011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_19 (.CI(n37412), .I0(n2705), .I1(n84), .CO(n37413));
    SB_LUT4 add_3032_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n37411), 
            .O(n7012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_18 (.CI(n37411), .I0(n2706), .I1(n85), .CO(n37412));
    SB_LUT4 add_3032_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n37410), 
            .O(n7013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_17 (.CI(n37410), .I0(n2707), .I1(n86), .CO(n37411));
    SB_LUT4 add_3032_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n37409), 
            .O(n7014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_16 (.CI(n37409), .I0(n2708), .I1(n87), .CO(n37410));
    SB_LUT4 add_3032_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n37408), 
            .O(n7015)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n36679), .I0(displacement_23__N_91[9]), 
            .I1(n16_adj_3969), .CO(n36680));
    SB_CARRY add_3032_15 (.CI(n37408), .I0(n2709), .I1(n88), .CO(n37409));
    SB_LUT4 add_3032_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n37407), 
            .O(n7016)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_14 (.CI(n37407), .I0(n2710), .I1(n89), .CO(n37408));
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_91[8]), 
            .I2(n17_adj_3968), .I3(n36678), .O(displacement_23__N_1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n37406), 
            .O(n7017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_13 (.CI(n37406), .I0(n2711), .I1(n90), .CO(n37407));
    SB_LUT4 add_3032_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n37405), 
            .O(n7018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_12 (.CI(n37405), .I0(n2712), .I1(n91), .CO(n37406));
    SB_LUT4 add_3032_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n37404), 
            .O(n7019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_11 (.CI(n37404), .I0(n2713), .I1(n92), .CO(n37405));
    SB_LUT4 add_3032_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n37403), 
            .O(n7020)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_10 (.CI(n37403), .I0(n2714), .I1(n93), .CO(n37404));
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n36678), .I0(displacement_23__N_91[8]), 
            .I1(n17_adj_3968), .CO(n36679));
    SB_LUT4 add_3032_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n37402), 
            .O(n7021)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_9 (.CI(n37402), .I0(n2715), .I1(n94), .CO(n37403));
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_91[7]), 
            .I2(n18_adj_3967), .I3(n36677), .O(displacement_23__N_1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n37401), 
            .O(n7022)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_8 (.CI(n37401), .I0(n2716), .I1(n95), .CO(n37402));
    SB_LUT4 add_3032_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n37400), 
            .O(n7023)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_7 (.CI(n37400), .I0(n2717), .I1(n96), .CO(n37401));
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n36677), .I0(displacement_23__N_91[7]), 
            .I1(n18_adj_3967), .CO(n36678));
    SB_LUT4 add_3032_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n37399), 
            .O(n7024)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_6 (.CI(n37399), .I0(n2718), .I1(n97), .CO(n37400));
    SB_LUT4 add_3032_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n37398), 
            .O(n7025)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_5 (.CI(n37398), .I0(n2719), .I1(n98), .CO(n37399));
    SB_LUT4 add_3032_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n37397), 
            .O(n7026)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_4 (.CI(n37397), .I0(n2720), .I1(n99), .CO(n37398));
    SB_LUT4 add_3032_3_lut (.I0(GND_net), .I1(n390), .I2(n558), .I3(n37396), 
            .O(n7027)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_3 (.CI(n37396), .I0(n390), .I1(n558), .CO(n37397));
    SB_CARRY add_3032_2 (.CI(VCC_net), .I0(n391), .I1(VCC_net), .CO(n37396));
    SB_LUT4 add_3031_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n37395), 
            .O(n6981)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3031_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n37394), 
            .O(n6982)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_22 (.CI(n37394), .I0(n2619), .I1(n80), .CO(n37395));
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_91[6]), 
            .I2(n19_adj_3966), .I3(n36676), .O(displacement_23__N_1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3031_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n37393), 
            .O(n6983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_21 (.CI(n37393), .I0(n2620), .I1(n81), .CO(n37394));
    SB_LUT4 add_3031_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n37392), 
            .O(n6984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_20 (.CI(n37392), .I0(n2621), .I1(n82), .CO(n37393));
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n36676), .I0(displacement_23__N_91[6]), 
            .I1(n19_adj_3966), .CO(n36677));
    SB_LUT4 div_12_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n389));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3031_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n37391), 
            .O(n6985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_19 (.CI(n37391), .I0(n2622), .I1(n83), .CO(n37392));
    SB_LUT4 add_3031_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n37390), 
            .O(n6986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_18 (.CI(n37390), .I0(n2623), .I1(n84), .CO(n37391));
    SB_LUT4 add_3031_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n37389), 
            .O(n6987)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_17 (.CI(n37389), .I0(n2624), .I1(n85), .CO(n37390));
    SB_LUT4 add_3031_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n37388), 
            .O(n6988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_16 (.CI(n37388), .I0(n2625), .I1(n86), .CO(n37389));
    SB_LUT4 add_3031_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n37387), 
            .O(n6989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_15 (.CI(n37387), .I0(n2626), .I1(n87), .CO(n37388));
    SB_LUT4 add_3031_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n37386), 
            .O(n6990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_14 (.CI(n37386), .I0(n2627), .I1(n88), .CO(n37387));
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_91[5]), 
            .I2(n20_adj_3965), .I3(n36675), .O(displacement_23__N_1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3031_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n37385), 
            .O(n6991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_13 (.CI(n37385), .I0(n2628), .I1(n89), .CO(n37386));
    SB_LUT4 add_3031_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n37384), 
            .O(n6992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_12 (.CI(n37384), .I0(n2629), .I1(n90), .CO(n37385));
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n36675), .I0(displacement_23__N_91[5]), 
            .I1(n20_adj_3965), .CO(n36676));
    SB_LUT4 div_12_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4299));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3031_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n37383), 
            .O(n6993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_11 (.CI(n37383), .I0(n2630), .I1(n91), .CO(n37384));
    SB_LUT4 add_3031_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n37382), 
            .O(n6994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_10 (.CI(n37382), .I0(n2631), .I1(n92), .CO(n37383));
    SB_LUT4 add_3031_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n37381), 
            .O(n6995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_9 (.CI(n37381), .I0(n2632), .I1(n93), .CO(n37382));
    SB_LUT4 add_3031_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n37380), 
            .O(n6996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_8 (.CI(n37380), .I0(n2633), .I1(n94), .CO(n37381));
    SB_LUT4 add_3031_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n37379), 
            .O(n6997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_7 (.CI(n37379), .I0(n2634), .I1(n95), .CO(n37380));
    SB_LUT4 add_3031_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n37378), 
            .O(n6998)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_6 (.CI(n37378), .I0(n2635), .I1(n96), .CO(n37379));
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_91[4]), 
            .I2(n21_adj_3964), .I3(n36674), .O(displacement_23__N_1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3031_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n37377), 
            .O(n6999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_5 (.CI(n37377), .I0(n2636), .I1(n97), .CO(n37378));
    SB_LUT4 add_3031_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n37376), 
            .O(n7000)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_4 (.CI(n37376), .I0(n2637), .I1(n98), .CO(n37377));
    SB_LUT4 add_3031_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n37375), 
            .O(n7001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n36674), .I0(displacement_23__N_91[4]), 
            .I1(n21_adj_3964), .CO(n36675));
    SB_LUT4 div_12_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4293));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3031_3 (.CI(n37375), .I0(n2638), .I1(n99), .CO(n37376));
    SB_LUT4 add_3031_2_lut (.I0(GND_net), .I1(n389), .I2(n558), .I3(VCC_net), 
            .O(n7002)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_2 (.CI(VCC_net), .I0(n389), .I1(n558), .CO(n37375));
    SB_LUT4 add_3030_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n37374), 
            .O(n6958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3030_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n37373), 
            .O(n6959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4294));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3030_21 (.CI(n37373), .I0(n2535), .I1(n81), .CO(n37374));
    SB_LUT4 add_3030_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n37372), 
            .O(n6960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_20 (.CI(n37372), .I0(n2536), .I1(n82), .CO(n37373));
    SB_LUT4 add_3030_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n37371), 
            .O(n6961)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_19 (.CI(n37371), .I0(n2537), .I1(n83), .CO(n37372));
    SB_LUT4 add_3030_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n37370), 
            .O(n6962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_18 (.CI(n37370), .I0(n2538), .I1(n84), .CO(n37371));
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_91[3]), 
            .I2(n22_adj_3963), .I3(n36673), .O(displacement_23__N_1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3030_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n37369), 
            .O(n6963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_17 (.CI(n37369), .I0(n2539), .I1(n85), .CO(n37370));
    SB_LUT4 add_3030_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n37368), 
            .O(n6964)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_16 (.CI(n37368), .I0(n2540), .I1(n86), .CO(n37369));
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n36673), .I0(displacement_23__N_91[3]), 
            .I1(n22_adj_3963), .CO(n36674));
    SB_LUT4 add_3030_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n37367), 
            .O(n6965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_15 (.CI(n37367), .I0(n2541), .I1(n87), .CO(n37368));
    SB_LUT4 add_3030_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n37366), 
            .O(n6966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_14 (.CI(n37366), .I0(n2542), .I1(n88), .CO(n37367));
    SB_LUT4 add_3030_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n37365), 
            .O(n6967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_13 (.CI(n37365), .I0(n2543), .I1(n89), .CO(n37366));
    SB_LUT4 add_3030_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n37364), 
            .O(n6968)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4281));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3030_12 (.CI(n37364), .I0(n2544), .I1(n90), .CO(n37365));
    SB_LUT4 add_3030_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n37363), 
            .O(n6969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_11 (.CI(n37363), .I0(n2545), .I1(n91), .CO(n37364));
    SB_LUT4 add_3030_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n37362), 
            .O(n6970)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_10 (.CI(n37362), .I0(n2546), .I1(n92), .CO(n37363));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_91[2]), 
            .I2(n23_adj_3962), .I3(n36672), .O(displacement_23__N_1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3030_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n37361), 
            .O(n6971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_9 (.CI(n37361), .I0(n2547), .I1(n93), .CO(n37362));
    SB_LUT4 add_3030_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n37360), 
            .O(n6972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_8 (.CI(n37360), .I0(n2548), .I1(n94), .CO(n37361));
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n36672), .I0(displacement_23__N_91[2]), 
            .I1(n23_adj_3962), .CO(n36673));
    SB_LUT4 div_12_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4291));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3030_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n37359), 
            .O(n6973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_7 (.CI(n37359), .I0(n2549), .I1(n95), .CO(n37360));
    SB_LUT4 add_3030_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n37358), 
            .O(n6974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_6 (.CI(n37358), .I0(n2550), .I1(n96), .CO(n37359));
    SB_LUT4 add_3030_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n37357), 
            .O(n6975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_5 (.CI(n37357), .I0(n2551), .I1(n97), .CO(n37358));
    SB_LUT4 add_3030_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n37356), 
            .O(n6976)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_4 (.CI(n37356), .I0(n2552), .I1(n98), .CO(n37357));
    SB_LUT4 div_12_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4292));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3030_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n37355), 
            .O(n6977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_3 (.CI(n37355), .I0(n2553), .I1(n99), .CO(n37356));
    SB_LUT4 add_3030_2_lut (.I0(GND_net), .I1(n388), .I2(n558), .I3(VCC_net), 
            .O(n6978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_91[1]), 
            .I2(n24_adj_3961), .I3(n36671), .O(displacement_23__N_1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_2 (.CI(VCC_net), .I0(n388), .I1(n558), .CO(n37355));
    SB_LUT4 add_3029_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n37354), 
            .O(n6936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3029_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n37353), 
            .O(n6937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_20 (.CI(n37353), .I0(n2448), .I1(n82), .CO(n37354));
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n36671), .I0(displacement_23__N_91[1]), 
            .I1(n24_adj_3961), .CO(n36672));
    SB_LUT4 add_3029_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n37352), 
            .O(n6938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4283));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3029_19 (.CI(n37352), .I0(n2449), .I1(n83), .CO(n37353));
    SB_LUT4 add_3029_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n37351), 
            .O(n6939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_18 (.CI(n37351), .I0(n2450), .I1(n84), .CO(n37352));
    SB_LUT4 add_3029_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n37350), 
            .O(n6940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_17 (.CI(n37350), .I0(n2451), .I1(n85), .CO(n37351));
    SB_LUT4 add_3029_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n37349), 
            .O(n6941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_16 (.CI(n37349), .I0(n2452), .I1(n86), .CO(n37350));
    SB_LUT4 add_3029_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n37348), 
            .O(n6942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_15 (.CI(n37348), .I0(n2453), .I1(n87), .CO(n37349));
    SB_LUT4 add_3029_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n37347), 
            .O(n6943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_14 (.CI(n37347), .I0(n2454), .I1(n88), .CO(n37348));
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_91[0]), 
            .I2(n25_adj_3960), .I3(VCC_net), .O(displacement_23__N_1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3029_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n37346), 
            .O(n6944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_13 (.CI(n37346), .I0(n2455), .I1(n89), .CO(n37347));
    SB_LUT4 add_3029_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n37345), 
            .O(n6945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_12 (.CI(n37345), .I0(n2456), .I1(n90), .CO(n37346));
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_91[0]), 
            .I1(n25_adj_3960), .CO(n36671));
    SB_LUT4 add_3029_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n37344), 
            .O(n6946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_11 (.CI(n37344), .I0(n2457), .I1(n91), .CO(n37345));
    SB_LUT4 add_3029_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n37343), 
            .O(n6947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_10 (.CI(n37343), .I0(n2458), .I1(n92), .CO(n37344));
    SB_LUT4 add_3029_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n37342), 
            .O(n6948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_9 (.CI(n37342), .I0(n2459), .I1(n93), .CO(n37343));
    SB_LUT4 add_3029_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n37341), 
            .O(n6949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_8 (.CI(n37341), .I0(n2460), .I1(n94), .CO(n37342));
    SB_LUT4 add_3029_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n37340), 
            .O(n6950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_7 (.CI(n37340), .I0(n2461), .I1(n95), .CO(n37341));
    SB_LUT4 add_3029_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n37339), 
            .O(n6951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_6 (.CI(n37339), .I0(n2462), .I1(n96), .CO(n37340));
    SB_LUT4 add_3029_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n37338), 
            .O(n6952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_5 (.CI(n37338), .I0(n2463), .I1(n97), .CO(n37339));
    SB_LUT4 add_3029_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n37337), 
            .O(n6953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_4 (.CI(n37337), .I0(n2464), .I1(n98), .CO(n37338));
    SB_LUT4 add_3029_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n37336), 
            .O(n6954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4285));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4287));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4288));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4295));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1764_3_lut_3_lut (.I0(n2642), .I1(n6991), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4290));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3029_3 (.CI(n37336), .I0(n2465), .I1(n99), .CO(n37337));
    SB_LUT4 add_3029_2_lut (.I0(GND_net), .I1(n387_adj_3993), .I2(n558), 
            .I3(VCC_net), .O(n6955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_2 (.CI(VCC_net), .I0(n387_adj_3993), .I1(n558), 
            .CO(n37336));
    SB_LUT4 div_12_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3028_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n37335), 
            .O(n6915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3028_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n37334), 
            .O(n6916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_19 (.CI(n37334), .I0(n2358), .I1(n83), .CO(n37335));
    SB_LUT4 add_3028_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n37333), 
            .O(n6917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_18 (.CI(n37333), .I0(n2359), .I1(n84), .CO(n37334));
    SB_LUT4 add_3028_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n37332), 
            .O(n6918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_17 (.CI(n37332), .I0(n2360), .I1(n85), .CO(n37333));
    SB_LUT4 add_3028_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n37331), 
            .O(n6919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31563_4_lut (.I0(n31_adj_4295), .I1(n19_adj_4288), .I2(n17_adj_4287), 
            .I3(n15_adj_4285), .O(n47077));
    defparam i31563_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3028_16 (.CI(n37331), .I0(n2361), .I1(n86), .CO(n37332));
    SB_LUT4 add_3028_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n37330), 
            .O(n6920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_15 (.CI(n37330), .I0(n2362), .I1(n87), .CO(n37331));
    SB_LUT4 add_3028_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n37329), 
            .O(n6921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_14 (.CI(n37329), .I0(n2363), .I1(n88), .CO(n37330));
    SB_LUT4 add_3028_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n37328), 
            .O(n6922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_13 (.CI(n37328), .I0(n2364), .I1(n89), .CO(n37329));
    SB_LUT4 add_3028_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n37327), 
            .O(n6923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_12 (.CI(n37327), .I0(n2365), .I1(n90), .CO(n37328));
    SB_LUT4 add_3028_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n37326), 
            .O(n6924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_11 (.CI(n37326), .I0(n2366), .I1(n91), .CO(n37327));
    SB_LUT4 add_3028_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n37325), 
            .O(n6925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_10 (.CI(n37325), .I0(n2367), .I1(n92), .CO(n37326));
    SB_LUT4 add_3028_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n37324), 
            .O(n6926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32187_4_lut (.I0(n13_adj_4283), .I1(n11_adj_4281), .I2(n2637), 
            .I3(n98), .O(n47701));
    defparam i32187_4_lut.LUT_INIT = 16'hfeef;
    SB_CARRY add_3028_9 (.CI(n37324), .I0(n2368), .I1(n93), .CO(n37325));
    SB_LUT4 add_3028_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n37323), 
            .O(n6927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_8 (.CI(n37323), .I0(n2369), .I1(n94), .CO(n37324));
    SB_LUT4 add_3028_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n37322), 
            .O(n6928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_7 (.CI(n37322), .I0(n2370), .I1(n95), .CO(n37323));
    SB_LUT4 add_3028_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n37321), 
            .O(n6929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_6 (.CI(n37321), .I0(n2371), .I1(n96), .CO(n37322));
    SB_LUT4 mux_23_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[0]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_3028_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n37320), 
            .O(n6930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_25[0]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3028_5 (.CI(n37320), .I0(n2372), .I1(n97), .CO(n37321));
    SB_LUT4 i32503_4_lut (.I0(n19_adj_4288), .I1(n17_adj_4287), .I2(n15_adj_4285), 
            .I3(n47701), .O(n48017));
    defparam i32503_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_3028_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n37319), 
            .O(n6931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_4 (.CI(n37319), .I0(n2373), .I1(n98), .CO(n37320));
    SB_LUT4 add_3028_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n37318), 
            .O(n6932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_3 (.CI(n37318), .I0(n2374), .I1(n99), .CO(n37319));
    SB_LUT4 add_3028_2_lut (.I0(GND_net), .I1(n386), .I2(n558), .I3(VCC_net), 
            .O(n6933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_2 (.CI(VCC_net), .I0(n386), .I1(n558), .CO(n37318));
    SB_LUT4 add_3027_19_lut (.I0(GND_net), .I1(n2264_adj_3994), .I2(n83), 
            .I3(n37317), .O(n6895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3027_18_lut (.I0(GND_net), .I1(n2265_adj_3995), .I2(n84), 
            .I3(n37316), .O(n6896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_18 (.CI(n37316), .I0(n2265_adj_3995), .I1(n84), 
            .CO(n37317));
    SB_LUT4 add_3027_17_lut (.I0(GND_net), .I1(n2266_adj_3996), .I2(n85), 
            .I3(n37315), .O(n6897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_17 (.CI(n37315), .I0(n2266_adj_3996), .I1(n85), 
            .CO(n37316));
    SB_LUT4 add_3027_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n37314), 
            .O(n6898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_16 (.CI(n37314), .I0(n2267), .I1(n86), .CO(n37315));
    SB_LUT4 add_3027_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n37313), 
            .O(n6899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10973_3_lut (.I0(n23783), .I1(r_Bit_Index[0]), .I2(n23649), 
            .I3(GND_net), .O(n24391));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10973_3_lut.LUT_INIT = 16'h1414;
    SB_CARRY add_3027_15 (.CI(n37313), .I0(n2268), .I1(n87), .CO(n37314));
    SB_LUT4 add_3027_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n37312), 
            .O(n6900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_14 (.CI(n37312), .I0(n2269), .I1(n88), .CO(n37313));
    SB_LUT4 add_3027_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n37311), 
            .O(n6901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_13 (.CI(n37311), .I0(n2270), .I1(n89), .CO(n37312));
    SB_LUT4 add_3027_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n37310), 
            .O(n6902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_12 (.CI(n37310), .I0(n2271), .I1(n90), .CO(n37311));
    SB_LUT4 add_3027_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n37309), 
            .O(n6903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_11 (.CI(n37309), .I0(n2272), .I1(n91), .CO(n37310));
    SB_LUT4 add_3027_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n37308), 
            .O(n6904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_10 (.CI(n37308), .I0(n2273), .I1(n92), .CO(n37309));
    SB_LUT4 add_3027_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n37307), 
            .O(n6905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_9 (.CI(n37307), .I0(n2274), .I1(n93), .CO(n37308));
    SB_LUT4 add_3027_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n37306), 
            .O(n6906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_8 (.CI(n37306), .I0(n2275), .I1(n94), .CO(n37307));
    SB_LUT4 add_3027_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n37305), 
            .O(n6907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_7 (.CI(n37305), .I0(n2276), .I1(n95), .CO(n37306));
    SB_LUT4 add_3027_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n37304), 
            .O(n6908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_6 (.CI(n37304), .I0(n2277), .I1(n96), .CO(n37305));
    SB_LUT4 i32501_4_lut (.I0(n25_adj_4292), .I1(n23_adj_4291), .I2(n21_adj_4290), 
            .I3(n48017), .O(n48015));
    defparam i32501_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31567_4_lut (.I0(n31_adj_4295), .I1(n29_adj_4294), .I2(n27_adj_4293), 
            .I3(n48015), .O(n47081));
    defparam i31567_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3027_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n37303), 
            .O(n6909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_5 (.CI(n37303), .I0(n2278), .I1(n97), .CO(n37304));
    SB_LUT4 add_3027_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n37302), 
            .O(n6910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1722_i8_4_lut (.I0(n389), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_4279));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY add_3027_4 (.CI(n37302), .I0(n2279), .I1(n98), .CO(n37303));
    SB_LUT4 add_3027_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n37301), 
            .O(n6911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_3 (.CI(n37301), .I0(n2280), .I1(n99), .CO(n37302));
    SB_LUT4 add_3027_2_lut (.I0(GND_net), .I1(n385), .I2(n558), .I3(VCC_net), 
            .O(n6912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32603_3_lut (.I0(n8_adj_4279), .I1(n87), .I2(n31_adj_4295), 
            .I3(GND_net), .O(n48117));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32603_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32604_3_lut (.I0(n48117), .I1(n86), .I2(n33_adj_4296), .I3(GND_net), 
            .O(n48118));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32604_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1722_i34_3_lut (.I0(n16_adj_4286), .I1(n83), 
            .I2(n39_adj_4300), .I3(GND_net), .O(n34_adj_4297));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31557_4_lut (.I0(n37_adj_4299), .I1(n35_adj_4298), .I2(n33_adj_4296), 
            .I3(n47077), .O(n47071));
    defparam i31557_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_i274_4_lut_4_lut (.I0(n392), .I1(n99), .I2(n2_adj_3955), 
            .I3(n5_adj_4363), .O(n43347));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i274_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i32985_4_lut (.I0(n34_adj_4297), .I1(n14_adj_4284), .I2(n39_adj_4300), 
            .I3(n47069), .O(n48499));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32985_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32052_3_lut (.I0(n48118), .I1(n85), .I2(n35_adj_4298), .I3(GND_net), 
            .O(n47566));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32052_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32605_3_lut (.I0(n10_adj_4280), .I1(n90), .I2(n25_adj_4292), 
            .I3(GND_net), .O(n48119));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32605_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32606_3_lut (.I0(n48119), .I1(n89), .I2(n27_adj_4293), .I3(GND_net), 
            .O(n48120));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32606_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32173_4_lut (.I0(n27_adj_4293), .I1(n25_adj_4292), .I2(n23_adj_4291), 
            .I3(n47089), .O(n47687));
    defparam i32173_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_12_LessThan_1722_i20_3_lut (.I0(n12_adj_4282), .I1(n91), 
            .I2(n23_adj_4291), .I3(GND_net), .O(n20_adj_4289));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32050_3_lut (.I0(n48120), .I1(n88), .I2(n29_adj_4294), .I3(GND_net), 
            .O(n47564));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32050_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32757_4_lut (.I0(n37_adj_4299), .I1(n35_adj_4298), .I2(n33_adj_4296), 
            .I3(n47081), .O(n48271));
    defparam i32757_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33096_4_lut (.I0(n47566), .I1(n48499), .I2(n39_adj_4300), 
            .I3(n47071), .O(n48610));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33096_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32451_4_lut (.I0(n47564), .I1(n20_adj_4289), .I2(n29_adj_4294), 
            .I3(n47687), .O(n47965));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32451_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33124_4_lut (.I0(n47965), .I1(n48610), .I2(n39_adj_4300), 
            .I3(n48271), .O(n48638));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33124_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33125_3_lut (.I0(n48638), .I1(n82), .I2(n2621), .I3(GND_net), 
            .O(n48639));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33125_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33117_3_lut (.I0(n48639), .I1(n81), .I2(n2620), .I3(GND_net), 
            .O(n48631));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33117_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i32802_3_lut (.I0(n48631), .I1(n80), .I2(n2619), .I3(GND_net), 
            .O(n48316));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32802_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut (.I0(n48316), .I1(n22633), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4276));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4278));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4274));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n388));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4277));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31697_3_lut_3_lut (.I0(n392), .I1(n558), .I2(n369), .I3(GND_net), 
            .O(n510));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31697_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_12_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4271));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4272));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4268));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4269));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4270));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_742_i36_4_lut (.I0(n375), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_LessThan_742_i40_3_lut (.I0(n38_adj_4081), .I1(n96), 
            .I2(n41), .I3(GND_net), .O(n40_adj_4082));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33022_4_lut (.I0(n40_adj_4082), .I1(n36), .I2(n41), .I3(n46873), 
            .O(n48536));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33022_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_12_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4259));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4261));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33023_3_lut (.I0(n48536), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n48537));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33023_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i32972_3_lut (.I0(n48537), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n48486));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32972_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1434 (.I0(n48486), .I1(n22591), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1434.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4263));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4265));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31692_3_lut_3_lut (.I0(n533), .I1(n558), .I2(n370), .I3(GND_net), 
            .O(n649));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31692_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_12_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4266));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3027_2 (.CI(VCC_net), .I0(n385), .I1(n558), .CO(n37301));
    SB_LUT4 div_12_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4273));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3026_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n37300), 
            .O(n6876)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i368_4_lut_4_lut (.I0(n533), .I1(n99), .I2(n2_adj_3954), 
            .I3(n510), .O(n648));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i368_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 add_3026_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n37299), 
            .O(n6877)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31605_4_lut (.I0(n33_adj_4273), .I1(n21_adj_4266), .I2(n19_adj_4265), 
            .I3(n17_adj_4263), .O(n47119));
    defparam i31605_4_lut.LUT_INIT = 16'haaab;
    SB_IO PIN_9_pad (.PACKAGE_PIN(PIN_9), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_9_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_9_pad.PIN_TYPE = 6'b000001;
    defparam PIN_9_pad.PULLUP = 1'b0;
    defparam PIN_9_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_3026_17 (.CI(n37299), .I0(n2169), .I1(n85), .CO(n37300));
    SB_LUT4 i32233_4_lut (.I0(n15_adj_4261), .I1(n13_adj_4259), .I2(n2552), 
            .I3(n98), .O(n47747));
    defparam i32233_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i32527_4_lut (.I0(n21_adj_4266), .I1(n19_adj_4265), .I2(n17_adj_4263), 
            .I3(n47747), .O(n48041));
    defparam i32527_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_3026_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n37298), 
            .O(n6878)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10500_3_lut (.I0(n23785), .I1(r_Bit_Index_adj_4404[0]), .I2(n23655), 
            .I3(GND_net), .O(n23918));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10500_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 div_12_i367_4_lut_4_lut (.I0(n533), .I1(n98), .I2(n4_adj_3953), 
            .I3(n43347), .O(n43349));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i367_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_CARRY add_3026_16 (.CI(n37298), .I0(n2170), .I1(n86), .CO(n37299));
    SB_LUT4 i32525_4_lut (.I0(n27_adj_4270), .I1(n25_adj_4269), .I2(n23_adj_4268), 
            .I3(n48041), .O(n48039));
    defparam i32525_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31609_4_lut (.I0(n33_adj_4273), .I1(n31_adj_4272), .I2(n29_adj_4271), 
            .I3(n48039), .O(n47123));
    defparam i31609_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1665_i10_4_lut (.I0(n388), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4257));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_3026_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n37297), 
            .O(n6879)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32611_3_lut (.I0(n10_adj_4257), .I1(n87), .I2(n33_adj_4273), 
            .I3(GND_net), .O(n48125));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32611_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10497_2_lut (.I0(n23914), .I1(n23913), .I2(GND_net), .I3(GND_net), 
            .O(n23915));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10497_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3026_15 (.CI(n37297), .I0(n2171), .I1(n87), .CO(n37298));
    SB_LUT4 add_3026_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n37296), 
            .O(n6880)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32612_3_lut (.I0(n48125), .I1(n86), .I2(n35_adj_4274), .I3(GND_net), 
            .O(n48126));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32612_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3026_14 (.CI(n37296), .I0(n2172), .I1(n88), .CO(n37297));
    SB_LUT4 add_3026_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n37295), 
            .O(n6881)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1665_i36_3_lut (.I0(n18_adj_4264), .I1(n83), 
            .I2(n41_adj_4278), .I3(GND_net), .O(n36_adj_4275));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31601_4_lut (.I0(n39_adj_4277), .I1(n37_adj_4276), .I2(n35_adj_4274), 
            .I3(n47119), .O(n47115));
    defparam i31601_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3026_13 (.CI(n37295), .I0(n2173), .I1(n89), .CO(n37296));
    SB_LUT4 add_3026_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n37294), 
            .O(n6882)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_12 (.CI(n37294), .I0(n2174), .I1(n90), .CO(n37295));
    SB_LUT4 add_3026_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n37293), 
            .O(n6883)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_11 (.CI(n37293), .I0(n2175), .I1(n91), .CO(n37294));
    SB_LUT4 add_3026_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n37292), 
            .O(n6884)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32983_4_lut (.I0(n36_adj_4275), .I1(n16_adj_4262), .I2(n41_adj_4278), 
            .I3(n47111), .O(n48497));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32983_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32040_3_lut (.I0(n48126), .I1(n85), .I2(n37_adj_4276), .I3(GND_net), 
            .O(n47554));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32040_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3026_10 (.CI(n37292), .I0(n2176), .I1(n92), .CO(n37293));
    SB_LUT4 add_3026_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n37291), 
            .O(n6885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_9 (.CI(n37291), .I0(n2177), .I1(n93), .CO(n37292));
    SB_LUT4 add_3026_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n37290), 
            .O(n6886)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_23_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[1]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_25[1]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3026_8 (.CI(n37290), .I0(n2178), .I1(n94), .CO(n37291));
    SB_LUT4 add_3026_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n37289), 
            .O(n6887)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_7 (.CI(n37289), .I0(n2179), .I1(n95), .CO(n37290));
    SB_LUT4 div_12_LessThan_1665_i22_3_lut (.I0(n14_adj_4260), .I1(n91), 
            .I2(n25_adj_4269), .I3(GND_net), .O(n22_adj_4267));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3026_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n37288), 
            .O(n6888)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32981_4_lut (.I0(n22_adj_4267), .I1(n12_adj_4258), .I2(n25_adj_4269), 
            .I3(n47135), .O(n48495));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32981_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3026_6 (.CI(n37288), .I0(n2180), .I1(n96), .CO(n37289));
    SB_LUT4 add_3026_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n37287), 
            .O(n6889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_5 (.CI(n37287), .I0(n2181), .I1(n97), .CO(n37288));
    SB_LUT4 i32982_3_lut (.I0(n48495), .I1(n90), .I2(n27_adj_4270), .I3(GND_net), 
            .O(n48496));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32982_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3026_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n37286), 
            .O(n6890)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_4 (.CI(n37286), .I0(n2182), .I1(n98), .CO(n37287));
    SB_LUT4 add_3026_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n37285), 
            .O(n6891)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32848_3_lut (.I0(n48496), .I1(n89), .I2(n29_adj_4271), .I3(GND_net), 
            .O(n48362));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32848_3_lut.LUT_INIT = 16'h3a3a;
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_8_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b000001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_3026_3 (.CI(n37285), .I0(n2183), .I1(n99), .CO(n37286));
    SB_LUT4 add_3026_2_lut (.I0(GND_net), .I1(n384), .I2(n558), .I3(VCC_net), 
            .O(n6892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_23_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[2]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32767_4_lut (.I0(n39_adj_4277), .I1(n37_adj_4276), .I2(n35_adj_4274), 
            .I3(n47123), .O(n48281));
    defparam i32767_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3026_2 (.CI(VCC_net), .I0(n384), .I1(n558), .CO(n37285));
    SB_LUT4 add_3025_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n37284), 
            .O(n6858)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33094_4_lut (.I0(n47554), .I1(n48497), .I2(n41_adj_4278), 
            .I3(n47115), .O(n48608));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33094_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3025_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n37283), 
            .O(n6859)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_25[2]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i460_4_lut_4_lut (.I0(n671), .I1(n99), .I2(n2), .I3(n649), 
            .O(n784));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i460_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_CARRY add_3025_16 (.CI(n37283), .I0(n2070), .I1(n86), .CO(n37284));
    SB_LUT4 add_3025_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n37282), 
            .O(n6860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_15 (.CI(n37282), .I0(n2071), .I1(n87), .CO(n37283));
    SB_LUT4 add_3025_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n37281), 
            .O(n6861)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_14 (.CI(n37281), .I0(n2072), .I1(n88), .CO(n37282));
    SB_LUT4 add_3025_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n37280), 
            .O(n6862)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_13 (.CI(n37280), .I0(n2073), .I1(n89), .CO(n37281));
    SB_LUT4 add_3025_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n37279), 
            .O(n6863)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_12 (.CI(n37279), .I0(n2074), .I1(n90), .CO(n37280));
    SB_LUT4 add_3025_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n37278), 
            .O(n6864)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_11 (.CI(n37278), .I0(n2075), .I1(n91), .CO(n37279));
    SB_LUT4 add_3025_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n37277), 
            .O(n6865)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_10 (.CI(n37277), .I0(n2076), .I1(n92), .CO(n37278));
    SB_LUT4 add_3025_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n37276), 
            .O(n6866)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_9 (.CI(n37276), .I0(n2077), .I1(n93), .CO(n37277));
    SB_LUT4 add_3025_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n37275), 
            .O(n6867)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_8 (.CI(n37275), .I0(n2078), .I1(n94), .CO(n37276));
    SB_LUT4 add_3025_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n37274), 
            .O(n6868)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_7 (.CI(n37274), .I0(n2079), .I1(n95), .CO(n37275));
    SB_LUT4 add_3025_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n37273), 
            .O(n6869)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32038_3_lut (.I0(n48362), .I1(n88), .I2(n31_adj_4272), .I3(GND_net), 
            .O(n47552));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32038_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3025_6 (.CI(n37273), .I0(n2080), .I1(n96), .CO(n37274));
    SB_LUT4 add_3025_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n37272), 
            .O(n6870)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_5 (.CI(n37272), .I0(n2081), .I1(n97), .CO(n37273));
    SB_LUT4 add_3025_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n37271), 
            .O(n6871)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_4 (.CI(n37271), .I0(n2082), .I1(n98), .CO(n37272));
    SB_LUT4 add_3025_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n37270), 
            .O(n6872)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_3 (.CI(n37270), .I0(n2083), .I1(n99), .CO(n37271));
    SB_LUT4 add_3025_2_lut (.I0(GND_net), .I1(n383), .I2(n558), .I3(VCC_net), 
            .O(n6873)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_2 (.CI(VCC_net), .I0(n383), .I1(n558), .CO(n37270));
    SB_LUT4 add_3024_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n37269), 
            .O(n6841)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3024_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n37268), 
            .O(n6842)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_15 (.CI(n37268), .I0(n1968), .I1(n87), .CO(n37269));
    SB_LUT4 add_3024_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n37267), 
            .O(n6843)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_14 (.CI(n37267), .I0(n1969), .I1(n88), .CO(n37268));
    SB_LUT4 add_3024_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n37266), 
            .O(n6844)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33122_4_lut (.I0(n47552), .I1(n48608), .I2(n41_adj_4278), 
            .I3(n48281), .O(n48636));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33122_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3024_13 (.CI(n37266), .I0(n1970), .I1(n89), .CO(n37267));
    SB_LUT4 mux_23_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[3]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_3024_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n37265), 
            .O(n6845)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_12 (.CI(n37265), .I0(n1971), .I1(n90), .CO(n37266));
    SB_LUT4 i33123_3_lut (.I0(n48636), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n48637));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33123_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 add_3024_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n37264), 
            .O(n6846)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_11_lut.LUT_INIT = 16'hC33C;
    SB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_6_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b011001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_24_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b000001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i33121_3_lut (.I0(n48637), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n48635));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33121_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1435 (.I0(n48635), .I1(n22630), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1435.LUT_INIT = 16'hceef;
    SB_CARRY add_3024_11 (.CI(n37264), .I0(n1972), .I1(n91), .CO(n37265));
    SB_LUT4 add_3024_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n37263), 
            .O(n6847)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_10 (.CI(n37263), .I0(n1973), .I1(n92), .CO(n37264));
    SB_LUT4 add_3024_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n37262), 
            .O(n6848)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i458_4_lut_4_lut (.I0(n671), .I1(n97), .I2(n6), .I3(n43349), 
            .O(n43351));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i458_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_12_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i31688_3_lut_3_lut (.I0(n671), .I1(n558), .I2(n371), .I3(GND_net), 
            .O(n785));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31688_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 mux_22_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_25[3]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3024_9 (.CI(n37262), .I0(n1974), .I1(n93), .CO(n37263));
    SB_LUT4 add_3024_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n37261), 
            .O(n6849)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_8 (.CI(n37261), .I0(n1975), .I1(n94), .CO(n37262));
    SB_LUT4 add_3024_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n37260), 
            .O(n6850)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n22531), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_3985));   // verilog/TinyFPGA_B.v(146[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_3024_7 (.CI(n37260), .I0(n1976), .I1(n95), .CO(n37261));
    SB_LUT4 div_12_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4254));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3024_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n37259), 
            .O(n6851)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_6 (.CI(n37259), .I0(n1977), .I1(n96), .CO(n37260));
    SB_LUT4 add_3024_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n37258), 
            .O(n6852)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1436 (.I0(control_mode[0]), .I1(n22531), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_3959));   // verilog/TinyFPGA_B.v(146[5:22])
    defparam i1_2_lut_3_lut_adj_1436.LUT_INIT = 16'hefef;
    SB_CARRY add_3024_5 (.CI(n37258), .I0(n1978), .I1(n97), .CO(n37259));
    SB_LUT4 add_3024_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n37257), 
            .O(n6853)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4252));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3024_4 (.CI(n37257), .I0(n1979), .I1(n98), .CO(n37258));
    SB_LUT4 add_3024_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n37256), 
            .O(n6854)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_3 (.CI(n37256), .I0(n1980), .I1(n99), .CO(n37257));
    SB_LUT4 div_12_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4256));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3024_2_lut (.I0(GND_net), .I1(n382), .I2(n558), .I3(VCC_net), 
            .O(n6855)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_2 (.CI(VCC_net), .I0(n382), .I1(n558), .CO(n37256));
    SB_LUT4 add_3023_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n37255), 
            .O(n6825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4255));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3023_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n37254), 
            .O(n6826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_23_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[4]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_3023_14 (.CI(n37254), .I0(n1863), .I1(n88), .CO(n37255));
    SB_LUT4 mux_22_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_25[4]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3023_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n37253), 
            .O(n6827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n387_adj_3993));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3023_13 (.CI(n37253), .I0(n1864), .I1(n89), .CO(n37254));
    SB_LUT4 add_3023_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n37252), 
            .O(n6828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_12 (.CI(n37252), .I0(n1865), .I1(n90), .CO(n37253));
    SB_LUT4 add_3023_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n37251), 
            .O(n6829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_11 (.CI(n37251), .I0(n1866), .I1(n91), .CO(n37252));
    SB_LUT4 add_3023_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n37250), 
            .O(n6830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_10 (.CI(n37250), .I0(n1867), .I1(n92), .CO(n37251));
    SB_LUT4 add_3023_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n37249), 
            .O(n6831)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4249));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3023_9 (.CI(n37249), .I0(n1868), .I1(n93), .CO(n37250));
    SB_LUT4 add_3023_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n37248), 
            .O(n6832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_8_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_4_pad (.PACKAGE_PIN(PIN_4), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_4_c_2)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_4_pad.PIN_TYPE = 6'b011001;
    defparam PIN_4_pad.PULLUP = 1'b0;
    defparam PIN_4_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_3_pad (.PACKAGE_PIN(PIN_3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_3_c_3)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_3_pad.PIN_TYPE = 6'b011001;
    defparam PIN_3_pad.PULLUP = 1'b0;
    defparam PIN_3_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_12_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4250));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3023_8 (.CI(n37248), .I0(n1869), .I1(n94), .CO(n37249));
    SB_LUT4 add_3023_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n37247), 
            .O(n6833)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_7 (.CI(n37247), .I0(n1870), .I1(n95), .CO(n37248));
    SB_LUT4 div_12_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4246));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 mux_23_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[5]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_12_LessThan_657_i38_4_lut (.I0(n374), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4247));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 mux_22_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_25[5]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4248));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3023_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n37246), 
            .O(n6834)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i459_4_lut_4_lut (.I0(n671), .I1(n98), .I2(n4), .I3(n648), 
            .O(n783));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i459_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_CARRY add_3023_6 (.CI(n37246), .I0(n1871), .I1(n96), .CO(n37247));
    SB_LUT4 mux_23_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[6]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_3023_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n37245), 
            .O(n6835)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_5 (.CI(n37245), .I0(n1872), .I1(n97), .CO(n37246));
    SB_LUT4 mux_22_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_25[6]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3023_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n37244), 
            .O(n6836)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4237));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3023_4 (.CI(n37244), .I0(n1873), .I1(n98), .CO(n37245));
    SB_LUT4 add_3023_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n37243), 
            .O(n6837)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_3 (.CI(n37243), .I0(n1874), .I1(n99), .CO(n37244));
    SB_LUT4 add_3023_2_lut (.I0(GND_net), .I1(n381), .I2(n558), .I3(VCC_net), 
            .O(n6838)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_23_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[7]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_12_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4239));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3023_2 (.CI(VCC_net), .I0(n381), .I1(n558), .CO(n37243));
    SB_LUT4 add_3021_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n37242), 
            .O(n6784)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_25[7]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4241));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3021_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n37241), 
            .O(n6785)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_13 (.CI(n37241), .I0(n1755), .I1(n89), .CO(n37242));
    SB_LUT4 add_3021_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n37240), 
            .O(n6786)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4243));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3021_12 (.CI(n37240), .I0(n1756), .I1(n90), .CO(n37241));
    SB_LUT4 add_3021_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n37239), 
            .O(n6787)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_11 (.CI(n37239), .I0(n1757), .I1(n91), .CO(n37240));
    SB_LUT4 div_12_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4244));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3021_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n37238), 
            .O(n6788)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4251));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31653_4_lut (.I0(n35_adj_4251), .I1(n23_adj_4244), .I2(n21_adj_4243), 
            .I3(n19_adj_4241), .O(n47167));
    defparam i31653_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3021_10 (.CI(n37238), .I0(n1758), .I1(n92), .CO(n37239));
    SB_LUT4 add_3021_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n37237), 
            .O(n6789)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_9 (.CI(n37237), .I0(n1759), .I1(n93), .CO(n37238));
    SB_LUT4 i32275_4_lut (.I0(n17_adj_4239), .I1(n15_adj_4237), .I2(n2464), 
            .I3(n98), .O(n47789));
    defparam i32275_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 add_3021_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n37236), 
            .O(n6790)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32545_4_lut (.I0(n23_adj_4244), .I1(n21_adj_4243), .I2(n19_adj_4241), 
            .I3(n47789), .O(n48059));
    defparam i32545_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_3021_8 (.CI(n37236), .I0(n1760), .I1(n94), .CO(n37237));
    SB_LUT4 add_3021_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n37235), 
            .O(n6791)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_7 (.CI(n37235), .I0(n1761), .I1(n95), .CO(n37236));
    SB_LUT4 add_3021_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n37234), 
            .O(n6792)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_6 (.CI(n37234), .I0(n1762), .I1(n96), .CO(n37235));
    SB_LUT4 add_3021_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n37233), 
            .O(n6793)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32541_4_lut (.I0(n29_adj_4248), .I1(n27_adj_4247), .I2(n25_adj_4246), 
            .I3(n48059), .O(n48055));
    defparam i32541_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_12_i1765_3_lut_3_lut (.I0(n2642), .I1(n6992), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31657_4_lut (.I0(n35_adj_4251), .I1(n33_adj_4250), .I2(n31_adj_4249), 
            .I3(n48055), .O(n47171));
    defparam i31657_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3021_5 (.CI(n37233), .I0(n1763), .I1(n97), .CO(n37234));
    SB_LUT4 div_12_LessThan_1606_i12_4_lut (.I0(n387_adj_3993), .I1(n99), 
            .I2(n2465), .I3(n558), .O(n12_adj_4235));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32615_3_lut (.I0(n12_adj_4235), .I1(n87), .I2(n35_adj_4251), 
            .I3(GND_net), .O(n48129));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32615_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3021_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n37232), 
            .O(n6794)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_23_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[8]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_3021_4 (.CI(n37232), .I0(n1764), .I1(n98), .CO(n37233));
    SB_LUT4 add_3021_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n37231), 
            .O(n6795)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_25[8]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3021_3 (.CI(n37231), .I0(n1765), .I1(n99), .CO(n37232));
    SB_LUT4 add_3021_2_lut (.I0(GND_net), .I1(n380), .I2(n558), .I3(VCC_net), 
            .O(n6796)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_2 (.CI(VCC_net), .I0(n380), .I1(n558), .CO(n37231));
    SB_LUT4 add_3019_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n37230), 
            .O(n6743)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3019_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n37229), 
            .O(n6744)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_12 (.CI(n37229), .I0(n1644), .I1(n90), .CO(n37230));
    SB_LUT4 add_3019_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n37228), 
            .O(n6745)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_11 (.CI(n37228), .I0(n1645), .I1(n91), .CO(n37229));
    SB_LUT4 div_12_LessThan_1606_i38_3_lut (.I0(n20_adj_4242), .I1(n83), 
            .I2(n43_adj_4256), .I3(GND_net), .O(n38_adj_4253));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3019_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n37227), 
            .O(n6746)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32616_3_lut (.I0(n48129), .I1(n86), .I2(n37_adj_4252), .I3(GND_net), 
            .O(n48130));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32616_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31647_4_lut (.I0(n41_adj_4255), .I1(n39_adj_4254), .I2(n37_adj_4252), 
            .I3(n47167), .O(n47161));
    defparam i31647_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3019_10 (.CI(n37227), .I0(n1646), .I1(n92), .CO(n37228));
    SB_LUT4 add_3019_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n37226), 
            .O(n6747)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_9 (.CI(n37226), .I0(n1647), .I1(n93), .CO(n37227));
    SB_LUT4 add_3019_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n37225), 
            .O(n6748)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_8 (.CI(n37225), .I0(n1648), .I1(n94), .CO(n37226));
    SB_LUT4 add_3019_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n37224), 
            .O(n6749)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_7 (.CI(n37224), .I0(n1649), .I1(n95), .CO(n37225));
    SB_LUT4 add_3019_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n37223), 
            .O(n6750)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32957_4_lut (.I0(n38_adj_4253), .I1(n18_adj_4240), .I2(n43_adj_4256), 
            .I3(n47157), .O(n48471));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32957_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3019_6 (.CI(n37223), .I0(n1650), .I1(n96), .CO(n37224));
    SB_LUT4 i32034_3_lut (.I0(n48130), .I1(n85), .I2(n39_adj_4254), .I3(GND_net), 
            .O(n47548));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32034_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3019_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n37222), 
            .O(n6751)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_657_i42_3_lut (.I0(n40_adj_4078), .I1(n96), 
            .I2(n43), .I3(GND_net), .O(n42_adj_4079));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3019_5 (.CI(n37222), .I0(n1651), .I1(n97), .CO(n37223));
    SB_LUT4 i32831_4_lut (.I0(n42_adj_4079), .I1(n38), .I2(n43), .I3(n46881), 
            .O(n48345));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32831_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32832_3_lut (.I0(n48345), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n48346));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32832_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_12_LessThan_1606_i24_3_lut (.I0(n16_adj_4238), .I1(n91), 
            .I2(n27_adj_4247), .I3(GND_net), .O(n24_adj_4245));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_4_lut_adj_1437 (.I0(n48346), .I1(n22588), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1437.LUT_INIT = 16'hceef;
    SB_LUT4 i22649_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4074), .I3(GND_net), 
            .O(n8_adj_4073));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22649_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 add_3019_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n37221), 
            .O(n6752)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32979_4_lut (.I0(n24_adj_4245), .I1(n14_adj_4236), .I2(n27_adj_4247), 
            .I3(n47181), .O(n48493));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32979_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32980_3_lut (.I0(n48493), .I1(n90), .I2(n29_adj_4248), .I3(GND_net), 
            .O(n48494));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32980_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32852_3_lut (.I0(n48494), .I1(n89), .I2(n31_adj_4249), .I3(GND_net), 
            .O(n48366));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32852_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3019_4 (.CI(n37221), .I0(n1652), .I1(n98), .CO(n37222));
    SB_LUT4 add_3019_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n37220), 
            .O(n6753)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32775_4_lut (.I0(n41_adj_4255), .I1(n39_adj_4254), .I2(n37_adj_4252), 
            .I3(n47171), .O(n48289));
    defparam i32775_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33080_4_lut (.I0(n47548), .I1(n48471), .I2(n43_adj_4256), 
            .I3(n47161), .O(n48594));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33080_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_12_i549_4_lut_4_lut (.I0(n806), .I1(n98), .I2(n4_adj_4075), 
            .I3(n784), .O(n916));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i549_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_CARRY add_3019_3 (.CI(n37220), .I0(n1653), .I1(n99), .CO(n37221));
    SB_LUT4 add_3019_2_lut (.I0(GND_net), .I1(n379), .I2(n558), .I3(VCC_net), 
            .O(n6754)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_2 (.CI(VCC_net), .I0(n379), .I1(n558), .CO(n37220));
    SB_LUT4 i32032_3_lut (.I0(n48366), .I1(n88), .I2(n33_adj_4250), .I3(GND_net), 
            .O(n47546));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32032_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3018_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n37219), 
            .O(n6730)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3018_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n37218), 
            .O(n6731)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_11 (.CI(n37218), .I0(n1530), .I1(n91), .CO(n37219));
    SB_LUT4 i33114_4_lut (.I0(n47546), .I1(n48594), .I2(n43_adj_4256), 
            .I3(n48289), .O(n48628));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33114_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i22641_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4075), .I3(GND_net), 
            .O(n6_adj_4074));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22641_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_12_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33115_3_lut (.I0(n48628), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n48629));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33115_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1438 (.I0(n48629), .I1(n22627), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1438.LUT_INIT = 16'hceef;
    SB_LUT4 i31687_3_lut_3_lut (.I0(n806), .I1(n558), .I2(n372), .I3(GND_net), 
            .O(n918));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31687_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 add_3018_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n37217), 
            .O(n6732)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_10 (.CI(n37217), .I0(n1531), .I1(n92), .CO(n37218));
    SB_LUT4 div_12_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n373));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3018_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n37216), 
            .O(n6733)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_9 (.CI(n37216), .I0(n1532), .I1(n93), .CO(n37217));
    SB_LUT4 div_12_i550_4_lut_4_lut (.I0(n806), .I1(n99), .I2(n2_adj_4080), 
            .I3(n785), .O(n917));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i550_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 add_3018_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n37215), 
            .O(n6734)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_8 (.CI(n37215), .I0(n1533), .I1(n94), .CO(n37216));
    SB_LUT4 add_3018_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n37214), 
            .O(n6735)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_7 (.CI(n37214), .I0(n1534), .I1(n95), .CO(n37215));
    SB_LUT4 add_3018_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n37213), 
            .O(n6736)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_6 (.CI(n37213), .I0(n1535), .I1(n96), .CO(n37214));
    SB_LUT4 div_12_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4232));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4234));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4230));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 mux_23_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[9]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_12_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4227));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 mux_22_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_25[9]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4228));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n386));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3018_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n37212), 
            .O(n6737)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10894_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24312));   // verilog/coms.v(125[12] 284[6])
    defparam i10894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rx_i_I_0_1_lut (.I0(rx_i), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(LED_c));   // verilog/TinyFPGA_B.v(73[16:21])
    defparam rx_i_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3018_5 (.CI(n37212), .I0(n1536), .I1(n97), .CO(n37213));
    SB_LUT4 add_3018_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n37211), 
            .O(n6738)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10983_3_lut (.I0(encoder1_position[2]), .I1(n2264), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24401));   // quad.v(35[10] 41[6])
    defparam i10983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10984_3_lut (.I0(encoder1_position[3]), .I1(n2263), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24402));   // quad.v(35[10] 41[6])
    defparam i10984_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3018_4 (.CI(n37211), .I0(n1537), .I1(n98), .CO(n37212));
    SB_LUT4 add_3018_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n37210), 
            .O(n6739)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4233));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3018_3 (.CI(n37210), .I0(n1538), .I1(n99), .CO(n37211));
    SB_LUT4 add_3018_2_lut (.I0(GND_net), .I1(n378), .I2(n558), .I3(VCC_net), 
            .O(n6740)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_2 (.CI(VCC_net), .I0(n378), .I1(n558), .CO(n37210));
    SB_LUT4 add_3016_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n37209), 
            .O(n6690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3016_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n37208), 
            .O(n6691)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_10 (.CI(n37208), .I0(n1413), .I1(n92), .CO(n37209));
    SB_LUT4 add_3016_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n37207), 
            .O(n6692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_9 (.CI(n37207), .I0(n1414), .I1(n93), .CO(n37208));
    SB_LUT4 add_3016_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n37206), 
            .O(n6693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_8 (.CI(n37206), .I0(n1415), .I1(n94), .CO(n37207));
    SB_LUT4 add_3016_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n37205), 
            .O(n6694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4224));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4225));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_3978));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10895_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24313));   // verilog/coms.v(125[12] 284[6])
    defparam i10895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4226));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3016_7 (.CI(n37205), .I0(n1416), .I1(n95), .CO(n37206));
    SB_LUT4 add_3016_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n37204), 
            .O(n6695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_6 (.CI(n37204), .I0(n1417), .I1(n96), .CO(n37205));
    SB_LUT4 add_3016_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n37203), 
            .O(n6696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_5 (.CI(n37203), .I0(n1418), .I1(n97), .CO(n37204));
    SB_LUT4 add_3016_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n37202), 
            .O(n6697)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_4 (.CI(n37202), .I0(n1419), .I1(n98), .CO(n37203));
    SB_LUT4 add_3016_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n37201), 
            .O(n6698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_3 (.CI(n37201), .I0(n1420), .I1(n99), .CO(n37202));
    SB_LUT4 add_3016_2_lut (.I0(GND_net), .I1(n377), .I2(n558), .I3(VCC_net), 
            .O(n6699)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_2 (.CI(VCC_net), .I0(n377), .I1(n558), .CO(n37201));
    SB_LUT4 div_12_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4215));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 mux_23_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[10]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_12_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4217));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3014_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n37200), 
            .O(n6650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_25[10]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3014_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n37199), 
            .O(n6651)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_9 (.CI(n37199), .I0(n1293), .I1(n93), .CO(n37200));
    SB_LUT4 add_3014_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n37198), 
            .O(n6652)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_8 (.CI(n37198), .I0(n1294), .I1(n94), .CO(n37199));
    SB_LUT4 add_3014_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n37197), 
            .O(n6653)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_7 (.CI(n37197), .I0(n1295), .I1(n95), .CO(n37198));
    SB_LUT4 add_3014_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n37196), 
            .O(n6654)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_6 (.CI(n37196), .I0(n1296), .I1(n96), .CO(n37197));
    SB_LUT4 add_3014_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n37195), 
            .O(n6655)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_5 (.CI(n37195), .I0(n1297), .I1(n97), .CO(n37196));
    SB_LUT4 add_3014_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n37194), 
            .O(n6656)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_4 (.CI(n37194), .I0(n1298), .I1(n98), .CO(n37195));
    SB_LUT4 add_3014_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n37193), 
            .O(n6657)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_3 (.CI(n37193), .I0(n1299), .I1(n99), .CO(n37194));
    SB_LUT4 add_3014_2_lut (.I0(GND_net), .I1(n376), .I2(n558), .I3(VCC_net), 
            .O(n6658)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_2 (.CI(VCC_net), .I0(n376), .I1(n558), .CO(n37193));
    SB_LUT4 div_12_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4219));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4221));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4222));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4229));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31698_4_lut (.I0(n37_adj_4229), .I1(n25_adj_4222), .I2(n23_adj_4221), 
            .I3(n21_adj_4219), .O(n47212));
    defparam i31698_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32311_4_lut (.I0(n19_adj_4217), .I1(n17_adj_4215), .I2(n2373), 
            .I3(n98), .O(n47825));
    defparam i32311_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i32565_4_lut (.I0(n25_adj_4222), .I1(n23_adj_4221), .I2(n21_adj_4219), 
            .I3(n47825), .O(n48079));
    defparam i32565_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32561_4_lut (.I0(n31_adj_4226), .I1(n29_adj_4225), .I2(n27_adj_4224), 
            .I3(n48079), .O(n48075));
    defparam i32561_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31700_4_lut (.I0(n37_adj_4229), .I1(n35_adj_4228), .I2(n33_adj_4227), 
            .I3(n48075), .O(n47214));
    defparam i31700_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_23_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[11]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_12_LessThan_1545_i14_4_lut (.I0(n386), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4213));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 mux_22_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_25[11]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32621_3_lut (.I0(n14_adj_4213), .I1(n87), .I2(n37_adj_4229), 
            .I3(GND_net), .O(n48135));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32621_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32622_3_lut (.I0(n48135), .I1(n86), .I2(n39_adj_4230), .I3(GND_net), 
            .O(n48136));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32622_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1545_i40_3_lut (.I0(n22_adj_4220), .I1(n83), 
            .I2(n45_adj_4234), .I3(GND_net), .O(n40_adj_4231));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31689_4_lut (.I0(n43_adj_4233), .I1(n41_adj_4232), .I2(n39_adj_4230), 
            .I3(n47212), .O(n47203));
    defparam i31689_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32725_4_lut (.I0(n40_adj_4231), .I1(n20_adj_4218), .I2(n45_adj_4234), 
            .I3(n47199), .O(n48239));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32725_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32028_3_lut (.I0(n48136), .I1(n85), .I2(n41_adj_4232), .I3(GND_net), 
            .O(n47542));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32028_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1545_i26_3_lut (.I0(n18_adj_4216), .I1(n91), 
            .I2(n29_adj_4225), .I3(GND_net), .O(n26_adj_4223));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_3974));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32977_4_lut (.I0(n26_adj_4223), .I1(n16_adj_4214), .I2(n29_adj_4225), 
            .I3(n47226), .O(n48491));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32977_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_23_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[12]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_25[12]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n374));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22625_2_lut (.I0(n372), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4080));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22625_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_12_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_570_i40_4_lut (.I0(n373), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_LessThan_570_i44_3_lut (.I0(n42_adj_4076), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44_adj_4077));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32425_4_lut (.I0(n44_adj_4077), .I1(n40), .I2(n45), .I3(n46887), 
            .O(n47939));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32425_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1439 (.I0(n47939), .I1(n22585), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1439.LUT_INIT = 16'hceef;
    SB_LUT4 add_3011_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n37162), 
            .O(n6579)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3011_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n37161), 
            .O(n6580)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_8 (.CI(n37161), .I0(n1170), .I1(n94), .CO(n37162));
    SB_LUT4 add_3011_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n37160), 
            .O(n6581)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_7 (.CI(n37160), .I0(n1171), .I1(n95), .CO(n37161));
    SB_LUT4 add_3011_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n37159), 
            .O(n6582)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_6 (.CI(n37159), .I0(n1172), .I1(n96), .CO(n37160));
    SB_LUT4 add_3011_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n37158), 
            .O(n6583)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_5 (.CI(n37158), .I0(n1173), .I1(n97), .CO(n37159));
    SB_LUT4 add_3011_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n37157), 
            .O(n6584)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_4 (.CI(n37157), .I0(n1174), .I1(n98), .CO(n37158));
    SB_LUT4 add_3011_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n37156), 
            .O(n6585)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32978_3_lut (.I0(n48491), .I1(n90), .I2(n31_adj_4226), .I3(GND_net), 
            .O(n48492));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32978_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3011_3 (.CI(n37156), .I0(n1175), .I1(n99), .CO(n37157));
    SB_LUT4 add_3011_2_lut (.I0(GND_net), .I1(n375), .I2(n558), .I3(VCC_net), 
            .O(n6586)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_2 (.CI(VCC_net), .I0(n375), .I1(n558), .CO(n37156));
    SB_IO PIN_2_pad (.PACKAGE_PIN(PIN_2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_2_c_4)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_2_pad.PIN_TYPE = 6'b011001;
    defparam PIN_2_pad.PULLUP = 1'b0;
    defparam PIN_2_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_3975));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22609_3_lut (.I0(n648), .I1(n98), .I2(n4), .I3(GND_net), 
            .O(n6));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22609_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_12_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_3956), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n372));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22593_2_lut (.I0(n371), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22593_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_12_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_481_i42_4_lut (.I0(n372), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32833_3_lut (.I0(n42), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n48347));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32833_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i32834_3_lut (.I0(n48347), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n48348));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32834_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1440 (.I0(n48348), .I1(n22582), .I2(n96), .I3(n43351), 
            .O(n806));
    defparam i1_4_lut_adj_1440.LUT_INIT = 16'hefce;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_3976));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22569_2_lut (.I0(n370), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3954));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22569_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_12_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n371));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32854_3_lut (.I0(n48492), .I1(n89), .I2(n33_adj_4227), .I3(GND_net), 
            .O(n48368));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32854_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32781_4_lut (.I0(n43_adj_4233), .I1(n41_adj_4232), .I2(n39_adj_4230), 
            .I3(n47214), .O(n48295));
    defparam i32781_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33003_4_lut (.I0(n47542), .I1(n48239), .I2(n45_adj_4234), 
            .I3(n47203), .O(n48517));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33003_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32026_3_lut (.I0(n48368), .I1(n88), .I2(n35_adj_4228), .I3(GND_net), 
            .O(n47540));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32026_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10985_3_lut (.I0(encoder1_position[4]), .I1(n2262), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24403));   // quad.v(35[10] 41[6])
    defparam i10985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i547_4_lut_4_lut (.I0(n806), .I1(n96), .I2(n8_adj_4073), 
            .I3(n43351), .O(n914));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i547_4_lut_4_lut.LUT_INIT = 16'h14eb;
    SB_LUT4 i33005_4_lut (.I0(n47540), .I1(n48517), .I2(n45_adj_4234), 
            .I3(n48295), .O(n48519));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33005_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1441 (.I0(n48519), .I1(n22624), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1441.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_23_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[13]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_25[13]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i548_4_lut_4_lut (.I0(n806), .I1(n97), .I2(n6_adj_4074), 
            .I3(n783), .O(n915));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i548_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_12_LessThan_390_i44_4_lut (.I0(n371), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32685_3_lut (.I0(n44), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n48199));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32685_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 mux_23_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[14]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_25[14]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i636_3_lut_3_lut (.I0(n938), .I1(n5828), .I2(n916), 
            .I3(GND_net), .O(n1045));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i636_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1442 (.I0(n48199), .I1(n22579), .I2(n97), .I3(n43349), 
            .O(n671));
    defparam i1_4_lut_adj_1442.LUT_INIT = 16'hefce;
    SB_LUT4 add_2986_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n36777), 
            .O(n5826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i637_3_lut_3_lut (.I0(n938), .I1(n5829), .I2(n917), 
            .I3(GND_net), .O(n1046));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i637_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10988_3_lut (.I0(encoder1_position[7]), .I1(n2259), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24406));   // quad.v(35[10] 41[6])
    defparam i10988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[15]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_3977));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_22_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_25[15]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2986_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n36776), 
            .O(n5827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_6 (.CI(n36776), .I0(n915), .I1(n96), .CO(n36777));
    SB_LUT4 add_2986_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n36775), 
            .O(n5828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_5 (.CI(n36775), .I0(n916), .I1(n97), .CO(n36776));
    SB_LUT4 div_12_i638_3_lut_3_lut (.I0(n938), .I1(n5830), .I2(n918), 
            .I3(GND_net), .O(n1047));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i638_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2986_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n36774), 
            .O(n5829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_4 (.CI(n36774), .I0(n917), .I1(n98), .CO(n36775));
    SB_LUT4 add_2986_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n36773), 
            .O(n5830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_3 (.CI(n36773), .I0(n918), .I1(n99), .CO(n36774));
    SB_LUT4 add_2986_2_lut (.I0(GND_net), .I1(n373), .I2(n558), .I3(VCC_net), 
            .O(n5831)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_2 (.CI(VCC_net), .I0(n373), .I1(n558), .CO(n36773));
    SB_LUT4 div_12_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_3957), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n370));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22553_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3955));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22553_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_12_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_297_i46_4_lut (.I0(n370), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_4_lut_adj_1443 (.I0(n46), .I1(n22576), .I2(n98), .I3(n43347), 
            .O(n533));
    defparam i1_4_lut_adj_1443.LUT_INIT = 16'hefce;
    SB_LUT4 i1_4_lut_adj_1444 (.I0(n224), .I1(n99), .I2(n22573), .I3(n558), 
            .O(n5_adj_4363));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i1_4_lut_adj_1444.LUT_INIT = 16'h555d;
    SB_LUT4 div_12_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_23_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[16]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31371_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n46540));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31371_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 mux_22_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_25[16]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i639_3_lut_3_lut (.I0(n938), .I1(n5831), .I2(n373), 
            .I3(GND_net), .O(n1048));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i639_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i634_3_lut_3_lut (.I0(n938), .I1(n5826), .I2(n914), 
            .I3(GND_net), .O(n1043));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i634_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_23_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[17]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_12_i635_3_lut_3_lut (.I0(n938), .I1(n5827), .I2(n915), 
            .I3(GND_net), .O(n1044));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i635_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_22_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_25[17]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_1[23]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_1[22]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_LUT4 div_12_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4076));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_1[21]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_1[20]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_1[19]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_1[18]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_1[17]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_1[16]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_1[15]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_1[14]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_1[13]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_1[12]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_1[11]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_1[10]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_1[9]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_1[8]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_1[7]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_1[6]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_1[5]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_1[4]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_1[3]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_1[2]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_1[1]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_LUT4 i2_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n22573), .O(n248));
    defparam i2_4_lut.LUT_INIT = 16'hff37;
    SB_LUT4 i1_4_lut_adj_1445 (.I0(n46540), .I1(n22573), .I2(n99), .I3(n5_adj_4363), 
            .O(n392));
    defparam i1_4_lut_adj_1445.LUT_INIT = 16'hefce;
    SB_LUT4 i33816_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n49328));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33816_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_3979));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_3992));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n22633));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1446 (.I0(n81), .I1(n22627), .I2(GND_net), .I3(GND_net), 
            .O(n22624));
    defparam i1_2_lut_adj_1446.LUT_INIT = 16'hdddd;
    SB_LUT4 i10896_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24314));   // verilog/coms.v(125[12] 284[6])
    defparam i10896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10897_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24315));   // verilog/coms.v(125[12] 284[6])
    defparam i10897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31374_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n46887));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31374_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4078));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31368_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n46881));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31368_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_i1595_3_lut_3_lut (.I0(n2381), .I1(n6927), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10898_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24316));   // verilog/coms.v(125[12] 284[6])
    defparam i10898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_IO PIN_1_pad (.PACKAGE_PIN(PIN_1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_1_c_5)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_1_pad.PIN_TYPE = 6'b011001;
    defparam PIN_1_pad.PULLUP = 1'b0;
    defparam PIN_1_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_12_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4049), .I3(n37553), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_12_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4050), .I3(n37552), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_24 (.CI(n37552), .I0(GND_net), .I1(n3_adj_4050), 
            .CO(n37553));
    SB_LUT4 div_12_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4051), .I3(n37551), .O(n4_adj_3957)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_23 (.CI(n37551), .I0(GND_net), .I1(n4_adj_4051), 
            .CO(n37552));
    SB_LUT4 div_12_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4052), .I3(n37550), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_22 (.CI(n37550), .I0(GND_net), .I1(n5_adj_4052), 
            .CO(n37551));
    SB_LUT4 div_12_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4053), .I3(n37549), .O(n6_adj_3956)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_21 (.CI(n37549), .I0(GND_net), .I1(n6_adj_4053), 
            .CO(n37550));
    SB_LUT4 div_12_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4054), .I3(n37548), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10899_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24317));   // verilog/coms.v(125[12] 284[6])
    defparam i10899_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_12_unary_minus_2_add_3_20 (.CI(n37548), .I0(GND_net), .I1(n7_adj_4054), 
            .CO(n37549));
    SB_LUT4 div_12_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4055), .I3(n37547), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_19 (.CI(n37547), .I0(GND_net), .I1(n8_adj_4055), 
            .CO(n37548));
    SB_LUT4 div_12_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4056), .I3(n37546), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_18 (.CI(n37546), .I0(GND_net), .I1(n9_adj_4056), 
            .CO(n37547));
    SB_LUT4 div_12_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4057), .I3(n37545), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_17 (.CI(n37545), .I0(GND_net), .I1(n10_adj_4057), 
            .CO(n37546));
    SB_LUT4 div_12_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4058), .I3(n37544), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_16 (.CI(n37544), .I0(GND_net), .I1(n11_adj_4058), 
            .CO(n37545));
    SB_LUT4 div_12_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4059), .I3(n37543), .O(n12)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_15 (.CI(n37543), .I0(GND_net), .I1(n12_adj_4059), 
            .CO(n37544));
    SB_LUT4 div_12_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4060), .I3(n37542), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_14 (.CI(n37542), .I0(GND_net), .I1(n13_adj_4060), 
            .CO(n37543));
    SB_LUT4 div_12_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4061), .I3(n37541), .O(n14)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_13 (.CI(n37541), .I0(GND_net), .I1(n14_adj_4061), 
            .CO(n37542));
    SB_LUT4 div_12_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4062), .I3(n37540), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_12 (.CI(n37540), .I0(GND_net), .I1(n15_adj_4062), 
            .CO(n37541));
    SB_LUT4 div_12_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4063), .I3(n37539), .O(n16)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_11 (.CI(n37539), .I0(GND_net), .I1(n16_adj_4063), 
            .CO(n37540));
    SB_LUT4 div_12_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4064), .I3(n37538), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_10 (.CI(n37538), .I0(GND_net), .I1(n17_adj_4064), 
            .CO(n37539));
    SB_LUT4 div_12_i1583_3_lut_3_lut (.I0(n2381), .I1(n6915), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4065), .I3(n37537), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_9 (.CI(n37537), .I0(GND_net), .I1(n18_adj_4065), 
            .CO(n37538));
    SB_LUT4 div_12_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4066), .I3(n37536), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_8 (.CI(n37536), .I0(GND_net), .I1(n19_adj_4066), 
            .CO(n37537));
    SB_LUT4 div_12_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4067), .I3(n37535), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_7 (.CI(n37535), .I0(GND_net), .I1(n20_adj_4067), 
            .CO(n37536));
    SB_LUT4 div_12_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4068), .I3(n37534), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_6 (.CI(n37534), .I0(GND_net), .I1(n21_adj_4068), 
            .CO(n37535));
    SB_LUT4 div_12_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4069), .I3(n37533), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_5 (.CI(n37533), .I0(GND_net), .I1(n22_adj_4069), 
            .CO(n37534));
    SB_LUT4 div_12_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4070), .I3(n37532), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_4 (.CI(n37532), .I0(GND_net), .I1(n23_adj_4070), 
            .CO(n37533));
    SB_LUT4 div_12_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4071), .I3(n37531), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_3 (.CI(n37531), .I0(GND_net), .I1(n24_adj_4071), 
            .CO(n37532));
    SB_LUT4 div_12_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4072), .I3(VCC_net), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4072), 
            .CO(n37531));
    SB_LUT4 div_12_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4025), .I3(n37530), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_12_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4026), .I3(n37529), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_24 (.CI(n37529), .I0(GND_net), .I1(n3_adj_4026), 
            .CO(n37530));
    SB_LUT4 div_12_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4027), .I3(n37528), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_23 (.CI(n37528), .I0(GND_net), .I1(n4_adj_4027), 
            .CO(n37529));
    SB_LUT4 div_12_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4028), .I3(n37527), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_22 (.CI(n37527), .I0(GND_net), .I1(n5_adj_4028), 
            .CO(n37528));
    SB_LUT4 div_12_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4029), .I3(n37526), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_21 (.CI(n37526), .I0(GND_net), .I1(n6_adj_4029), 
            .CO(n37527));
    SB_LUT4 div_12_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4030), .I3(n37525), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_20 (.CI(n37525), .I0(GND_net), .I1(n7_adj_4030), 
            .CO(n37526));
    SB_LUT4 div_12_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4031), .I3(n37524), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_19 (.CI(n37524), .I0(GND_net), .I1(n8_adj_4031), 
            .CO(n37525));
    SB_LUT4 div_12_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4032), .I3(n37523), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_18 (.CI(n37523), .I0(GND_net), .I1(n9_adj_4032), 
            .CO(n37524));
    SB_LUT4 div_12_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4033), .I3(n37522), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_17 (.CI(n37522), .I0(GND_net), .I1(n10_adj_4033), 
            .CO(n37523));
    SB_LUT4 div_12_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4034), .I3(n37521), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_23_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b000001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY div_12_unary_minus_4_add_3_16 (.CI(n37521), .I0(GND_net), .I1(n11_adj_4034), 
            .CO(n37522));
    SB_LUT4 div_12_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4035), .I3(n37520), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_15 (.CI(n37520), .I0(GND_net), .I1(n12_adj_4035), 
            .CO(n37521));
    SB_LUT4 div_12_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4036), .I3(n37519), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_14 (.CI(n37519), .I0(GND_net), .I1(n13_adj_4036), 
            .CO(n37520));
    SB_LUT4 div_12_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4037), .I3(n37518), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_13 (.CI(n37518), .I0(GND_net), .I1(n14_adj_4037), 
            .CO(n37519));
    SB_LUT4 div_12_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4038), .I3(n37517), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_12 (.CI(n37517), .I0(GND_net), .I1(n15_adj_4038), 
            .CO(n37518));
    SB_LUT4 div_12_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4039), .I3(n37516), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_11 (.CI(n37516), .I0(GND_net), .I1(n16_adj_4039), 
            .CO(n37517));
    SB_LUT4 div_12_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4040), .I3(n37515), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1584_3_lut_3_lut (.I0(n2381), .I1(n6916), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_12_unary_minus_4_add_3_10 (.CI(n37515), .I0(GND_net), .I1(n17_adj_4040), 
            .CO(n37516));
    SB_LUT4 div_12_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4041), .I3(n37514), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_9 (.CI(n37514), .I0(GND_net), .I1(n18_adj_4041), 
            .CO(n37515));
    SB_LUT4 div_12_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4042), .I3(n37513), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_8 (.CI(n37513), .I0(GND_net), .I1(n19_adj_4042), 
            .CO(n37514));
    SB_LUT4 div_12_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4043), .I3(n37512), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_7 (.CI(n37512), .I0(GND_net), .I1(n20_adj_4043), 
            .CO(n37513));
    SB_LUT4 div_12_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4044), .I3(n37511), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_6 (.CI(n37511), .I0(GND_net), .I1(n21_adj_4044), 
            .CO(n37512));
    SB_LUT4 div_12_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4045), .I3(n37510), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_5 (.CI(n37510), .I0(GND_net), .I1(n22_adj_4045), 
            .CO(n37511));
    SB_LUT4 div_12_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4046), .I3(n37509), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_4 (.CI(n37509), .I0(GND_net), .I1(n23_adj_4046), 
            .CO(n37510));
    SB_LUT4 div_12_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4047), .I3(n37508), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_3 (.CI(n37508), .I0(GND_net), .I1(n24_adj_4047), 
            .CO(n37509));
    SB_LUT4 div_12_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4048), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4048), 
            .CO(n37508));
    SB_LUT4 div_12_i1773_3_lut_3_lut (.I0(n2642), .I1(n7000), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1587_3_lut_3_lut (.I0(n2381), .I1(n6919), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1588_3_lut_3_lut (.I0(n2381), .I1(n6920), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1774_3_lut_3_lut (.I0(n2642), .I1(n7001), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4209));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2999_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n36941), 
            .O(n6218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1482_i43_2_lut (.I0(n2266_adj_3996), .I1(n85), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4212));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2999_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n36940), 
            .O(n6219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_7 (.CI(n36940), .I0(n1044), .I1(n95), .CO(n36941));
    SB_LUT4 add_2999_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n36939), 
            .O(n6220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_6 (.CI(n36939), .I0(n1045), .I1(n96), .CO(n36940));
    SB_LUT4 add_2999_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n36938), 
            .O(n6221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_5 (.CI(n36938), .I0(n1046), .I1(n97), .CO(n36939));
    SB_LUT4 div_12_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4211));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2999_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n36937), 
            .O(n6222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10866_4_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n5023), .I3(n22498), .O(n24284));   // verilog/coms.v(125[12] 284[6])
    defparam i10866_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY add_2999_4 (.CI(n36937), .I0(n1047), .I1(n98), .CO(n36938));
    SB_LUT4 div_12_i1585_3_lut_3_lut (.I0(n2381), .I1(n6917), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2999_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n36936), 
            .O(n6223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_3 (.CI(n36936), .I0(n1048), .I1(n99), .CO(n36937));
    SB_LUT4 add_2999_2_lut (.I0(GND_net), .I1(n374), .I2(n558), .I3(VCC_net), 
            .O(n6224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4210));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2999_2 (.CI(VCC_net), .I0(n374), .I1(n558), .CO(n36936));
    SB_LUT4 div_12_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n385));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_556_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(pwm[3]), 
            .I2(pwm[2]), .I3(GND_net), .O(n6_adj_4012));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_556_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_12_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4206));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4207));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10872_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24290));   // verilog/coms.v(125[12] 284[6])
    defparam i10872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4208));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10873_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24291));   // verilog/coms.v(125[12] 284[6])
    defparam i10873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31430_3_lut_4_lut (.I0(pwm_count[3]), .I1(pwm[3]), .I2(pwm[2]), 
            .I3(pwm_count[2]), .O(n46943));   // verilog/motorControl.v(58[19:32])
    defparam i31430_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_12_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4203));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1586_3_lut_3_lut (.I0(n2381), .I1(n6918), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_1[0]));   // verilog/TinyFPGA_B.v(170[10] 172[6])
    SB_LUT4 div_12_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4205));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10874_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24292));   // verilog/coms.v(125[12] 284[6])
    defparam i10874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10875_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24293));   // verilog/coms.v(125[12] 284[6])
    defparam i10875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4197));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4199));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i808_3_lut_3_lut (.I0(n1193), .I1(n6585), .I2(n1175), 
            .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i808_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i807_3_lut_3_lut (.I0(n1193), .I1(n6584), .I2(n1174), 
            .I3(GND_net), .O(n1297));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i807_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10876_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24294));   // verilog/coms.v(125[12] 284[6])
    defparam i10876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i809_3_lut_3_lut (.I0(n1193), .I1(n6586), .I2(n375), 
            .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i809_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10877_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24295));   // verilog/coms.v(125[12] 284[6])
    defparam i10877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1447 (.I0(n84), .I1(n22618), .I2(GND_net), .I3(GND_net), 
            .O(n22615));
    defparam i1_2_lut_adj_1447.LUT_INIT = 16'hdddd;
    SB_LUT4 i10878_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24296));   // verilog/coms.v(125[12] 284[6])
    defparam i10878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4201));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4202));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10879_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24297));   // verilog/coms.v(125[12] 284[6])
    defparam i10879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i805_3_lut_3_lut (.I0(n1193), .I1(n6582), .I2(n1172), 
            .I3(GND_net), .O(n1295));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i805_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1601_3_lut_3_lut (.I0(n2381), .I1(n6933), .I2(n386), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10880_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24298));   // verilog/coms.v(125[12] 284[6])
    defparam i10880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4195));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31771_4_lut (.I0(n23_adj_4201), .I1(n21_adj_4199), .I2(n19_adj_4197), 
            .I3(n17_adj_4195), .O(n47285));
    defparam i31771_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i10881_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24299));   // verilog/coms.v(125[12] 284[6])
    defparam i10881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31761_4_lut (.I0(n29_adj_4205), .I1(n27_adj_4203), .I2(n25_adj_4202), 
            .I3(n47285), .O(n47275));
    defparam i31761_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32791_4_lut (.I0(n35_adj_4208), .I1(n33_adj_4207), .I2(n31_adj_4206), 
            .I3(n47275), .O(n48305));
    defparam i32791_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_12_LessThan_1482_i16_4_lut (.I0(n385), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_4194));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i10882_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24300));   // verilog/coms.v(125[12] 284[6])
    defparam i10882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i804_3_lut_3_lut (.I0(n1193), .I1(n6581), .I2(n1171), 
            .I3(GND_net), .O(n1294));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i804_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10883_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24301));   // verilog/coms.v(125[12] 284[6])
    defparam i10883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32629_3_lut (.I0(n16_adj_4194), .I1(n87), .I2(n39_adj_4210), 
            .I3(GND_net), .O(n48143));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32629_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32630_3_lut (.I0(n48143), .I1(n86), .I2(n41_adj_4211), .I3(GND_net), 
            .O(n48144));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32630_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i806_3_lut_3_lut (.I0(n1193), .I1(n6583), .I2(n1173), 
            .I3(GND_net), .O(n1296));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i806_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32323_4_lut (.I0(n41_adj_4211), .I1(n39_adj_4210), .I2(n27_adj_4203), 
            .I3(n47281), .O(n47837));
    defparam i32323_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_12_i803_3_lut_3_lut (.I0(n1193), .I1(n6580), .I2(n1170), 
            .I3(GND_net), .O(n1293));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i803_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32723_3_lut (.I0(n22_adj_4200), .I1(n93), .I2(n27_adj_4203), 
            .I3(GND_net), .O(n48237));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32723_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10884_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24302));   // verilog/coms.v(125[12] 284[6])
    defparam i10884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32018_3_lut (.I0(n48144), .I1(n85), .I2(n43_adj_4212), .I3(GND_net), 
            .O(n47532));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32018_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i802_3_lut_3_lut (.I0(n1193), .I1(n6579), .I2(n1169), 
            .I3(GND_net), .O(n1292));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i802_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10885_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24303));   // verilog/coms.v(125[12] 284[6])
    defparam i10885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4081));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1597_3_lut_3_lut (.I0(n2381), .I1(n6929), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1482_i28_3_lut (.I0(n20_adj_4198), .I1(n91), 
            .I2(n31_adj_4206), .I3(GND_net), .O(n28_adj_4204));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10886_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24304));   // verilog/coms.v(125[12] 284[6])
    defparam i10886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32975_4_lut (.I0(n28_adj_4204), .I1(n18_adj_4196), .I2(n31_adj_4206), 
            .I3(n47268), .O(n48489));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32975_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i10887_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24305));   // verilog/coms.v(125[12] 284[6])
    defparam i10887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31360_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n46873));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31360_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i32976_3_lut (.I0(n48489), .I1(n90), .I2(n33_adj_4207), .I3(GND_net), 
            .O(n48490));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32976_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32860_3_lut (.I0(n48490), .I1(n89), .I2(n35_adj_4208), .I3(GND_net), 
            .O(n48374));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32860_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32327_4_lut (.I0(n41_adj_4211), .I1(n39_adj_4210), .I2(n37_adj_4209), 
            .I3(n48305), .O(n47841));
    defparam i32327_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_12_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10888_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24306));   // verilog/coms.v(125[12] 284[6])
    defparam i10888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i889_3_lut_3_lut (.I0(n1316), .I1(n6656), .I2(n1298), 
            .I3(GND_net), .O(n1418));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i889_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i890_3_lut_3_lut (.I0(n1316), .I1(n6657), .I2(n1299), 
            .I3(GND_net), .O(n1419));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i890_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32857_4_lut (.I0(n47532), .I1(n48237), .I2(n43_adj_4212), 
            .I3(n47837), .O(n48371));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32857_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32016_3_lut (.I0(n48374), .I1(n88), .I2(n37_adj_4209), .I3(GND_net), 
            .O(n47530));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32016_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33043_4_lut (.I0(n47530), .I1(n48371), .I2(n43_adj_4212), 
            .I3(n47841), .O(n48557));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33043_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10989_3_lut (.I0(encoder1_position[8]), .I1(n2258), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24407));   // quad.v(35[10] 41[6])
    defparam i10989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33044_3_lut (.I0(n48557), .I1(n84), .I2(n2265_adj_3995), 
            .I3(GND_net), .O(n48558));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33044_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1448 (.I0(n48558), .I1(n22621), .I2(n83), .I3(n2264_adj_3994), 
            .O(n2288));
    defparam i1_4_lut_adj_1448.LUT_INIT = 16'hceef;
    SB_LUT4 i1_2_lut_adj_1449 (.I0(n87), .I1(n22609), .I2(GND_net), .I3(GND_net), 
            .O(n22606));
    defparam i1_2_lut_adj_1449.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_i891_3_lut_3_lut (.I0(n1316), .I1(n6658), .I2(n376), 
            .I3(GND_net), .O(n1420));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i891_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10990_3_lut (.I0(encoder1_position[9]), .I1(n2257), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24408));   // quad.v(35[10] 41[6])
    defparam i10990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1598_3_lut_3_lut (.I0(n2381), .I1(n6930), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10991_3_lut (.I0(encoder1_position[10]), .I1(n2256), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24409));   // quad.v(35[10] 41[6])
    defparam i10991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4190));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1594_3_lut_3_lut (.I0(n2381), .I1(n6926), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i887_3_lut_3_lut (.I0(n1316), .I1(n6654), .I2(n1296), 
            .I3(GND_net), .O(n1416));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i887_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10992_3_lut (.I0(encoder1_position[11]), .I1(n2255), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24410));   // quad.v(35[10] 41[6])
    defparam i10992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10993_3_lut (.I0(encoder1_position[12]), .I1(n2254), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24411));   // quad.v(35[10] 41[6])
    defparam i10993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10994_3_lut (.I0(encoder1_position[13]), .I1(n2253), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24412));   // quad.v(35[10] 41[6])
    defparam i10994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_91[23]), 
            .I2(n3_adj_3992), .I3(n36693), .O(displacement_23__N_1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_91[22]), 
            .I2(n3_adj_3992), .I3(n36692), .O(displacement_23__N_1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4193));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10995_3_lut (.I0(encoder1_position[14]), .I1(n2252), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24413));   // quad.v(35[10] 41[6])
    defparam i10995_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n36692), .I0(displacement_23__N_91[22]), 
            .I1(n3_adj_3992), .CO(n36693));
    SB_LUT4 div_12_i886_3_lut_3_lut (.I0(n1316), .I1(n6653), .I2(n1295), 
            .I3(GND_net), .O(n1415));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i886_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_91[21]), 
            .I2(n3_adj_3992), .I3(n36691), .O(displacement_23__N_1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n36691), .I0(displacement_23__N_91[21]), 
            .I1(n3_adj_3992), .CO(n36692));
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_91[20]), 
            .I2(n3_adj_3992), .I3(n36690), .O(displacement_23__N_1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10996_3_lut (.I0(encoder1_position[15]), .I1(n2251), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24414));   // quad.v(35[10] 41[6])
    defparam i10996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1593_3_lut_3_lut (.I0(n2381), .I1(n6925), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4192));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4191));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10997_3_lut (.I0(encoder1_position[16]), .I1(n2250), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24415));   // quad.v(35[10] 41[6])
    defparam i10997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10998_3_lut (.I0(encoder1_position[17]), .I1(n2249), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24416));   // quad.v(35[10] 41[6])
    defparam i10998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i888_3_lut_3_lut (.I0(n1316), .I1(n6655), .I2(n1297), 
            .I3(GND_net), .O(n1417));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i888_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i885_3_lut_3_lut (.I0(n1316), .I1(n6652), .I2(n1294), 
            .I3(GND_net), .O(n1414));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i885_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10999_3_lut (.I0(encoder1_position[18]), .I1(n2248), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24417));   // quad.v(35[10] 41[6])
    defparam i10999_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 div_12_i1592_3_lut_3_lut (.I0(n2381), .I1(n6924), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i11000_3_lut (.I0(encoder1_position[19]), .I1(n2247), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24418));   // quad.v(35[10] 41[6])
    defparam i11000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n384));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11001_3_lut (.I0(encoder1_position[20]), .I1(n2246), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24419));   // quad.v(35[10] 41[6])
    defparam i11001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4187));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4188));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i883_3_lut_3_lut (.I0(n1316), .I1(n6650), .I2(n1292), 
            .I3(GND_net), .O(n1412));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i883_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4189));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11002_3_lut (.I0(encoder1_position[21]), .I1(n2245), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24420));   // quad.v(35[10] 41[6])
    defparam i11002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11003_3_lut (.I0(encoder1_position[22]), .I1(n2244), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24421));   // quad.v(35[10] 41[6])
    defparam i11003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11004_3_lut (.I0(encoder1_position[23]), .I1(n2243), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24422));   // quad.v(35[10] 41[6])
    defparam i11004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4184));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4186));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4183));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11005_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n44475), 
            .I3(GND_net), .O(n24423));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i884_3_lut_3_lut (.I0(n1316), .I1(n6651), .I2(n1293), 
            .I3(GND_net), .O(n1413));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i884_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33800_4_lut (.I0(r_SM_Main[2]), .I1(n46590), .I2(n46591), 
            .I3(r_SM_Main[1]), .O(n29023));
    defparam i33800_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i10473_2_lut (.I0(n28694), .I1(n23889), .I2(GND_net), .I3(GND_net), 
            .O(n23891));   // verilog/coms.v(125[12] 284[6])
    defparam i10473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4177));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4179));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4181));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11008_4_lut (.I0(pwm_23__N_2948), .I1(n470), .I2(PWMLimit[1]), 
            .I3(n387), .O(n24426));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11008_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4175));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31129_4_lut (.I0(n25_adj_4181), .I1(n23_adj_4179), .I2(n21_adj_4177), 
            .I3(n19_adj_4175), .O(n46641));
    defparam i31129_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31125_4_lut (.I0(n31_adj_4186), .I1(n29_adj_4184), .I2(n27_adj_4183), 
            .I3(n46641), .O(n46637));
    defparam i31125_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i11012_4_lut (.I0(pwm_23__N_2948), .I1(n469), .I2(PWMLimit[2]), 
            .I3(n387), .O(n24430));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11012_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i32597_4_lut (.I0(n37_adj_4189), .I1(n35_adj_4188), .I2(n33_adj_4187), 
            .I3(n46637), .O(n48111));
    defparam i32597_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11013_4_lut (.I0(pwm_23__N_2948), .I1(n468), .I2(PWMLimit[3]), 
            .I3(n387), .O(n24431));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11013_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i14768_3_lut (.I0(\PID_CONTROLLER.result [4]), .I1(n416), .I2(n421), 
            .I3(GND_net), .O(n28170));
    defparam i14768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1417_i18_4_lut (.I0(n384), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4174));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i31317_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n46829));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31317_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i14826_3_lut (.I0(\PID_CONTROLLER.result [5]), .I1(n415), .I2(n421), 
            .I3(GND_net), .O(n28227));
    defparam i14826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32633_3_lut (.I0(n18_adj_4174), .I1(n87), .I2(n41_adj_4191), 
            .I3(GND_net), .O(n48147));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32633_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32634_3_lut (.I0(n48147), .I1(n86), .I2(n43_adj_4192), .I3(GND_net), 
            .O(n48148));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32634_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1591_3_lut_3_lut (.I0(n2381), .I1(n6923), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32351_4_lut (.I0(n43_adj_4192), .I1(n41_adj_4191), .I2(n29_adj_4184), 
            .I3(n46639), .O(n47865));
    defparam i32351_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_12_i1590_3_lut_3_lut (.I0(n2381), .I1(n6922), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1417_i26_3_lut (.I0(n24_adj_4180), .I1(n93), 
            .I2(n29_adj_4184), .I3(GND_net), .O(n26_adj_4182));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32010_3_lut (.I0(n48148), .I1(n85), .I2(n45_adj_4193), .I3(GND_net), 
            .O(n47524));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32010_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i11016_4_lut (.I0(pwm_23__N_2948), .I1(n465), .I2(PWMLimit[6]), 
            .I3(n387), .O(n24434));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11016_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4083));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i5_3_lut (.I0(\PID_CONTROLLER.result [7]), .I1(n413), .I2(n421), 
            .I3(GND_net), .O(n1));
    defparam i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1417_i30_3_lut (.I0(n22_adj_4178), .I1(n91), 
            .I2(n33_adj_4187), .I3(GND_net), .O(n30_adj_4185));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33034_4_lut (.I0(n30_adj_4185), .I1(n20_adj_4176), .I2(n33_adj_4187), 
            .I3(n46635), .O(n48548));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33034_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33035_3_lut (.I0(n48548), .I1(n90), .I2(n35_adj_4188), .I3(GND_net), 
            .O(n48549));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33035_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i11018_4_lut (.I0(pwm_23__N_2948), .I1(n463), .I2(PWMLimit[8]), 
            .I3(n387), .O(n24436));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11018_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i11019_4_lut (.I0(pwm_23__N_2948), .I1(n462), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24437));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11019_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_i1596_3_lut_3_lut (.I0(n2381), .I1(n6928), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32960_3_lut (.I0(n48549), .I1(n89), .I2(n37_adj_4189), .I3(GND_net), 
            .O(n48474));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32960_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31809_4_lut (.I0(n43_adj_4192), .I1(n41_adj_4191), .I2(n39_adj_4190), 
            .I3(n48111), .O(n47323));
    defparam i31809_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i11020_4_lut (.I0(pwm_23__N_2948), .I1(n461), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24438));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11020_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i32721_4_lut (.I0(n47524), .I1(n26_adj_4182), .I2(n45_adj_4193), 
            .I3(n47865), .O(n48235));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32721_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32894_3_lut (.I0(n48474), .I1(n88), .I2(n39_adj_4190), .I3(GND_net), 
            .O(n48408));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32894_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33001_4_lut (.I0(n48408), .I1(n48235), .I2(n45_adj_4193), 
            .I3(n47323), .O(n48515));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33001_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1450 (.I0(n48515), .I1(n22618), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1450.LUT_INIT = 16'hceef;
    SB_LUT4 i11021_4_lut (.I0(pwm_23__N_2948), .I1(n460), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24439));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11021_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10986_3_lut (.I0(encoder1_position[5]), .I1(n2261), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24404));   // quad.v(35[10] 41[6])
    defparam i10986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10987_3_lut (.I0(encoder1_position[6]), .I1(n2260), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24405));   // quad.v(35[10] 41[6])
    defparam i10987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11022_4_lut (.I0(pwm_23__N_2948), .I1(n459), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24440));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11022_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i11023_4_lut (.I0(pwm_23__N_2948), .I1(n458), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24441));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11023_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i11024_4_lut (.I0(pwm_23__N_2948), .I1(n457), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24442));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11024_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i11025_4_lut (.I0(pwm_23__N_2948), .I1(n456), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24443));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11025_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i11026_4_lut (.I0(pwm_23__N_2948), .I1(n455), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24444));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11026_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4173));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1589_3_lut_3_lut (.I0(n2381), .I1(n6921), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4172));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1451 (.I0(pwm_23__N_2948), .I1(n46604), .I2(PWMLimit[9]), 
            .I3(n387), .O(n41480));   // verilog/motorControl.v(31[14] 52[8])
    defparam i1_4_lut_adj_1451.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4171));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4170));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11029_4_lut (.I0(pwm_23__N_2948), .I1(n46565), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24447));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11029_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n383));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11030_4_lut (.I0(pwm_23__N_2948), .I1(n46567), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24448));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11030_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4160));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4162));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11031_4_lut (.I0(pwm_23__N_2948), .I1(n46569), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24449));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11031_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4164));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11032_4_lut (.I0(pwm_23__N_2948), .I1(n46571), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24450));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11032_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4166));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4167));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4169));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11033_4_lut (.I0(pwm_23__N_2948), .I1(n46573), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24451));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11033_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1600_3_lut_3_lut (.I0(n2381), .I1(n6932), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4158));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11034_3_lut (.I0(quadA_debounced_adj_3982), .I1(reg_B_adj_4411[1]), 
            .I2(n44154), .I3(GND_net), .O(n24452));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11034_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31149_4_lut (.I0(n27_adj_4164), .I1(n25_adj_4162), .I2(n23_adj_4160), 
            .I3(n21_adj_4158), .O(n46661));
    defparam i31149_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31145_4_lut (.I0(n33_adj_4169), .I1(n31_adj_4167), .I2(n29_adj_4166), 
            .I3(n46661), .O(n46657));
    defparam i31145_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i11035_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_3980), 
            .I3(n22534), .O(n24453));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11035_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i7_2_lut (.I0(pwm_23__N_2951[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4004));   // verilog/motorControl.v(25[23:29])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_LessThan_1350_i20_4_lut (.I0(n383), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4157));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_LessThan_1350_i28_3_lut (.I0(n26_adj_4163), .I1(n93), 
            .I2(n31_adj_4167), .I3(GND_net), .O(n28_adj_4165));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i9_2_lut (.I0(deadband[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4001));   // verilog/motorControl.v(25[23:29])
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14_2_lut (.I0(deadband[4]), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4000));   // verilog/motorControl.v(25[23:29])
    defparam i14_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_LessThan_1350_i32_3_lut (.I0(n24_adj_4161), .I1(n91), 
            .I2(n35_adj_4170), .I3(GND_net), .O(n32_adj_4168));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33030_4_lut (.I0(n32_adj_4168), .I1(n22_adj_4159), .I2(n35_adj_4170), 
            .I3(n46655), .O(n48544));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33030_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33031_3_lut (.I0(n48544), .I1(n90), .I2(n37_adj_4171), .I3(GND_net), 
            .O(n48545));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33031_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32964_3_lut (.I0(n48545), .I1(n89), .I2(n39_adj_4172), .I3(GND_net), 
            .O(n48478));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32964_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32607_4_lut (.I0(n39_adj_4172), .I1(n37_adj_4171), .I2(n35_adj_4170), 
            .I3(n46657), .O(n48121));
    defparam i32607_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32913_4_lut (.I0(n28_adj_4165), .I1(n20_adj_4157), .I2(n31_adj_4167), 
            .I3(n46659), .O(n48427));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32913_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32890_3_lut (.I0(n48478), .I1(n88), .I2(n41_adj_4173), .I3(GND_net), 
            .O(n48404));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32890_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33032_4_lut (.I0(n48404), .I1(n48427), .I2(n41_adj_4173), 
            .I3(n48121), .O(n48546));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33032_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33033_3_lut (.I0(n48546), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n48547));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33033_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_12_i1599_3_lut_3_lut (.I0(n2381), .I1(n6931), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32962_3_lut (.I0(n48547), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n48476));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32962_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1452 (.I0(n48476), .I1(n22615), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1452.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4156));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4154));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4153));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4152));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n382));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4148));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4149));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4151));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4142));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4144));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4146));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4140));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31172_4_lut (.I0(n29_adj_4146), .I1(n27_adj_4144), .I2(n25_adj_4142), 
            .I3(n23_adj_4140), .O(n46684));
    defparam i31172_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31163_4_lut (.I0(n35_adj_4151), .I1(n33_adj_4149), .I2(n31_adj_4148), 
            .I3(n46684), .O(n46675));
    defparam i31163_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1281_i22_4_lut (.I0(n382), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4139));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_LessThan_1281_i30_3_lut (.I0(n28_adj_4145), .I1(n93), 
            .I2(n33_adj_4149), .I3(GND_net), .O(n30_adj_4147));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1281_i34_3_lut (.I0(n26_adj_4143), .I1(n91), 
            .I2(n37_adj_4152), .I3(GND_net), .O(n34_adj_4150));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33028_4_lut (.I0(n34_adj_4150), .I1(n24_adj_4141), .I2(n37_adj_4152), 
            .I3(n46673), .O(n48542));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33028_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33029_3_lut (.I0(n48542), .I1(n90), .I2(n39_adj_4153), .I3(GND_net), 
            .O(n48543));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33029_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32966_3_lut (.I0(n48543), .I1(n89), .I2(n41_adj_4154), .I3(GND_net), 
            .O(n48480));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32966_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32617_4_lut (.I0(n41_adj_4154), .I1(n39_adj_4153), .I2(n37_adj_4152), 
            .I3(n46675), .O(n48131));
    defparam i32617_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32591_4_lut (.I0(n30_adj_4147), .I1(n22_adj_4139), .I2(n33_adj_4149), 
            .I3(n46682), .O(n48105));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32591_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32888_3_lut (.I0(n48480), .I1(n88), .I2(n43_adj_4156), .I3(GND_net), 
            .O(n42_adj_4155));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32888_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32809_4_lut (.I0(n42_adj_4155), .I1(n48105), .I2(n43_adj_4156), 
            .I3(n48131), .O(n48323));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32809_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32810_3_lut (.I0(n48323), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n48324));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32810_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1453 (.I0(n48324), .I1(n22612), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1453.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i1763_3_lut_3_lut (.I0(n2642), .I1(n6990), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1210_i43_2_lut (.I0(n1864), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4136));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i45_2_lut (.I0(n1863), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4138));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i41_2_lut (.I0(n1865), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4135));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4134));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1649_3_lut_3_lut (.I0(n2471), .I1(n6943), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n381));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4130));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4131));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4133));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10_2_lut (.I0(pwm_23__N_2951[4]), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4002));   // verilog/motorControl.v(25[23:29])
    defparam i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i7_2_lut_adj_1454 (.I0(pwm_23__N_2951[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4003));   // verilog/motorControl.v(25[23:29])
    defparam i7_2_lut_adj_1454.LUT_INIT = 16'h6666;
    SB_LUT4 i8_2_lut (.I0(PWMLimit[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4007));   // verilog/motorControl.v(25[23:29])
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4124));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13_2_lut (.I0(PWMLimit[4]), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4005));   // verilog/motorControl.v(25[23:29])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4126));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i5_2_lut (.I0(PWMLimit[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4006));   // verilog/motorControl.v(25[23:29])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4128));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i970_3_lut_3_lut (.I0(n1436), .I1(n6698), .I2(n1420), 
            .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i970_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1642_3_lut_3_lut (.I0(n2471), .I1(n6936), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4122));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31198_4_lut (.I0(n31_adj_4128), .I1(n29_adj_4126), .I2(n27_adj_4124), 
            .I3(n25_adj_4122), .O(n46710));
    defparam i31198_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31190_4_lut (.I0(n37_adj_4133), .I1(n35_adj_4131), .I2(n33_adj_4130), 
            .I3(n46710), .O(n46702));
    defparam i31190_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1210_i24_4_lut (.I0(n381), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4121));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_i1643_3_lut_3_lut (.I0(n2471), .I1(n6937), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1210_i32_3_lut (.I0(n30_adj_4127), .I1(n93), 
            .I2(n35_adj_4131), .I3(GND_net), .O(n32_adj_4129));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i967_3_lut_3_lut (.I0(n1436), .I1(n6695), .I2(n1417), 
            .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i967_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1210_i36_3_lut (.I0(n28_adj_4125), .I1(n91), 
            .I2(n39_adj_4134), .I3(GND_net), .O(n36_adj_4132));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i968_3_lut_3_lut (.I0(n1436), .I1(n6696), .I2(n1418), 
            .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i968_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33026_4_lut (.I0(n36_adj_4132), .I1(n26_adj_4123), .I2(n39_adj_4134), 
            .I3(n46700), .O(n48540));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33026_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_12_i1644_3_lut_3_lut (.I0(n2471), .I1(n6938), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33027_3_lut (.I0(n48540), .I1(n90), .I2(n41_adj_4135), .I3(GND_net), 
            .O(n48541));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33027_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32968_3_lut (.I0(n48541), .I1(n89), .I2(n43_adj_4136), .I3(GND_net), 
            .O(n48482));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32968_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32627_4_lut (.I0(n43_adj_4136), .I1(n41_adj_4135), .I2(n39_adj_4134), 
            .I3(n46702), .O(n48141));
    defparam i32627_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32441_4_lut (.I0(n32_adj_4129), .I1(n24_adj_4121), .I2(n35_adj_4131), 
            .I3(n46706), .O(n47955));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32441_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32886_3_lut (.I0(n48482), .I1(n88), .I2(n45_adj_4138), .I3(GND_net), 
            .O(n44_adj_4137));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32886_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32443_4_lut (.I0(n44_adj_4137), .I1(n47955), .I2(n45_adj_4138), 
            .I3(n48141), .O(n47957));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32443_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1455 (.I0(n47957), .I1(n22609), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1455.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i1647_3_lut_3_lut (.I0(n2471), .I1(n6941), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1645_3_lut_3_lut (.I0(n2471), .I1(n6939), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4117));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i964_3_lut_3_lut (.I0(n1436), .I1(n6692), .I2(n1414), 
            .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i964_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4116));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1648_3_lut_3_lut (.I0(n2471), .I1(n6942), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n380));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4120));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4119));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1661_3_lut_3_lut (.I0(n2471), .I1(n6955), .I2(n387_adj_3993), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4112));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4114));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4115));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i963_3_lut_3_lut (.I0(n1436), .I1(n6691), .I2(n1413), 
            .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i963_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31239_4_lut (.I0(n33_adj_4115), .I1(n31_adj_4114), .I2(n29_adj_4112), 
            .I3(n27), .O(n46751));
    defparam i31239_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1137_i38_3_lut (.I0(n30_adj_4113), .I1(n91), 
            .I2(n41_adj_4120), .I3(GND_net), .O(n38_adj_4118));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1137_i26_4_lut (.I0(n380), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_i966_3_lut_3_lut (.I0(n1436), .I1(n6694), .I2(n1416), 
            .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i966_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32817_3_lut (.I0(n26), .I1(n95), .I2(n33_adj_4115), .I3(GND_net), 
            .O(n48331));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32817_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i971_3_lut_3_lut (.I0(n1436), .I1(n6699), .I2(n377), 
            .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i971_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32818_3_lut (.I0(n48331), .I1(n94), .I2(n35_adj_4116), .I3(GND_net), 
            .O(n48332));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32818_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31224_4_lut (.I0(n39_adj_4119), .I1(n37_adj_4117), .I2(n35_adj_4116), 
            .I3(n46751), .O(n46736));
    defparam i31224_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33024_4_lut (.I0(n38_adj_4118), .I1(n28_adj_4111), .I2(n41_adj_4120), 
            .I3(n46730), .O(n48538));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33024_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32706_3_lut (.I0(n48332), .I1(n93), .I2(n37_adj_4117), .I3(GND_net), 
            .O(n48220));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32706_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33110_4_lut (.I0(n48220), .I1(n48538), .I2(n41_adj_4120), 
            .I3(n46736), .O(n48624));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33110_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33111_3_lut (.I0(n48624), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n48625));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33111_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33083_3_lut (.I0(n48625), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n48597));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33083_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1456 (.I0(n48597), .I1(n22606), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1456.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i965_3_lut_3_lut (.I0(n1436), .I1(n6693), .I2(n1415), 
            .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i965_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4107));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i962_3_lut_3_lut (.I0(n1436), .I1(n6690), .I2(n1412), 
            .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i962_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4106));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10_2_lut_adj_1457 (.I0(n413), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4010));   // verilog/motorControl.v(25[23:29])
    defparam i10_2_lut_adj_1457.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_i1646_3_lut_3_lut (.I0(n2471), .I1(n6940), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n379));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4110));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4109));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4102));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4104));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1650_3_lut_3_lut (.I0(n2471), .I1(n6944), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1651_3_lut_3_lut (.I0(n2471), .I1(n6945), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4105));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11_2_lut (.I0(n416), .I1(\PID_CONTROLLER.result [4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4008));   // verilog/motorControl.v(25[23:29])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i6_2_lut (.I0(n415), .I1(\PID_CONTROLLER.result [5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4009));   // verilog/motorControl.v(25[23:29])
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31263_4_lut (.I0(n35_adj_4105), .I1(n33_adj_4104), .I2(n31_adj_4102), 
            .I3(n29), .O(n46775));
    defparam i31263_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_i1657_3_lut_3_lut (.I0(n2471), .I1(n6951), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1062_i40_3_lut (.I0(n32_adj_4103), .I1(n91), 
            .I2(n43_adj_4110), .I3(GND_net), .O(n40_adj_4108));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1062_i28_4_lut (.I0(n379), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32821_3_lut (.I0(n28), .I1(n95), .I2(n35_adj_4105), .I3(GND_net), 
            .O(n48335));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32821_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32822_3_lut (.I0(n48335), .I1(n94), .I2(n37_adj_4106), .I3(GND_net), 
            .O(n48336));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32822_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31255_4_lut (.I0(n41_adj_4109), .I1(n39_adj_4107), .I2(n37_adj_4106), 
            .I3(n46775), .O(n46767));
    defparam i31255_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32819_4_lut (.I0(n40_adj_4108), .I1(n30_adj_4101), .I2(n43_adj_4110), 
            .I3(n46765), .O(n48333));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32819_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32702_3_lut (.I0(n48336), .I1(n93), .I2(n39_adj_4107), .I3(GND_net), 
            .O(n48216));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32702_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33057_4_lut (.I0(n48216), .I1(n48333), .I2(n43_adj_4110), 
            .I3(n46767), .O(n48571));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33057_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33058_3_lut (.I0(n48571), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n48572));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33058_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1458 (.I0(n48572), .I1(n22603), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1458.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i1658_3_lut_3_lut (.I0(n2471), .I1(n6952), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4097));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n378));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4096));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4100));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i969_3_lut_3_lut (.I0(n1436), .I1(n6697), .I2(n1419), 
            .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i969_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1659_3_lut_3_lut (.I0(n2471), .I1(n6953), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4099));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11036_4_lut (.I0(pwm_23__N_2948), .I1(n471), .I2(PWMLimit[0]), 
            .I3(n387), .O(n24454));   // verilog/motorControl.v(31[14] 52[8])
    defparam i11036_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4095));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31308_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n46820));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i31308_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11038_3_lut (.I0(setpoint[1]), .I1(n3801), .I2(n44107), .I3(GND_net), 
            .O(n24456));   // verilog/coms.v(125[12] 284[6])
    defparam i11038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31281_4_lut (.I0(n37_adj_4095), .I1(n35), .I2(n33), .I3(n31), 
            .O(n46793));
    defparam i31281_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i11039_3_lut (.I0(setpoint[2]), .I1(n3802), .I2(n44107), .I3(GND_net), 
            .O(n24457));   // verilog/coms.v(125[12] 284[6])
    defparam i11039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1654_3_lut_3_lut (.I0(n2471), .I1(n6948), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i11040_3_lut (.I0(setpoint[3]), .I1(n3803), .I2(n44107), .I3(GND_net), 
            .O(n24458));   // verilog/coms.v(125[12] 284[6])
    defparam i11040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4089));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i11041_3_lut (.I0(setpoint[4]), .I1(n3804), .I2(n44107), .I3(GND_net), 
            .O(n24459));   // verilog/coms.v(125[12] 284[6])
    defparam i11041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_985_i42_3_lut (.I0(n34_adj_4094), .I1(n91), 
            .I2(n45_adj_4100), .I3(GND_net), .O(n42_adj_4098));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_985_i30_4_lut (.I0(n378), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32879_3_lut (.I0(n30), .I1(n95), .I2(n37_adj_4095), .I3(GND_net), 
            .O(n48393));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32879_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1048_3_lut_3_lut (.I0(n1553), .I1(n6739), .I2(n1538), 
            .I3(GND_net), .O(n1652));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1048_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i11042_3_lut (.I0(setpoint[5]), .I1(n3805), .I2(n44107), .I3(GND_net), 
            .O(n24460));   // verilog/coms.v(125[12] 284[6])
    defparam i11042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32880_3_lut (.I0(n48393), .I1(n94), .I2(n39_adj_4096), .I3(GND_net), 
            .O(n48394));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32880_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31275_4_lut (.I0(n43_adj_4099), .I1(n41_adj_4097), .I2(n39_adj_4096), 
            .I3(n46793), .O(n46787));
    defparam i31275_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i11043_3_lut (.I0(setpoint[6]), .I1(n3806), .I2(n44107), .I3(GND_net), 
            .O(n24461));   // verilog/coms.v(125[12] 284[6])
    defparam i11043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32435_4_lut (.I0(n42_adj_4098), .I1(n32_adj_4093), .I2(n45_adj_4100), 
            .I3(n46783), .O(n47949));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32435_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32700_3_lut (.I0(n48394), .I1(n93), .I2(n41_adj_4097), .I3(GND_net), 
            .O(n48214));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32700_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1653_3_lut_3_lut (.I0(n2471), .I1(n6947), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32881_4_lut (.I0(n48214), .I1(n47949), .I2(n45_adj_4100), 
            .I3(n46787), .O(n48395));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32881_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11044_3_lut (.I0(setpoint[7]), .I1(n3807), .I2(n44107), .I3(GND_net), 
            .O(n24462));   // verilog/coms.v(125[12] 284[6])
    defparam i11044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1459 (.I0(n48395), .I1(n22600), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1459.LUT_INIT = 16'hceef;
    SB_LUT4 i11045_3_lut (.I0(setpoint[8]), .I1(n3808), .I2(n44107), .I3(GND_net), 
            .O(n24463));   // verilog/coms.v(125[12] 284[6])
    defparam i11045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11046_3_lut (.I0(setpoint[9]), .I1(n3809), .I2(n44107), .I3(GND_net), 
            .O(n24464));   // verilog/coms.v(125[12] 284[6])
    defparam i11046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4092));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1045_3_lut_3_lut (.I0(n1553), .I1(n6736), .I2(n1535), 
            .I3(GND_net), .O(n1649));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1045_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11047_3_lut (.I0(setpoint[10]), .I1(n3810), .I2(n44107), 
            .I3(GND_net), .O(n24465));   // verilog/coms.v(125[12] 284[6])
    defparam i11047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1046_3_lut_3_lut (.I0(n1553), .I1(n6737), .I2(n1536), 
            .I3(GND_net), .O(n1650));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1046_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4091));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11048_3_lut (.I0(setpoint[11]), .I1(n3811), .I2(n44107), 
            .I3(GND_net), .O(n24466));   // verilog/coms.v(125[12] 284[6])
    defparam i11048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10390_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n23808));   // verilog/coms.v(125[12] 284[6])
    defparam i10390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4090));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11049_3_lut (.I0(setpoint[12]), .I1(n3812), .I2(n44107), 
            .I3(GND_net), .O(n24467));   // verilog/coms.v(125[12] 284[6])
    defparam i11049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10394_3_lut (.I0(\PID_CONTROLLER.err_prev [0]), .I1(\PID_CONTROLLER.err [0]), 
            .I2(n44066), .I3(GND_net), .O(n23812));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10394_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29081_4_lut (.I0(n22512), .I1(n22525), .I2(n737), .I3(n2854), 
            .O(n44592));
    defparam i29081_4_lut.LUT_INIT = 16'hfac8;
    SB_LUT4 div_12_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n377));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1460 (.I0(n43773), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n44557), .I3(n20156), .O(n42006));   // verilog/coms.v(125[12] 284[6])
    defparam i1_4_lut_adj_1460.LUT_INIT = 16'hd5f5;
    SB_LUT4 i11050_3_lut (.I0(setpoint[13]), .I1(n3813), .I2(n44107), 
            .I3(GND_net), .O(n24468));   // verilog/coms.v(125[12] 284[6])
    defparam i11050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10396_3_lut (.I0(encoder0_position[0]), .I1(n2316), .I2(count_enable), 
            .I3(GND_net), .O(n23814));   // quad.v(35[10] 41[6])
    defparam i10396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10397_3_lut (.I0(encoder1_position[0]), .I1(n2266), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n23815));   // quad.v(35[10] 41[6])
    defparam i10397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10398_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n44475), 
            .I3(GND_net), .O(n23816));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11051_3_lut (.I0(setpoint[14]), .I1(n3814), .I2(n44107), 
            .I3(GND_net), .O(n24469));   // verilog/coms.v(125[12] 284[6])
    defparam i11051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_906_i32_4_lut (.I0(n377), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32825_3_lut (.I0(n32), .I1(n95), .I2(n39_adj_4090), .I3(GND_net), 
            .O(n48339));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32825_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10399_4_lut (.I0(r_SM_Main[2]), .I1(n1_adj_4351), .I2(n28989), 
            .I3(r_SM_Main[1]), .O(n23817));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10399_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i32826_3_lut (.I0(n48339), .I1(n94), .I2(n41_adj_4091), .I3(GND_net), 
            .O(n48340));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32826_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31949_4_lut (.I0(n41_adj_4091), .I1(n39_adj_4090), .I2(n37), 
            .I3(n46820), .O(n47463));
    defparam i31949_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32433_3_lut (.I0(n34_adj_4089), .I1(n96), .I2(n37), .I3(GND_net), 
            .O(n47947));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32433_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10403_3_lut (.I0(quadB_debounced_adj_3983), .I1(reg_B_adj_4411[0]), 
            .I2(n44154), .I3(GND_net), .O(n23821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1652_3_lut_3_lut (.I0(n2471), .I1(n6946), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i11052_3_lut (.I0(setpoint[15]), .I1(n3815), .I2(n44107), 
            .I3(GND_net), .O(n24470));   // verilog/coms.v(125[12] 284[6])
    defparam i11052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11053_3_lut (.I0(setpoint[16]), .I1(n3816), .I2(n44107), 
            .I3(GND_net), .O(n24471));   // verilog/coms.v(125[12] 284[6])
    defparam i11053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32696_3_lut (.I0(n48340), .I1(n93), .I2(n43_adj_4092), .I3(GND_net), 
            .O(n48210));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32696_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32823_4_lut (.I0(n48210), .I1(n47947), .I2(n43_adj_4092), 
            .I3(n47463), .O(n48337));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32823_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32824_3_lut (.I0(n48337), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n48338));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32824_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1461 (.I0(n48338), .I1(n22597), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1461.LUT_INIT = 16'hceef;
    SB_LUT4 i11054_3_lut (.I0(setpoint[17]), .I1(n3817), .I2(n44107), 
            .I3(GND_net), .O(n24472));   // verilog/coms.v(125[12] 284[6])
    defparam i11054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1042_3_lut_3_lut (.I0(n1553), .I1(n6733), .I2(n1532), 
            .I3(GND_net), .O(n1646));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1042_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1656_3_lut_3_lut (.I0(n2471), .I1(n6950), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10410_3_lut (.I0(setpoint[0]), .I1(n3800), .I2(n44107), .I3(GND_net), 
            .O(n23828));   // verilog/coms.v(125[12] 284[6])
    defparam i10410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11055_3_lut (.I0(setpoint[18]), .I1(n3818), .I2(n44107), 
            .I3(GND_net), .O(n24473));   // verilog/coms.v(125[12] 284[6])
    defparam i11055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_3971));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11056_3_lut (.I0(setpoint[19]), .I1(n3819), .I2(n44107), 
            .I3(GND_net), .O(n24474));   // verilog/coms.v(125[12] 284[6])
    defparam i11056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4088));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11057_3_lut (.I0(setpoint[20]), .I1(n3820), .I2(n44107), 
            .I3(GND_net), .O(n24475));   // verilog/coms.v(125[12] 284[6])
    defparam i11057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11058_3_lut (.I0(setpoint[21]), .I1(n3821), .I2(n44107), 
            .I3(GND_net), .O(n24476));   // verilog/coms.v(125[12] 284[6])
    defparam i11058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4086));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4085));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i11059_3_lut (.I0(setpoint[22]), .I1(n3822), .I2(n44107), 
            .I3(GND_net), .O(n24477));   // verilog/coms.v(125[12] 284[6])
    defparam i11059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1462 (.I0(n90), .I1(n22600), .I2(GND_net), .I3(GND_net), 
            .O(n22597));
    defparam i1_2_lut_adj_1462.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n376));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11060_3_lut (.I0(setpoint[23]), .I1(n3823), .I2(n44107), 
            .I3(GND_net), .O(n24478));   // verilog/coms.v(125[12] 284[6])
    defparam i11060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1655_3_lut_3_lut (.I0(n2471), .I1(n6949), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1660_3_lut_3_lut (.I0(n2471), .I1(n6954), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_825_i34_4_lut (.I0(n376), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_i1041_3_lut_3_lut (.I0(n1553), .I1(n6732), .I2(n1531), 
            .I3(GND_net), .O(n1645));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1041_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10464_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n28517), 
            .I3(n22539), .O(n23882));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10464_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i10465_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n28517), 
            .I3(n22534), .O(n23883));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10465_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 div_12_i1049_3_lut_3_lut (.I0(n1553), .I1(n6740), .I2(n378), 
            .I3(GND_net), .O(n1653));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1049_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32827_3_lut (.I0(n34), .I1(n95), .I2(n41_adj_4085), .I3(GND_net), 
            .O(n48341));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32827_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32828_3_lut (.I0(n48341), .I1(n94), .I2(n43_adj_4086), .I3(GND_net), 
            .O(n48342));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32828_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10466_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_3986), 
            .I3(n22539), .O(n23884));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10466_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31969_4_lut (.I0(n43_adj_4086), .I1(n41_adj_4085), .I2(n39), 
            .I3(n46829), .O(n47483));
    defparam i31969_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i10467_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_3986), 
            .I3(n22534), .O(n23885));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10467_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_12_LessThan_825_i38_3_lut (.I0(n36_adj_4083), .I1(n96), 
            .I2(n39), .I3(GND_net), .O(n38_adj_4084));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32694_3_lut (.I0(n48342), .I1(n93), .I2(n45_adj_4088), .I3(GND_net), 
            .O(n44_adj_4087));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32694_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32431_4_lut (.I0(n44_adj_4087), .I1(n38_adj_4084), .I2(n45_adj_4088), 
            .I3(n47483), .O(n47945));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32431_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1463 (.I0(n47945), .I1(n22594), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1463.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i725_3_lut_3_lut (.I0(n1067), .I1(n6224), .I2(n374), 
            .I3(GND_net), .O(n1175));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i725_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_3972));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10468_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_3981), 
            .I3(n22539), .O(n23886));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10468_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_12_i1044_3_lut_3_lut (.I0(n1553), .I1(n6735), .I2(n1534), 
            .I3(GND_net), .O(n1648));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1044_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10469_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_3981), 
            .I3(n22534), .O(n23887));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10469_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_12_i724_3_lut_3_lut (.I0(n1067), .I1(n6223), .I2(n1048), 
            .I3(GND_net), .O(n1174));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i724_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1043_3_lut_3_lut (.I0(n1553), .I1(n6734), .I2(n1533), 
            .I3(GND_net), .O(n1647));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1043_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_3973));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11064_4_lut (.I0(n28694), .I1(byte_transmit_counter[0]), .I2(n2241), 
            .I3(n3840), .O(n24482));   // verilog/coms.v(125[12] 284[6])
    defparam i11064_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10491_2_lut (.I0(n28694), .I1(n23907), .I2(GND_net), .I3(GND_net), 
            .O(n23909));   // verilog/coms.v(125[12] 284[6])
    defparam i10491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10488_2_lut (.I0(n28694), .I1(n23904), .I2(GND_net), .I3(GND_net), 
            .O(n23906));   // verilog/coms.v(125[12] 284[6])
    defparam i10488_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10485_2_lut (.I0(n28694), .I1(n23901), .I2(GND_net), .I3(GND_net), 
            .O(n23903));   // verilog/coms.v(125[12] 284[6])
    defparam i10485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10482_2_lut (.I0(n28694), .I1(n23898), .I2(GND_net), .I3(GND_net), 
            .O(n23900));   // verilog/coms.v(125[12] 284[6])
    defparam i10482_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1040_3_lut_3_lut (.I0(n1553), .I1(n6731), .I2(n1530), 
            .I3(GND_net), .O(n1644));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1040_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i722_3_lut_3_lut (.I0(n1067), .I1(n6221), .I2(n1046), 
            .I3(GND_net), .O(n1172));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i722_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1039_3_lut_3_lut (.I0(n1553), .I1(n6730), .I2(n1529), 
            .I3(GND_net), .O(n1643));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1039_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n375));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1047_3_lut_3_lut (.I0(n1553), .I1(n6738), .I2(n1537), 
            .I3(GND_net), .O(n1651));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1047_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1124_3_lut_3_lut (.I0(n1667), .I1(n6753), .I2(n1653), 
            .I3(GND_net), .O(n1764));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1124_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10463_4_lut (.I0(n23783), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n23649), .O(n23881));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10463_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_12_i1121_3_lut_3_lut (.I0(n1667), .I1(n6750), .I2(n1650), 
            .I3(GND_net), .O(n1761));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1121_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1122_3_lut_3_lut (.I0(n1667), .I1(n6751), .I2(n1651), 
            .I3(GND_net), .O(n1762));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1122_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i721_3_lut_3_lut (.I0(n1067), .I1(n6220), .I2(n1045), 
            .I3(GND_net), .O(n1171));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i721_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1118_3_lut_3_lut (.I0(n1667), .I1(n6747), .I2(n1647), 
            .I3(GND_net), .O(n1758));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1118_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i720_3_lut_3_lut (.I0(n1067), .I1(n6219), .I2(n1044), 
            .I3(GND_net), .O(n1170));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i720_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10460_4_lut (.I0(n23783), .I1(r_Bit_Index[2]), .I2(n4016), 
            .I3(n23649), .O(n23878));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10460_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_12_i1117_3_lut_3_lut (.I0(n1667), .I1(n6746), .I2(n1646), 
            .I3(GND_net), .O(n1757));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1117_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1125_3_lut_3_lut (.I0(n1667), .I1(n6754), .I2(n379), 
            .I3(GND_net), .O(n1765));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1125_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10457_4_lut (.I0(n23785), .I1(r_Bit_Index_adj_4404[1]), .I2(r_Bit_Index_adj_4404[0]), 
            .I3(n23655), .O(n23875));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10457_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_12_i1120_3_lut_3_lut (.I0(n1667), .I1(n6749), .I2(n1649), 
            .I3(GND_net), .O(n1760));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1120_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1119_3_lut_3_lut (.I0(n1667), .I1(n6748), .I2(n1648), 
            .I3(GND_net), .O(n1759));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1119_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1116_3_lut_3_lut (.I0(n1667), .I1(n6745), .I2(n1645), 
            .I3(GND_net), .O(n1756));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1116_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1114_3_lut_3_lut (.I0(n1667), .I1(n6743), .I2(n1643), 
            .I3(GND_net), .O(n1754));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1114_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1115_3_lut_3_lut (.I0(n1667), .I1(n6744), .I2(n1644), 
            .I3(GND_net), .O(n1755));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1115_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1123_3_lut_3_lut (.I0(n1667), .I1(n6752), .I2(n1652), 
            .I3(GND_net), .O(n1763));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1123_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i719_3_lut_3_lut (.I0(n1067), .I1(n6218), .I2(n1043), 
            .I3(GND_net), .O(n1169));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1198_3_lut_3_lut (.I0(n1778), .I1(n6795), .I2(n1765), 
            .I3(GND_net), .O(n1873));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1198_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10454_4_lut (.I0(n23785), .I1(r_Bit_Index_adj_4404[2]), .I2(n4038), 
            .I3(n23655), .O(n23872));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10454_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_12_i1189_3_lut_3_lut (.I0(n1778), .I1(n6786), .I2(n1756), 
            .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1189_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1187_3_lut_3_lut (.I0(n1778), .I1(n6784), .I2(n1754), 
            .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1187_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1197_3_lut_3_lut (.I0(n1778), .I1(n6794), .I2(n1764), 
            .I3(GND_net), .O(n1872));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1197_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1196_3_lut_3_lut (.I0(n1778), .I1(n6793), .I2(n1763), 
            .I3(GND_net), .O(n1871));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1196_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10450_2_lut (.I0(n23914), .I1(n23866), .I2(GND_net), .I3(GND_net), 
            .O(n23868));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10450_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1195_3_lut_3_lut (.I0(n1778), .I1(n6792), .I2(n1762), 
            .I3(GND_net), .O(n1870));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1195_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1193_3_lut_3_lut (.I0(n1778), .I1(n6790), .I2(n1760), 
            .I3(GND_net), .O(n1868));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1193_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1194_3_lut_3_lut (.I0(n1778), .I1(n6791), .I2(n1761), 
            .I3(GND_net), .O(n1869));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1194_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1192_3_lut_3_lut (.I0(n1778), .I1(n6789), .I2(n1759), 
            .I3(GND_net), .O(n1867));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1192_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i723_3_lut_3_lut (.I0(n1067), .I1(n6222), .I2(n1047), 
            .I3(GND_net), .O(n1173));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i723_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10447_2_lut (.I0(n23914), .I1(n23863), .I2(GND_net), .I3(GND_net), 
            .O(n23865));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10444_2_lut (.I0(n23914), .I1(n23860), .I2(GND_net), .I3(GND_net), 
            .O(n23862));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10444_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1199_3_lut_3_lut (.I0(n1778), .I1(n6796), .I2(n380), 
            .I3(GND_net), .O(n1874));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1199_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10441_2_lut (.I0(n23914), .I1(n23857), .I2(GND_net), .I3(GND_net), 
            .O(n23859));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10441_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1191_3_lut_3_lut (.I0(n1778), .I1(n6788), .I2(n1758), 
            .I3(GND_net), .O(n1866));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1191_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1190_3_lut_3_lut (.I0(n1778), .I1(n6787), .I2(n1757), 
            .I3(GND_net), .O(n1865));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1190_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10438_2_lut (.I0(n23914), .I1(n23854), .I2(GND_net), .I3(GND_net), 
            .O(n23856));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1188_3_lut_3_lut (.I0(n1778), .I1(n6785), .I2(n1755), 
            .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1188_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1270_3_lut_3_lut (.I0(n1886), .I1(n6837), .I2(n1874), 
            .I3(GND_net), .O(n1979));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1270_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10435_2_lut (.I0(n23914), .I1(n23851), .I2(GND_net), .I3(GND_net), 
            .O(n23853));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10435_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1260_3_lut_3_lut (.I0(n1886), .I1(n6827), .I2(n1864), 
            .I3(GND_net), .O(n1969));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1260_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10432_2_lut (.I0(n23914), .I1(n23848), .I2(GND_net), .I3(GND_net), 
            .O(n23850));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1258_3_lut_3_lut (.I0(n1886), .I1(n6825), .I2(n1862), 
            .I3(GND_net), .O(n1967));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1258_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1259_3_lut_3_lut (.I0(n1886), .I1(n6826), .I2(n1863), 
            .I3(GND_net), .O(n1968));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1259_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1269_3_lut_3_lut (.I0(n1886), .I1(n6836), .I2(n1873), 
            .I3(GND_net), .O(n1978));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1269_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1267_3_lut_3_lut (.I0(n1886), .I1(n6834), .I2(n1871), 
            .I3(GND_net), .O(n1976));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1267_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i1268_3_lut_3_lut (.I0(n1886), .I1(n6835), .I2(n1872), 
            .I3(GND_net), .O(n1977));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1268_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1265_3_lut_3_lut (.I0(n1886), .I1(n6832), .I2(n1869), 
            .I3(GND_net), .O(n1974));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1265_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10429_2_lut (.I0(n23914), .I1(n23845), .I2(GND_net), .I3(GND_net), 
            .O(n23847));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10429_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1266_3_lut_3_lut (.I0(n1886), .I1(n6833), .I2(n1870), 
            .I3(GND_net), .O(n1975));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1266_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1264_3_lut_3_lut (.I0(n1886), .I1(n6831), .I2(n1868), 
            .I3(GND_net), .O(n1973));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1264_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1271_3_lut_3_lut (.I0(n1886), .I1(n6838), .I2(n381), 
            .I3(GND_net), .O(n1980));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1271_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10479_2_lut (.I0(n28694), .I1(n23895), .I2(GND_net), .I3(GND_net), 
            .O(n23897));   // verilog/coms.v(125[12] 284[6])
    defparam i10479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10470_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_3980), 
            .I3(n22539), .O(n23888));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10470_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_12_i1263_3_lut_3_lut (.I0(n1886), .I1(n6830), .I2(n1867), 
            .I3(GND_net), .O(n1972));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1263_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1262_3_lut_3_lut (.I0(n1886), .I1(n6829), .I2(n1866), 
            .I3(GND_net), .O(n1971));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1262_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10889_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24307));   // verilog/coms.v(125[12] 284[6])
    defparam i10889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10890_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24308));   // verilog/coms.v(125[12] 284[6])
    defparam i10890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1261_3_lut_3_lut (.I0(n1886), .I1(n6828), .I2(n1865), 
            .I3(GND_net), .O(n1970));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1261_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10891_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24309));   // verilog/coms.v(125[12] 284[6])
    defparam i10891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10892_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24310));   // verilog/coms.v(125[12] 284[6])
    defparam i10892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1340_3_lut_3_lut (.I0(n1991), .I1(n6854), .I2(n1980), 
            .I3(GND_net), .O(n2082));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1340_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1712_3_lut_3_lut (.I0(n2558), .I1(n6971), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1331_3_lut_3_lut (.I0(n1991), .I1(n6845), .I2(n1971), 
            .I3(GND_net), .O(n2073));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1331_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1328_3_lut_3_lut (.I0(n1991), .I1(n6842), .I2(n1968), 
            .I3(GND_net), .O(n2070));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1328_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1330_3_lut_3_lut (.I0(n1991), .I1(n6844), .I2(n1970), 
            .I3(GND_net), .O(n2072));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1330_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1327_3_lut_3_lut (.I0(n1991), .I1(n6841), .I2(n1967), 
            .I3(GND_net), .O(n2069));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1327_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1329_3_lut_3_lut (.I0(n1991), .I1(n6843), .I2(n1969), 
            .I3(GND_net), .O(n2071));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1329_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_23_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[18]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_12_i1699_3_lut_3_lut (.I0(n2558), .I1(n6958), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_22_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_25[18]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1700_3_lut_3_lut (.I0(n2558), .I1(n6959), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1336_3_lut_3_lut (.I0(n1991), .I1(n6850), .I2(n1976), 
            .I3(GND_net), .O(n2078));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1336_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1334_3_lut_3_lut (.I0(n1991), .I1(n6848), .I2(n1974), 
            .I3(GND_net), .O(n2076));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1334_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1335_3_lut_3_lut (.I0(n1991), .I1(n6849), .I2(n1975), 
            .I3(GND_net), .O(n2077));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1335_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1339_3_lut_3_lut (.I0(n1991), .I1(n6853), .I2(n1979), 
            .I3(GND_net), .O(n2081));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1339_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1338_3_lut_3_lut (.I0(n1991), .I1(n6852), .I2(n1978), 
            .I3(GND_net), .O(n2080));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1338_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1337_3_lut_3_lut (.I0(n1991), .I1(n6851), .I2(n1977), 
            .I3(GND_net), .O(n2079));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1337_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1341_3_lut_3_lut (.I0(n1991), .I1(n6855), .I2(n382), 
            .I3(GND_net), .O(n2083));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1341_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1333_3_lut_3_lut (.I0(n1991), .I1(n6847), .I2(n1973), 
            .I3(GND_net), .O(n2075));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1333_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1702_3_lut_3_lut (.I0(n2558), .I1(n6961), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_23_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[19]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_12_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_22_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_25[19]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1332_3_lut_3_lut (.I0(n1991), .I1(n6846), .I2(n1972), 
            .I3(GND_net), .O(n2074));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1332_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1408_3_lut_3_lut (.I0(n2093), .I1(n6872), .I2(n2083), 
            .I3(GND_net), .O(n2182));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1408_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1399_3_lut_3_lut (.I0(n2093), .I1(n6863), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1409_3_lut_3_lut (.I0(n2093), .I1(n6873), .I2(n383), 
            .I3(GND_net), .O(n2183));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1409_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1397_3_lut_3_lut (.I0(n2093), .I1(n6861), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_adj_1464 (.I0(n93), .I1(n22591), .I2(GND_net), .I3(GND_net), 
            .O(n22588));
    defparam i1_2_lut_adj_1464.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_23_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[20]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14_4_lut (.I0(n21_adj_4357), .I1(n23_adj_4355), .I2(n22_adj_4356), 
            .I3(n24_adj_4354), .O(n30_adj_4352));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_22_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_25[20]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1396_3_lut_3_lut (.I0(n2093), .I1(n6860), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13_4_lut (.I0(n17_adj_4361), .I1(n19_adj_4359), .I2(n18_adj_4360), 
            .I3(n20_adj_4358), .O(n29_adj_4353));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_12_i1395_3_lut_3_lut (.I0(n2093), .I1(n6859), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1398_3_lut_3_lut (.I0(n2093), .I1(n6862), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 LessThan_556_i15_2_lut (.I0(pwm_count[7]), .I1(pwm[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4017));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_556_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_556_i9_2_lut (.I0(pwm_count[4]), .I1(pwm[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4014));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_556_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_556_i13_2_lut (.I0(pwm_count[6]), .I1(pwm[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4016));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_556_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_556_i11_2_lut (.I0(pwm_count[5]), .I1(pwm[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4015));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_556_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i1394_3_lut_3_lut (.I0(n2093), .I1(n6858), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1407_3_lut_3_lut (.I0(n2093), .I1(n6871), .I2(n2082), 
            .I3(GND_net), .O(n2181));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1407_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1405_3_lut_3_lut (.I0(n2093), .I1(n6869), .I2(n2080), 
            .I3(GND_net), .O(n2179));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1405_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32641_3_lut (.I0(n4_adj_4011), .I1(pwm[5]), .I2(n11_adj_4015), 
            .I3(GND_net), .O(n48155));   // verilog/motorControl.v(58[19:32])
    defparam i32641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32642_3_lut (.I0(n48155), .I1(pwm[6]), .I2(n13_adj_4016), 
            .I3(GND_net), .O(n48156));   // verilog/motorControl.v(58[19:32])
    defparam i32642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1406_3_lut_3_lut (.I0(n2093), .I1(n6870), .I2(n2081), 
            .I3(GND_net), .O(n2180));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1406_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32081_4_lut (.I0(n13_adj_4016), .I1(n11_adj_4015), .I2(n9_adj_4014), 
            .I3(n46943), .O(n47595));
    defparam i32081_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_556_i8_3_lut (.I0(n6_adj_4012), .I1(pwm[4]), .I2(n9_adj_4014), 
            .I3(GND_net), .O(n8_adj_4013));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_556_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31978_3_lut (.I0(n48156), .I1(pwm[7]), .I2(n15_adj_4017), 
            .I3(GND_net), .O(n47492));   // verilog/motorControl.v(58[19:32])
    defparam i31978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32679_4_lut (.I0(n47492), .I1(n8_adj_4013), .I2(n15_adj_4017), 
            .I3(n47595), .O(n48193));   // verilog/motorControl.v(58[19:32])
    defparam i32679_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_12_i1404_3_lut_3_lut (.I0(n2093), .I1(n6868), .I2(n2079), 
            .I3(GND_net), .O(n2178));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1404_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1701_3_lut_3_lut (.I0(n2558), .I1(n6960), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1403_3_lut_3_lut (.I0(n2093), .I1(n6867), .I2(n2078), 
            .I3(GND_net), .O(n2177));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1403_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1402_3_lut_3_lut (.I0(n2093), .I1(n6866), .I2(n2077), 
            .I3(GND_net), .O(n2176));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1402_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10501_3_lut (.I0(encoder0_position[23]), .I1(n2293), .I2(count_enable), 
            .I3(GND_net), .O(n23919));   // quad.v(35[10] 41[6])
    defparam i10501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1400_3_lut_3_lut (.I0(n2093), .I1(n6864), .I2(n2075), 
            .I3(GND_net), .O(n2174));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1400_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10502_3_lut (.I0(encoder0_position[22]), .I1(n2294), .I2(count_enable), 
            .I3(GND_net), .O(n23920));   // quad.v(35[10] 41[6])
    defparam i10502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1401_3_lut_3_lut (.I0(n2093), .I1(n6865), .I2(n2076), 
            .I3(GND_net), .O(n2175));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1401_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10503_3_lut (.I0(encoder0_position[21]), .I1(n2295), .I2(count_enable), 
            .I3(GND_net), .O(n23921));   // quad.v(35[10] 41[6])
    defparam i10503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10504_3_lut (.I0(encoder0_position[20]), .I1(n2296), .I2(count_enable), 
            .I3(GND_net), .O(n23922));   // quad.v(35[10] 41[6])
    defparam i10504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10505_3_lut (.I0(encoder0_position[19]), .I1(n2297), .I2(count_enable), 
            .I3(GND_net), .O(n23923));   // quad.v(35[10] 41[6])
    defparam i10505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10506_3_lut (.I0(encoder0_position[18]), .I1(n2298), .I2(count_enable), 
            .I3(GND_net), .O(n23924));   // quad.v(35[10] 41[6])
    defparam i10506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10507_3_lut (.I0(encoder0_position[17]), .I1(n2299), .I2(count_enable), 
            .I3(GND_net), .O(n23925));   // quad.v(35[10] 41[6])
    defparam i10507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10508_3_lut (.I0(encoder0_position[16]), .I1(n2300), .I2(count_enable), 
            .I3(GND_net), .O(n23926));   // quad.v(35[10] 41[6])
    defparam i10508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10509_3_lut (.I0(encoder0_position[15]), .I1(n2301), .I2(count_enable), 
            .I3(GND_net), .O(n23927));   // quad.v(35[10] 41[6])
    defparam i10509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10510_3_lut (.I0(encoder0_position[14]), .I1(n2302), .I2(count_enable), 
            .I3(GND_net), .O(n23928));   // quad.v(35[10] 41[6])
    defparam i10510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10511_3_lut (.I0(encoder0_position[13]), .I1(n2303), .I2(count_enable), 
            .I3(GND_net), .O(n23929));   // quad.v(35[10] 41[6])
    defparam i10511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[21]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10512_3_lut (.I0(encoder0_position[12]), .I1(n2304), .I2(count_enable), 
            .I3(GND_net), .O(n23930));   // quad.v(35[10] 41[6])
    defparam i10512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_25[21]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10513_3_lut (.I0(encoder0_position[11]), .I1(n2305), .I2(count_enable), 
            .I3(GND_net), .O(n23931));   // quad.v(35[10] 41[6])
    defparam i10513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10514_3_lut (.I0(encoder0_position[10]), .I1(n2306), .I2(count_enable), 
            .I3(GND_net), .O(n23932));   // quad.v(35[10] 41[6])
    defparam i10514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10515_3_lut (.I0(encoder0_position[9]), .I1(n2307), .I2(count_enable), 
            .I3(GND_net), .O(n23933));   // quad.v(35[10] 41[6])
    defparam i10515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10516_3_lut (.I0(encoder0_position[8]), .I1(n2308), .I2(count_enable), 
            .I3(GND_net), .O(n23934));   // quad.v(35[10] 41[6])
    defparam i10516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10517_3_lut (.I0(encoder0_position[7]), .I1(n2309), .I2(count_enable), 
            .I3(GND_net), .O(n23935));   // quad.v(35[10] 41[6])
    defparam i10517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10518_3_lut (.I0(encoder0_position[6]), .I1(n2310), .I2(count_enable), 
            .I3(GND_net), .O(n23936));   // quad.v(35[10] 41[6])
    defparam i10518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10519_3_lut (.I0(encoder0_position[5]), .I1(n2311), .I2(count_enable), 
            .I3(GND_net), .O(n23937));   // quad.v(35[10] 41[6])
    defparam i10519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10520_3_lut (.I0(encoder0_position[4]), .I1(n2312), .I2(count_enable), 
            .I3(GND_net), .O(n23938));   // quad.v(35[10] 41[6])
    defparam i10520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10900_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24318));   // verilog/coms.v(125[12] 284[6])
    defparam i10900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10521_3_lut (.I0(encoder0_position[3]), .I1(n2313), .I2(count_enable), 
            .I3(GND_net), .O(n23939));   // quad.v(35[10] 41[6])
    defparam i10521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10522_3_lut (.I0(encoder0_position[2]), .I1(n2314), .I2(count_enable), 
            .I3(GND_net), .O(n23940));   // quad.v(35[10] 41[6])
    defparam i10522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10523_3_lut (.I0(encoder0_position[1]), .I1(n2315), .I2(count_enable), 
            .I3(GND_net), .O(n23941));   // quad.v(35[10] 41[6])
    defparam i10523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1465 (.I0(n5_adj_3999), .I1(n122), .I2(n2119), 
            .I3(n63_adj_3998), .O(n6_adj_4366));   // verilog/coms.v(125[12] 284[6])
    defparam i1_4_lut_adj_1465.LUT_INIT = 16'heaaa;
    SB_LUT4 i3_4_lut (.I0(n50013), .I1(n6_adj_4366), .I2(n22511), .I3(n3758), 
            .O(n8_adj_3997));   // verilog/coms.v(125[12] 284[6])
    defparam i3_4_lut.LUT_INIT = 16'hcfce;
    SB_LUT4 mux_23_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[22]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i4_4_lut (.I0(n122), .I1(n8_adj_3997), .I2(n43773), .I3(n5_adj_4365), 
            .O(n49493));   // verilog/coms.v(125[12] 284[6])
    defparam i4_4_lut.LUT_INIT = 16'hefcf;
    SB_LUT4 mux_22_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_25[22]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1471_3_lut_3_lut (.I0(n2192), .I1(n6888), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10525_3_lut (.I0(\PID_CONTROLLER.err_prev [31]), .I1(\PID_CONTROLLER.err [31]), 
            .I2(n44066), .I3(GND_net), .O(n23943));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1705_3_lut_3_lut (.I0(n2558), .I1(n6964), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10526_3_lut (.I0(\PID_CONTROLLER.err_prev [23]), .I1(\PID_CONTROLLER.err [23]), 
            .I2(n44066), .I3(GND_net), .O(n23944));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10526_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10527_3_lut (.I0(\PID_CONTROLLER.err_prev [22]), .I1(\PID_CONTROLLER.err [22]), 
            .I2(n44066), .I3(GND_net), .O(n23945));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10527_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10528_3_lut (.I0(\PID_CONTROLLER.err_prev [21]), .I1(\PID_CONTROLLER.err [21]), 
            .I2(n44066), .I3(GND_net), .O(n23946));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10528_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10529_3_lut (.I0(\PID_CONTROLLER.err_prev [20]), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n44066), .I3(GND_net), .O(n23947));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10529_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10530_3_lut (.I0(\PID_CONTROLLER.err_prev [19]), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n44066), .I3(GND_net), .O(n23948));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10530_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10531_3_lut (.I0(\PID_CONTROLLER.err_prev [18]), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n44066), .I3(GND_net), .O(n23949));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10531_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10901_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24319));   // verilog/coms.v(125[12] 284[6])
    defparam i10901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10532_3_lut (.I0(\PID_CONTROLLER.err_prev [17]), .I1(\PID_CONTROLLER.err [17]), 
            .I2(n44066), .I3(GND_net), .O(n23950));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10532_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10533_3_lut (.I0(\PID_CONTROLLER.err_prev [16]), .I1(\PID_CONTROLLER.err [16]), 
            .I2(n44066), .I3(GND_net), .O(n23951));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10533_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10902_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24320));   // verilog/coms.v(125[12] 284[6])
    defparam i10902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10534_3_lut (.I0(\PID_CONTROLLER.err_prev [15]), .I1(\PID_CONTROLLER.err [15]), 
            .I2(n44066), .I3(GND_net), .O(n23952));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10534_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10535_3_lut (.I0(\PID_CONTROLLER.err_prev [14]), .I1(\PID_CONTROLLER.err [14]), 
            .I2(n44066), .I3(GND_net), .O(n23953));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10535_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10536_3_lut (.I0(\PID_CONTROLLER.err_prev [13]), .I1(\PID_CONTROLLER.err [13]), 
            .I2(n44066), .I3(GND_net), .O(n23954));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10536_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1459_3_lut_3_lut (.I0(n2192), .I1(n6876), .I2(n2168), 
            .I3(GND_net), .O(n2264_adj_3994));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10537_3_lut (.I0(\PID_CONTROLLER.err_prev [12]), .I1(\PID_CONTROLLER.err [12]), 
            .I2(n44066), .I3(GND_net), .O(n23955));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10537_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10538_3_lut (.I0(\PID_CONTROLLER.err_prev [11]), .I1(\PID_CONTROLLER.err [11]), 
            .I2(n44066), .I3(GND_net), .O(n23956));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10538_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10539_3_lut (.I0(\PID_CONTROLLER.err_prev [10]), .I1(\PID_CONTROLLER.err [10]), 
            .I2(n44066), .I3(GND_net), .O(n23957));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10539_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10540_3_lut (.I0(\PID_CONTROLLER.err_prev [9]), .I1(\PID_CONTROLLER.err [9]), 
            .I2(n44066), .I3(GND_net), .O(n23958));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10540_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10541_3_lut (.I0(\PID_CONTROLLER.err_prev [8]), .I1(\PID_CONTROLLER.err [8]), 
            .I2(n44066), .I3(GND_net), .O(n23959));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10541_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10542_3_lut (.I0(\PID_CONTROLLER.err_prev [7]), .I1(\PID_CONTROLLER.err [7]), 
            .I2(n44066), .I3(GND_net), .O(n23960));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10542_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10543_3_lut (.I0(\PID_CONTROLLER.err_prev [6]), .I1(\PID_CONTROLLER.err [6]), 
            .I2(n44066), .I3(GND_net), .O(n23961));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10543_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10544_3_lut (.I0(\PID_CONTROLLER.err_prev [5]), .I1(\PID_CONTROLLER.err [5]), 
            .I2(n44066), .I3(GND_net), .O(n23962));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10544_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1470_3_lut_3_lut (.I0(n2192), .I1(n6887), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1467_3_lut_3_lut (.I0(n2192), .I1(n6884), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10545_3_lut (.I0(\PID_CONTROLLER.err_prev [4]), .I1(\PID_CONTROLLER.err [4]), 
            .I2(n44066), .I3(GND_net), .O(n23963));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10545_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10546_3_lut (.I0(\PID_CONTROLLER.err_prev [3]), .I1(\PID_CONTROLLER.err [3]), 
            .I2(n44066), .I3(GND_net), .O(n23964));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10546_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1465_3_lut_3_lut (.I0(n2192), .I1(n6882), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1475_3_lut_3_lut (.I0(n2192), .I1(n6892), .I2(n384), 
            .I3(GND_net), .O(n2280));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10547_3_lut (.I0(\PID_CONTROLLER.err_prev [2]), .I1(\PID_CONTROLLER.err [2]), 
            .I2(n44066), .I3(GND_net), .O(n23965));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10547_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10548_3_lut (.I0(\PID_CONTROLLER.err_prev [1]), .I1(\PID_CONTROLLER.err [1]), 
            .I2(n44066), .I3(GND_net), .O(n23966));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10548_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1466 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_4362));   // verilog/TinyFPGA_B.v(147[5:22])
    defparam i4_4_lut_adj_1466.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1467 (.I0(control_mode[6]), .I1(n10_adj_4362), 
            .I2(control_mode[2]), .I3(GND_net), .O(n22531));   // verilog/TinyFPGA_B.v(147[5:22])
    defparam i5_3_lut_adj_1467.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n22531), 
            .I3(GND_net), .O(n15_adj_3958));   // verilog/TinyFPGA_B.v(147[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_23_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_3958), .I3(n15_adj_3959), .O(motor_state_23__N_25[23]));   // verilog/TinyFPGA_B.v(147[5] 150[10])
    defparam mux_23_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_25[23]), 
            .I2(n15_adj_3985), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(146[5] 150[10])
    defparam mux_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1463_3_lut_3_lut (.I0(n2192), .I1(n6880), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1462_3_lut_3_lut (.I0(n2192), .I1(n6879), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1703_3_lut_3_lut (.I0(n2558), .I1(n6962), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1461_3_lut_3_lut (.I0(n2192), .I1(n6878), .I2(n2170), 
            .I3(GND_net), .O(n2266_adj_3996));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1706_3_lut_3_lut (.I0(n2558), .I1(n6965), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_3960));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1464_3_lut_3_lut (.I0(n2192), .I1(n6881), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_3961));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1460_3_lut_3_lut (.I0(n2192), .I1(n6877), .I2(n2169), 
            .I3(GND_net), .O(n2265_adj_3995));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1474_3_lut_3_lut (.I0(n2192), .I1(n6891), .I2(n2183), 
            .I3(GND_net), .O(n2279));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1472_3_lut_3_lut (.I0(n2192), .I1(n6889), .I2(n2181), 
            .I3(GND_net), .O(n2277));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1473_3_lut_3_lut (.I0(n2192), .I1(n6890), .I2(n2182), 
            .I3(GND_net), .O(n2278));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_3962));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1719_3_lut_3_lut (.I0(n2558), .I1(n6978), .I2(n388), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1469_3_lut_3_lut (.I0(n2192), .I1(n6886), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1468_3_lut_3_lut (.I0(n2192), .I1(n6885), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1466_3_lut_3_lut (.I0(n2192), .I1(n6883), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_3963));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1704_3_lut_3_lut (.I0(n2558), .I1(n6963), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4048));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_3964));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1533_3_lut_3_lut (.I0(n2288), .I1(n6906), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_3965));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4047));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4046));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4045));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_3966));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4044));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4043));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1522_3_lut_3_lut (.I0(n2288), .I1(n6895), .I2(n2264_adj_3994), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_3967));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1525_3_lut_3_lut (.I0(n2288), .I1(n6898), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_3968));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4042));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1523_3_lut_3_lut (.I0(n2288), .I1(n6896), .I2(n2265_adj_3995), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4041));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4040));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4039));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_3969));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4038));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_3970));   // verilog/TinyFPGA_B.v(171[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1526_3_lut_3_lut (.I0(n2288), .I1(n6899), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4037));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n7009), 
            .I3(n2724), .O(n39_adj_4346));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n7008), 
            .I3(n2724), .O(n41_adj_4348));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4036));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n391));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n7006), 
            .I3(n2724), .O(n45_adj_4350));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n7007), 
            .I3(n2724), .O(n43_adj_4349));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4035));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n7010), 
            .I3(n2724), .O(n37_adj_4345));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4034));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n7014), 
            .I3(n2724), .O(n29_adj_4340));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n7013), 
            .I3(n2724), .O(n31_adj_4342));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n7018), 
            .I3(n2724), .O(n21_adj_4335));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n7017), 
            .I3(n2724), .O(n23_adj_4336));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4033));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1770_3_lut_3_lut (.I0(n2642), .I1(n6997), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n7016), 
            .I3(n2724), .O(n25_adj_4338));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n7020), 
            .I3(n2724), .O(n17_adj_4333));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n7019), 
            .I3(n2724), .O(n19_adj_4334));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4032));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n7025), 
            .I3(n2724), .O(n7_adj_4324));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n7011), 
            .I3(n2724), .O(n35_adj_4344));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n7012), 
            .I3(n2724), .O(n33_adj_4343));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_i1534_3_lut_3_lut (.I0(n2288), .I1(n6907), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n7024), 
            .I3(n2724), .O(n9_adj_4326));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n7023), 
            .I3(n2724), .O(n11_adj_4328));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n7022), 
            .I3(n2724), .O(n13_adj_4330));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4031));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4030));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n7021), 
            .I3(n2724), .O(n15_adj_4331));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n7015), 
            .I3(n2724), .O(n27_adj_4339));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31324_4_lut (.I0(n27_adj_4339), .I1(n15_adj_4331), .I2(n13_adj_4330), 
            .I3(n11_adj_4328), .O(n46836));
    defparam i31324_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4343), 
            .I3(GND_net), .O(n12_adj_4329));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i31284_2_lut (.I0(n33_adj_4343), .I1(n15_adj_4331), .I2(GND_net), 
            .I3(GND_net), .O(n46796));
    defparam i31284_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_12_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_4330), 
            .I3(GND_net), .O(n10_adj_4327));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_1830_i30_3_lut (.I0(n12_adj_4329), .I1(n83), 
            .I2(n35_adj_4344), .I3(GND_net), .O(n30_adj_4341));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1709_3_lut_3_lut (.I0(n2558), .I1(n6968), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1828_3_lut (.I0(n2720), .I1(n7026), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31424_3_lut (.I0(n7_adj_4324), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n46937));
    defparam i31424_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 i32073_4_lut (.I0(n13_adj_4330), .I1(n11_adj_4328), .I2(n9_adj_4326), 
            .I3(n46937), .O(n47587));
    defparam i32073_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32011_4_lut (.I0(n19_adj_4334), .I1(n17_adj_4333), .I2(n15_adj_4331), 
            .I3(n47587), .O(n47525));
    defparam i32011_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32875_4_lut (.I0(n25_adj_4338), .I1(n23_adj_4336), .I2(n21_adj_4335), 
            .I3(n47525), .O(n48389));
    defparam i32875_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32419_4_lut (.I0(n31_adj_4342), .I1(n29_adj_4340), .I2(n27_adj_4339), 
            .I3(n48389), .O(n47933));
    defparam i32419_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32991_4_lut (.I0(n37_adj_4345), .I1(n35_adj_4344), .I2(n33_adj_4343), 
            .I3(n47933), .O(n48505));
    defparam i32991_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_12_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4349), 
            .I3(GND_net), .O(n16_adj_4332));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4324), 
            .I3(GND_net), .O(n6_adj_4323));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i32797_3_lut (.I0(n6_adj_4323), .I1(n90), .I2(n21_adj_4335), 
            .I3(GND_net), .O(n48311));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32797_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32798_3_lut (.I0(n48311), .I1(n89), .I2(n23_adj_4336), .I3(GND_net), 
            .O(n48312));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32798_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31378_4_lut (.I0(n21_adj_4335), .I1(n19_adj_4334), .I2(n17_adj_4333), 
            .I3(n9_adj_4326), .O(n46891));
    defparam i31378_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31257_2_lut (.I0(n43_adj_4349), .I1(n19_adj_4334), .I2(GND_net), 
            .I3(GND_net), .O(n46769));
    defparam i31257_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_12_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4029));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4028));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4027));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4026));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1708_3_lut_3_lut (.I0(n2558), .I1(n6967), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1717_3_lut_3_lut (.I0(n2558), .I1(n6976), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4333), 
            .I3(GND_net), .O(n8_adj_4325));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4025));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1830_i24_3_lut (.I0(n16_adj_4332), .I1(n78), 
            .I2(n45_adj_4350), .I3(GND_net), .O(n24_adj_4337));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31261_4_lut (.I0(n43_adj_4349), .I1(n25_adj_4338), .I2(n23_adj_4336), 
            .I3(n46891), .O(n46773));
    defparam i31261_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_i1532_3_lut_3_lut (.I0(n2288), .I1(n6905), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1531_3_lut_3_lut (.I0(n2288), .I1(n6904), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32455_4_lut (.I0(n24_adj_4337), .I1(n8_adj_4325), .I2(n45_adj_4350), 
            .I3(n46769), .O(n47969));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32455_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32734_3_lut (.I0(n48312), .I1(n88), .I2(n25_adj_4338), .I3(GND_net), 
            .O(n48248));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32734_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4072));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1829_3_lut (.I0(n390), .I1(n7027), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4071));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4070));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4069));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1830_i4_4_lut (.I0(n391), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4322));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4068));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32795_3_lut (.I0(n4_adj_4322), .I1(n87), .I2(n27_adj_4339), 
            .I3(GND_net), .O(n48309));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32795_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4067));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1530_3_lut_3_lut (.I0(n2288), .I1(n6903), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32796_3_lut (.I0(n48309), .I1(n86), .I2(n29_adj_4340), .I3(GND_net), 
            .O(n48310));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32796_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4066));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31296_4_lut (.I0(n33_adj_4343), .I1(n31_adj_4342), .I2(n29_adj_4340), 
            .I3(n46836), .O(n46808));
    defparam i31296_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4065));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33037_4_lut (.I0(n30_adj_4341), .I1(n10_adj_4327), .I2(n35_adj_4344), 
            .I3(n46796), .O(n48551));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33037_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32736_3_lut (.I0(n48310), .I1(n85), .I2(n31_adj_4342), .I3(GND_net), 
            .O(n48250));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32736_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1524_3_lut_3_lut (.I0(n2288), .I1(n6897), .I2(n2266_adj_3996), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33112_4_lut (.I0(n48250), .I1(n48551), .I2(n35_adj_4344), 
            .I3(n46808), .O(n48626));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33112_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33113_3_lut (.I0(n48626), .I1(n82), .I2(n37_adj_4345), .I3(GND_net), 
            .O(n48627));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33113_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1539_3_lut_3_lut (.I0(n2288), .I1(n6912), .I2(n385), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33079_3_lut (.I0(n48627), .I1(n81), .I2(n39_adj_4346), .I3(GND_net), 
            .O(n48593));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33079_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31265_4_lut (.I0(n43_adj_4349), .I1(n41_adj_4348), .I2(n39_adj_4346), 
            .I3(n48505), .O(n46777));
    defparam i31265_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32901_4_lut (.I0(n48248), .I1(n47969), .I2(n45_adj_4350), 
            .I3(n46773), .O(n48415));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32901_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33065_3_lut (.I0(n48593), .I1(n80), .I2(n41_adj_4348), .I3(GND_net), 
            .O(n40_adj_4347));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33065_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4064));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1529_3_lut_3_lut (.I0(n2288), .I1(n6902), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1807_3_lut (.I0(n2699), .I1(n7005), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32903_4_lut (.I0(n40_adj_4347), .I1(n48415), .I2(n45_adj_4350), 
            .I3(n46777), .O(n48417));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32903_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32904_3_lut (.I0(n48417), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32904_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_12_i1528_3_lut_3_lut (.I0(n2288), .I1(n6901), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1527_3_lut_3_lut (.I0(n2288), .I1(n6900), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i1535_3_lut_3_lut (.I0(n2288), .I1(n6908), .I2(n2277), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1538_3_lut_3_lut (.I0(n2288), .I1(n6911), .I2(n2280), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_adj_1468 (.I0(n96), .I1(n22582), .I2(GND_net), .I3(GND_net), 
            .O(n22579));
    defparam i1_2_lut_adj_1468.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4319));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1537_3_lut_3_lut (.I0(n2288), .I1(n6910), .I2(n2279), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4317));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4321));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4063));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4062));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4061));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4060));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4059));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1536_3_lut_3_lut (.I0(n2288), .I1(n6909), .I2(n2278), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4320));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4058));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4057));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4312));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4056));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4313));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n390));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4055));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4314));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4315));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4303));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4305));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4054));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4311));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4053));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4052));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4307));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4309));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4310));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4316));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31482_4_lut (.I0(n29_adj_4316), .I1(n17_adj_4310), .I2(n15_adj_4309), 
            .I3(n13_adj_4307), .O(n46996));
    defparam i31482_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32143_4_lut (.I0(n11_adj_4305), .I1(n9_adj_4303), .I2(n2719), 
            .I3(n98), .O(n47657));
    defparam i32143_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i32481_4_lut (.I0(n17_adj_4310), .I1(n15_adj_4309), .I2(n13_adj_4307), 
            .I3(n47657), .O(n47995));
    defparam i32481_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32479_4_lut (.I0(n23_adj_4313), .I1(n21_adj_4312), .I2(n19_adj_4311), 
            .I3(n47995), .O(n47993));
    defparam i32479_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31499_4_lut (.I0(n29_adj_4316), .I1(n27_adj_4315), .I2(n25_adj_4314), 
            .I3(n47993), .O(n47013));
    defparam i31499_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1777_i6_4_lut (.I0(n390), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_4301));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32595_3_lut (.I0(n6_adj_4301), .I1(n87), .I2(n29_adj_4316), 
            .I3(GND_net), .O(n48109));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32595_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1777_i32_3_lut (.I0(n14_adj_4308), .I1(n83), 
            .I2(n37_adj_4321), .I3(GND_net), .O(n32_adj_4318));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32596_3_lut (.I0(n48109), .I1(n86), .I2(n31_adj_4317), .I3(GND_net), 
            .O(n48110));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32596_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31455_4_lut (.I0(n35_adj_4320), .I1(n33_adj_4319), .I2(n31_adj_4317), 
            .I3(n46996), .O(n46968));
    defparam i31455_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32987_4_lut (.I0(n32_adj_4318), .I1(n12_adj_4306), .I2(n37_adj_4321), 
            .I3(n46964), .O(n48501));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32987_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32062_3_lut (.I0(n48110), .I1(n85), .I2(n33_adj_4319), .I3(GND_net), 
            .O(n47576));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32062_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32599_3_lut (.I0(n8_adj_4302), .I1(n90), .I2(n23_adj_4313), 
            .I3(GND_net), .O(n48113));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32599_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32600_3_lut (.I0(n48113), .I1(n89), .I2(n25_adj_4314), .I3(GND_net), 
            .O(n48114));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32600_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4051));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4050));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32127_4_lut (.I0(n25_adj_4314), .I1(n23_adj_4313), .I2(n21_adj_4312), 
            .I3(n47026), .O(n47641));
    defparam i32127_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32453_3_lut (.I0(n10_adj_4304), .I1(n91), .I2(n21_adj_4312), 
            .I3(GND_net), .O(n47967));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32453_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4049));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_adj_1469 (.I0(\FRAME_MATCHER.state [2]), .I1(n22513), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n22528), .O(n43773));
    defparam i3_4_lut_adj_1469.LUT_INIT = 16'hffef;
    SB_LUT4 i32060_3_lut (.I0(n48114), .I1(n88), .I2(n27_adj_4315), .I3(GND_net), 
            .O(n47574));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32060_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32745_4_lut (.I0(n35_adj_4320), .I1(n33_adj_4319), .I2(n31_adj_4317), 
            .I3(n47013), .O(n48259));
    defparam i32745_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33092_4_lut (.I0(n47576), .I1(n48501), .I2(n37_adj_4321), 
            .I3(n46968), .O(n48606));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33092_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32799_4_lut (.I0(n47574), .I1(n47967), .I2(n27_adj_4315), 
            .I3(n47641), .O(n48313));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32799_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33126_4_lut (.I0(n48313), .I1(n48606), .I2(n37_adj_4321), 
            .I3(n48259), .O(n48640));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33126_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33127_3_lut (.I0(n48640), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n48641));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33127_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33119_3_lut (.I0(n48641), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n48633));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i33119_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i32955_3_lut (.I0(n48633), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n48469));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32955_3_lut.LUT_INIT = 16'h2b2b;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    SB_LUT4 i32956_3_lut (.I0(n48469), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n48470));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i32956_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1834_4_lut (.I0(n48470), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i1834_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 i10893_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24311));   // verilog/coms.v(125[12] 284[6])
    defparam i10893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(n98), .I1(n97), .I2(n96), .I3(n22582), 
            .O(n22573));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1470 (.I0(n97), .I1(n96), .I2(n22582), 
            .I3(GND_net), .O(n22576));
    defparam i1_2_lut_3_lut_adj_1470.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_4302));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_4306));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31451_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n46964));
    defparam i31451_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_4308));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4304));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1718_3_lut_3_lut (.I0(n2558), .I1(n6977), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31512_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n47026));
    defparam i31512_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_i1714_3_lut_3_lut (.I0(n2558), .I1(n6973), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1471 (.I0(n95), .I1(n94), .I2(n93), .I3(n22591), 
            .O(n22582));
    defparam i1_2_lut_4_lut_adj_1471.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1472 (.I0(n94), .I1(n93), .I2(n22591), 
            .I3(GND_net), .O(n22585));
    defparam i1_2_lut_3_lut_adj_1472.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1473 (.I0(n92), .I1(n91), .I2(n90), .I3(n22600), 
            .O(n22591));
    defparam i1_2_lut_4_lut_adj_1473.LUT_INIT = 16'hff7f;
    SB_LUT4 div_12_i1707_3_lut_3_lut (.I0(n2558), .I1(n6966), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1716_3_lut_3_lut (.I0(n2558), .I1(n6975), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i1711_3_lut_3_lut (.I0(n2558), .I1(n6970), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 LessThan_559_i15_2_lut (.I0(pwm_count[7]), .I1(n869), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4024));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_559_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_559_i9_2_lut (.I0(pwm_count[4]), .I1(n872), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4021));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_559_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_559_i13_2_lut (.I0(pwm_count[6]), .I1(n870), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4023));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_559_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_559_i11_2_lut (.I0(pwm_count[5]), .I1(n871), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4022));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_559_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_559_i4_3_lut (.I0(n46539), .I1(n875), .I2(pwm_count[1]), 
            .I3(GND_net), .O(n4_adj_4018));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_559_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_12_i1710_3_lut_3_lut (.I0(n2558), .I1(n6969), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32635_3_lut (.I0(n4_adj_4018), .I1(n871), .I2(n11_adj_4022), 
            .I3(GND_net), .O(n48149));   // verilog/motorControl.v(77[28:44])
    defparam i32635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32636_3_lut (.I0(n48149), .I1(n870), .I2(n13_adj_4023), .I3(GND_net), 
            .O(n48150));   // verilog/motorControl.v(77[28:44])
    defparam i32636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32007_4_lut (.I0(n13_adj_4023), .I1(n11_adj_4022), .I2(n9_adj_4021), 
            .I3(n46927), .O(n47521));
    defparam i32007_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_559_i8_3_lut (.I0(n6_adj_4019), .I1(n872), .I2(n9_adj_4021), 
            .I3(GND_net), .O(n8_adj_4020));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_559_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31998_3_lut (.I0(n48150), .I1(n869), .I2(n15_adj_4024), .I3(GND_net), 
            .O(n47512));   // verilog/motorControl.v(77[28:44])
    defparam i31998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32681_4_lut (.I0(n47512), .I1(n8_adj_4020), .I2(n15_adj_4024), 
            .I3(n47521), .O(n48195));   // verilog/motorControl.v(77[28:44])
    defparam i32681_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32682_3_lut (.I0(n48195), .I1(n868), .I2(pwm_count[8]), .I3(GND_net), 
            .O(n48196));   // verilog/motorControl.v(77[28:44])
    defparam i32682_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_1474 (.I0(n91), .I1(n90), .I2(n22600), 
            .I3(GND_net), .O(n22594));
    defparam i1_2_lut_3_lut_adj_1474.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4093));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31271_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n46783));
    defparam i31271_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4094));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1715_3_lut_3_lut (.I0(n2558), .I1(n6974), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1713_3_lut_3_lut (.I0(n2558), .I1(n6972), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1769_3_lut_3_lut (.I0(n2642), .I1(n6996), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4101));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31253_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n46765));
    defparam i31253_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4103));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1754_3_lut_3_lut (.I0(n2642), .I1(n6981), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1475 (.I0(n89), .I1(n88), .I2(n87), .I3(n22609), 
            .O(n22600));
    defparam i1_2_lut_4_lut_adj_1475.LUT_INIT = 16'hff7f;
    SB_LUT4 div_12_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4111));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31218_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n46730));
    defparam i31218_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4113));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1756_3_lut_3_lut (.I0(n2642), .I1(n6983), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10476_2_lut (.I0(n28694), .I1(n23892), .I2(GND_net), .I3(GND_net), 
            .O(n23894));   // verilog/coms.v(125[12] 284[6])
    defparam i10476_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10970_3_lut (.I0(encoder1_position[1]), .I1(n2265), .I2(count_enable_adj_3984), 
            .I3(GND_net), .O(n24388));   // quad.v(35[10] 41[6])
    defparam i10970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4123));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31188_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n46700));
    defparam i31188_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_i1757_3_lut_3_lut (.I0(n2642), .I1(n6984), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4125));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31194_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n46706));
    defparam i31194_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_4127));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4141));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31161_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n46673));
    defparam i31161_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4143));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1772_3_lut_3_lut (.I0(n2642), .I1(n6999), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31170_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n46682));
    defparam i31170_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_4145));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4159));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31143_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n46655));
    defparam i31143_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_i1758_3_lut_3_lut (.I0(n2642), .I1(n6985), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4161));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31147_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n46659));
    defparam i31147_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_4163));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4176));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31123_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n46635));
    defparam i31123_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4178));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_4180));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1755_3_lut_3_lut (.I0(n2642), .I1(n6982), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31127_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n46639));
    defparam i31127_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i1_2_lut_3_lut_adj_1476 (.I0(n88), .I1(n87), .I2(n22609), 
            .I3(GND_net), .O(n22603));
    defparam i1_2_lut_3_lut_adj_1476.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1477 (.I0(n86), .I1(n85), .I2(n84), .I3(n22618), 
            .O(n22609));
    defparam i1_2_lut_4_lut_adj_1477.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1478 (.I0(n85), .I1(n84), .I2(n22618), 
            .I3(GND_net), .O(n22612));
    defparam i1_2_lut_3_lut_adj_1478.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_4196));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31754_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n47268));
    defparam i31754_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4198));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_4200));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1761_3_lut_3_lut (.I0(n2642), .I1(n6988), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31767_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n47281));
    defparam i31767_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i10871_3_lut_4_lut (.I0(\data_out_frame[0] [2]), .I1(n3362), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n23616), .O(n24289));   // verilog/coms.v(125[12] 284[6])
    defparam i10871_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i10870_3_lut_4_lut (.I0(\data_out_frame[0] [3]), .I1(n3362), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n23616), .O(n24288));   // verilog/coms.v(125[12] 284[6])
    defparam i10870_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i1_2_lut_4_lut_adj_1479 (.I0(n83), .I1(n82), .I2(n81), .I3(n22627), 
            .O(n22618));
    defparam i1_2_lut_4_lut_adj_1479.LUT_INIT = 16'hff7f;
    SB_LUT4 i10869_3_lut_4_lut (.I0(\data_out_frame[0] [4]), .I1(n3362), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n23616), .O(n24287));   // verilog/coms.v(125[12] 284[6])
    defparam i10869_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i1_2_lut_3_lut_adj_1480 (.I0(n82), .I1(n81), .I2(n22627), 
            .I3(GND_net), .O(n22621));
    defparam i1_2_lut_3_lut_adj_1480.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_i1762_3_lut_3_lut (.I0(n2642), .I1(n6989), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1759_3_lut_3_lut (.I0(n2642), .I1(n6986), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1760_3_lut_3_lut (.I0(n2642), .I1(n6987), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_adj_1481 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n22627));
    defparam i1_2_lut_4_lut_adj_1481.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1482 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n22630));
    defparam i1_2_lut_3_lut_adj_1482.LUT_INIT = 16'hf7f7;
    SB_LUT4 i22577_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n370), .I3(n558), 
            .O(n4_adj_3953));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22577_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i22601_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n371), .I3(n558), 
            .O(n4));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22601_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i22633_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n372), .I3(n558), 
            .O(n4_adj_4075));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam i22633_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_12_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4214));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31712_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n47226));
    defparam i31712_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4216));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_4218));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1768_3_lut_3_lut (.I0(n2642), .I1(n6995), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31685_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n47199));
    defparam i31685_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4220));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4236));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31667_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n47181));
    defparam i31667_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_i1766_3_lut_3_lut (.I0(n2642), .I1(n6993), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31414_3_lut_4_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(pwm_count[2]), .O(n46927));   // verilog/motorControl.v(77[28:44])
    defparam i31414_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_559_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(GND_net), .O(n6_adj_4019));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_559_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_12_i1771_3_lut_3_lut (.I0(n2642), .I1(n6998), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4238));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_4240));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31643_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n47157));
    defparam i31643_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4242));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n22573), 
            .O(n249));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    coms c0 (.clk32MHz(clk32MHz), .n22513(n22513), .GND_net(GND_net), 
         .\Kd[7] (Kd[7]), .gearBoxRatio({gearBoxRatio}), .rx_data({rx_data}), 
         .IntegralLimit({IntegralLimit}), .n24320(n24320), .\data_in[0] ({\data_in[0] }), 
         .n24319(n24319), .n24318(n24318), .\deadband[9] (deadband[9]), 
         .\deadband[8] (deadband[8]), .\deadband[7] (deadband[7]), .\deadband[6] (deadband[6]), 
         .\deadband[5] (deadband[5]), .\deadband[4] (deadband[4]), .\deadband[3] (deadband[3]), 
         .\deadband[2] (deadband[2]), .n24482(n24482), .VCC_net(VCC_net), 
         .byte_transmit_counter({Open_0, Open_1, Open_2, Open_3, Open_4, 
         Open_5, Open_6, byte_transmit_counter[0]}), .\deadband[1] (deadband[1]), 
         .n24478(n24478), .setpoint({setpoint}), .n24477(n24477), .n24476(n24476), 
         .n24475(n24475), .n24474(n24474), .n24473(n24473), .n24472(n24472), 
         .n24471(n24471), .n24470(n24470), .n24469(n24469), .n24468(n24468), 
         .n24467(n24467), .n24466(n24466), .n24465(n24465), .n24464(n24464), 
         .n24463(n24463), .n24462(n24462), .n24461(n24461), .n24460(n24460), 
         .n24459(n24459), .n24458(n24458), .n24457(n24457), .n24456(n24456), 
         .n23891(n23891), .n24306(n24306), .\data_in[1] ({\data_in[1] }), 
         .n24305(n24305), .\data_in[2] ({\data_in[2] }), .n24304(n24304), 
         .n24303(n24303), .n24302(n24302), .n24301(n24301), .n24300(n24300), 
         .n24299(n24299), .n24298(n24298), .n24297(n24297), .\data_in[3] ({\data_in[3] }), 
         .n24296(n24296), .n24295(n24295), .n24294(n24294), .n24293(n24293), 
         .n24292(n24292), .n24291(n24291), .n24290(n24290), .n24289(n24289), 
         .\data_out_frame[0][2] (\data_out_frame[0] [2]), .n24288(n24288), 
         .\data_out_frame[0][3] (\data_out_frame[0] [3]), .n24287(n24287), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .n24284(n24284), 
         .\data_out_frame[5][2] (\data_out_frame[5] [2]), .n24317(n24317), 
         .n24316(n24316), .n24315(n24315), .n24314(n24314), .rx_data_ready(rx_data_ready), 
         .n24313(n24313), .n24312(n24312), .\Kp[1] (Kp[1]), .\Kp[2] (Kp[2]), 
         .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), .n22525(n22525), 
         .n24158(n24158), .\data_out_frame[22] ({Open_7, Open_8, Open_9, 
         Open_10, Open_11, Open_12, \data_out_frame[22] [1], Open_13}), 
         .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\FRAME_MATCHER.state[2] (\FRAME_MATCHER.state [2]), 
         .n22498(n22498), .encoder0_position({encoder0_position}), .displacement({displacement}), 
         .\Kp[5] (Kp[5]), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .n22528(n22528), .n23894(n23894), .pwm({pwm}), .encoder1_position({encoder1_position}), 
         .control_mode({control_mode}), .n23907(n23907), .n3840(n3840), 
         .n23904(n23904), .n23901(n23901), .n24311(n24311), .\Kp[6] (Kp[6]), 
         .n23898(n23898), .n41946(n41946), .n23895(n23895), .n23892(n23892), 
         .n23889(n23889), .n2241(n2241), .\PWMLimit[1] (PWMLimit[1]), 
         .\PWMLimit[2] (PWMLimit[2]), .\PWMLimit[3] (PWMLimit[3]), .\PWMLimit[4] (PWMLimit[4]), 
         .\PWMLimit[5] (PWMLimit[5]), .\PWMLimit[6] (PWMLimit[6]), .\PWMLimit[7] (PWMLimit[7]), 
         .\PWMLimit[8] (PWMLimit[8]), .\PWMLimit[9] (PWMLimit[9]), .n49493(n49493), 
         .\Kp[7] (Kp[7]), .\Ki[1] (Ki[1]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), 
         .n24310(n24310), .n24309(n24309), .\Ki[4] (Ki[4]), .n5025(n5025), 
         .n5023(n5023), .n23616(n23616), .n24308(n24308), .n3362(n3362), 
         .n24307(n24307), .\Ki[5] (Ki[5]), .n23897(n23897), .n23900(n23900), 
         .n23903(n23903), .n23906(n23906), .n23909(n23909), .\Ki[6] (Ki[6]), 
         .\Ki[7] (Ki[7]), .\Kd[1] (Kd[1]), .\Kd[2] (Kd[2]), .\Kd[3] (Kd[3]), 
         .\Kd[4] (Kd[4]), .\Kd[5] (Kd[5]), .\Kd[6] (Kd[6]), .\deadband[0] (deadband[0]), 
         .n23828(n23828), .n42006(n42006), .\PWMLimit[0] (PWMLimit[0]), 
         .n23808(n23808), .\Kd[0] (Kd[0]), .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), 
         .n3800(n3800), .n3801(n3801), .n3802(n3802), .n3803(n3803), 
         .n3804(n3804), .n3805(n3805), .n3806(n3806), .n3807(n3807), 
         .n3808(n3808), .n3809(n3809), .n3810(n3810), .n3811(n3811), 
         .n3812(n3812), .n3813(n3813), .n3814(n3814), .n3815(n3815), 
         .n3816(n3816), .n3817(n3817), .n3818(n3818), .n3819(n3819), 
         .n3820(n3820), .n3821(n3821), .n3823(n3823), .n3822(n3822), 
         .n44107(n44107), .n28694(n28694), .n122(n122), .n2854(n2854), 
         .n63(n63_adj_3998), .n5(n5_adj_3999), .n50013(n50013), .n39599(n39599), 
         .\FRAME_MATCHER.state_31__N_1860[1] (\FRAME_MATCHER.state_31__N_1860 [1]), 
         .n43447(n43447), .n22512(n22512), .n43773(n43773), .n2119(n2119), 
         .n3758(n3758), .n737(n737), .n20156(n20156), .n3(n3_adj_4364), 
         .n22511(n22511), .n5_adj_3(n5_adj_4365), .n23847(n23847), .n23850(n23850), 
         .n23853(n23853), .n23856(n23856), .n23859(n23859), .n23862(n23862), 
         .n23865(n23865), .n23868(n23868), .n23872(n23872), .r_Bit_Index({r_Bit_Index_adj_4404}), 
         .n23875(n23875), .n23845(n23845), .n23848(n23848), .n23851(n23851), 
         .n23915(n23915), .n23918(n23918), .n23854(n23854), .n23857(n23857), 
         .n23860(n23860), .n23863(n23863), .n23866(n23866), .n23913(n23913), 
         .tx_o(tx_o), .n23655(n23655), .n23785(n23785), .n4038(n4038), 
         .n23914(n23914), .tx_enable(tx_enable), .n23878(n23878), .r_Bit_Index_adj_9({r_Bit_Index}), 
         .n23881(n23881), .n24453(n24453), .n29023(n29023), .\r_SM_Main[1] (r_SM_Main[1]), 
         .r_Rx_Data(r_Rx_Data), .LED_c(LED_c), .n24391(n24391), .\r_SM_Main[2] (r_SM_Main[2]), 
         .n23888(n23888), .n23887(n23887), .n23886(n23886), .n23885(n23885), 
         .n23884(n23884), .n23883(n23883), .n23882(n23882), .n23817(n23817), 
         .n46591(n46591), .n22534(n22534), .n4(n4_adj_3980), .n28989(n28989), 
         .n28517(n28517), .n4_adj_7(n4_adj_3986), .n4_adj_8(n4_adj_3981), 
         .n23649(n23649), .n23783(n23783), .n4016(n4016), .n22539(n22539), 
         .n1(n1_adj_4351), .n46590(n46590)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(88[8] 107[4])
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n24406(n24406), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n24405(n24405), .n24404(n24404), .n24422(n24422), 
            .n24421(n24421), .n24420(n24420), .n24419(n24419), .n24418(n24418), 
            .n24417(n24417), .n24416(n24416), .n24415(n24415), .n24414(n24414), 
            .n24413(n24413), .n24412(n24412), .n24411(n24411), .n24410(n24410), 
            .n24409(n24409), .n24408(n24408), .n24407(n24407), .n24403(n24403), 
            .data_o({quadA_debounced_adj_3982, quadB_debounced_adj_3983}), 
            .n24402(n24402), .n24401(n24401), .n24388(n24388), .count_enable(count_enable_adj_3984), 
            .n2242({n2243, n2244, n2245, n2246, n2247, n2248, n2249, 
            n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, 
            n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, 
            n2266}), .GND_net(GND_net), .n23815(n23815), .n24452(n24452), 
            .PIN_23_c_0(PIN_23_c_0), .reg_B({reg_B_adj_4411}), .PIN_24_c_1(PIN_24_c_1), 
            .n23821(n23821), .n44154(n44154)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(183[15] 188[4])
    SB_LUT4 div_12_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4258));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31621_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n47135));
    defparam i31621_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4260));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1767_3_lut_3_lut (.I0(n2642), .I1(n6994), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1775_3_lut_3_lut (.I0(n2642), .I1(n7002), .I2(n389), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_4262));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31597_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n47111));
    defparam i31597_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4264));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i3_3_lut_4_lut (.I0(n2119), .I1(n3_adj_4364), .I2(n44592), 
            .I3(n43447), .O(n44557));   // verilog/coms.v(125[12] 284[6])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_1483 (.I0(n2119), .I1(n3_adj_4364), .I2(\FRAME_MATCHER.state_31__N_1860 [1]), 
            .I3(GND_net), .O(n41946));   // verilog/coms.v(125[12] 284[6])
    defparam i1_2_lut_3_lut_adj_1483.LUT_INIT = 16'he0e0;
    SB_LUT4 div_12_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_4280));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_4284));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31555_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n47069));
    defparam i31555_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_4286));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_4282));   // verilog/TinyFPGA_B.v(171[21:53])
    defparam div_12_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31575_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n47089));
    defparam i31575_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i10740_3_lut_4_lut (.I0(\data_out_frame[22] [1]), .I1(n39599), 
            .I2(n5025), .I3(n5023), .O(n24158));   // verilog/coms.v(125[12] 284[6])
    defparam i10740_3_lut_4_lut.LUT_INIT = 16'ha3aa;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n2292, encoder0_position, GND_net, 
            data_o, clk32MHz, n23941, n23940, n23939, n23938, n23937, 
            n23936, n23935, n23934, n23933, n23932, n23931, n23930, 
            n23929, n23928, n23927, n23926, n23925, n23924, n23923, 
            n23922, n23921, n23920, n23919, n23814, count_enable, 
            n24423, PIN_8_c_1, reg_B, PIN_9_c_0, n23816, n44475) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]n2292;
    output [23:0]encoder0_position;
    input GND_net;
    output [1:0]data_o;
    input clk32MHz;
    input n23941;
    input n23940;
    input n23939;
    input n23938;
    input n23937;
    input n23936;
    input n23935;
    input n23934;
    input n23933;
    input n23932;
    input n23931;
    input n23930;
    input n23929;
    input n23928;
    input n23927;
    input n23926;
    input n23925;
    input n23924;
    input n23923;
    input n23922;
    input n23921;
    input n23920;
    input n23919;
    input n23814;
    output count_enable;
    input n24423;
    input PIN_8_c_1;
    output [1:0]reg_B;
    input PIN_9_c_0;
    input n23816;
    output n44475;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n2288, n36512, n36513, n36511, n36510, n36509, count_direction, 
        n36508, B_delayed, A_delayed, n36531, n36530, n36529, n36528, 
        n36527, n36526, n36525, n36524, n36523, n36522, n36521, 
        n36520, n36519, n36518, n36517, n36516, n36514, n36515;
    
    SB_LUT4 add_550_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2288), 
            .I3(n36512), .O(n2292[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_6 (.CI(n36512), .I0(encoder0_position[4]), .I1(n2288), 
            .CO(n36513));
    SB_LUT4 add_550_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2288), 
            .I3(n36511), .O(n2292[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_5 (.CI(n36511), .I0(encoder0_position[3]), .I1(n2288), 
            .CO(n36512));
    SB_LUT4 add_550_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2288), 
            .I3(n36510), .O(n2292[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_4 (.CI(n36510), .I0(encoder0_position[2]), .I1(n2288), 
            .CO(n36511));
    SB_LUT4 add_550_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2288), 
            .I3(n36509), .O(n2292[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_3 (.CI(n36509), .I0(encoder0_position[1]), .I1(n2288), 
            .CO(n36510));
    SB_LUT4 add_550_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n36508), .O(n2292[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_2 (.CI(n36508), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n36509));
    SB_CARRY add_550_1 (.CI(GND_net), .I0(n2288), .I1(n2288), .CO(n36508));
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_550_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2288), 
            .I3(n36531), .O(n2292[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_550_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2288), 
            .I3(n36530), .O(n2292[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_24 (.CI(n36530), .I0(encoder0_position[22]), .I1(n2288), 
            .CO(n36531));
    SB_LUT4 add_550_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2288), 
            .I3(n36529), .O(n2292[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_23 (.CI(n36529), .I0(encoder0_position[21]), .I1(n2288), 
            .CO(n36530));
    SB_LUT4 add_550_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2288), 
            .I3(n36528), .O(n2292[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_22 (.CI(n36528), .I0(encoder0_position[20]), .I1(n2288), 
            .CO(n36529));
    SB_LUT4 add_550_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2288), 
            .I3(n36527), .O(n2292[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_21 (.CI(n36527), .I0(encoder0_position[19]), .I1(n2288), 
            .CO(n36528));
    SB_LUT4 add_550_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2288), 
            .I3(n36526), .O(n2292[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_20 (.CI(n36526), .I0(encoder0_position[18]), .I1(n2288), 
            .CO(n36527));
    SB_LUT4 add_550_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2288), 
            .I3(n36525), .O(n2292[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_19 (.CI(n36525), .I0(encoder0_position[17]), .I1(n2288), 
            .CO(n36526));
    SB_LUT4 add_550_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2288), 
            .I3(n36524), .O(n2292[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_18 (.CI(n36524), .I0(encoder0_position[16]), .I1(n2288), 
            .CO(n36525));
    SB_LUT4 add_550_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2288), 
            .I3(n36523), .O(n2292[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_17 (.CI(n36523), .I0(encoder0_position[15]), .I1(n2288), 
            .CO(n36524));
    SB_LUT4 add_550_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2288), 
            .I3(n36522), .O(n2292[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_16 (.CI(n36522), .I0(encoder0_position[14]), .I1(n2288), 
            .CO(n36523));
    SB_LUT4 add_550_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2288), 
            .I3(n36521), .O(n2292[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_15 (.CI(n36521), .I0(encoder0_position[13]), .I1(n2288), 
            .CO(n36522));
    SB_LUT4 add_550_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2288), 
            .I3(n36520), .O(n2292[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_14 (.CI(n36520), .I0(encoder0_position[12]), .I1(n2288), 
            .CO(n36521));
    SB_LUT4 add_550_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2288), 
            .I3(n36519), .O(n2292[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_13 (.CI(n36519), .I0(encoder0_position[11]), .I1(n2288), 
            .CO(n36520));
    SB_LUT4 add_550_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2288), 
            .I3(n36518), .O(n2292[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_12 (.CI(n36518), .I0(encoder0_position[10]), .I1(n2288), 
            .CO(n36519));
    SB_LUT4 add_550_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2288), 
            .I3(n36517), .O(n2292[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_11 (.CI(n36517), .I0(encoder0_position[9]), .I1(n2288), 
            .CO(n36518));
    SB_LUT4 add_550_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2288), 
            .I3(n36516), .O(n2292[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_10 (.CI(n36516), .I0(encoder0_position[8]), .I1(n2288), 
            .CO(n36517));
    SB_LUT4 add_550_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2288), 
            .I3(n36513), .O(n2292[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_8 (.CI(n36514), .I0(encoder0_position[6]), .I1(n2288), 
            .CO(n36515));
    SB_LUT4 add_550_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2288), 
            .I3(n36514), .O(n2292[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_9 (.CI(n36515), .I0(encoder0_position[7]), .I1(n2288), 
            .CO(n36516));
    SB_LUT4 add_550_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2288), 
            .I3(n36515), .O(n2292[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_550_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_550_7 (.CI(n36513), .I0(encoder0_position[5]), .I1(n2288), 
            .CO(n36514));
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n23941));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n23940));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n23939));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n23938));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n23937));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n23936));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n23935));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n23934));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n23933));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n23932));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n23931));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n23930));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n23929));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n23928));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n23927));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n23926));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n23925));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n23924));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n23923));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n23922));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n23921));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n23920));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n23919));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n23814));   // quad.v(35[10] 41[6])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i767_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2288));   // quad.v(37[5] 40[8])
    defparam i767_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n24423(n24423), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .PIN_8_c_1(PIN_8_c_1), .reg_B({reg_B}), 
            .PIN_9_c_0(PIN_9_c_0), .n23816(n23816), .n44475(n44475), .GND_net(GND_net)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n24423, data_o, clk32MHz, PIN_8_c_1, 
            reg_B, PIN_9_c_0, n23816, n44475, GND_net) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n24423;
    output [1:0]data_o;
    input clk32MHz;
    input PIN_8_c_1;
    output [1:0]reg_B;
    input PIN_9_c_0;
    input n23816;
    output n44475;
    input GND_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n1;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3104;
    wire [2:0]n17;
    
    wire n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n24423));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_8_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1050__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n1), .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_9_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1050__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1050__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n23816));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[2]), 
            .I3(GND_net), .O(n44475));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i22862_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22862_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22855_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22855_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n44475), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i1275_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(170[42:59])
    defparam i1275_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, VCC_net, \PID_CONTROLLER.err[31] , \Kd[1] , 
            \Kd[0] , \Kd[2] , \Kd[3] , \deadband[3] , \Kd[4] , \Kd[5] , 
            \Kd[6] , \motor_state[23] , \deadband[4] , \Kd[7] , \motor_state[22] , 
            setpoint, \motor_state[21] , \motor_state[20] , \Kp[1] , 
            \PID_CONTROLLER.err[23] , \Kp[0] , \Kp[2] , \motor_state[19] , 
            \Kp[3] , \Kp[4] , \motor_state[18] , \Kp[5] , n24454, 
            pwm, clk32MHz, n24451, n24450, n24449, n24448, n24447, 
            n41480, n24444, n24443, n24442, n24441, n24440, n24439, 
            n24438, n24437, n24436, n24434, n24431, n24430, n24426, 
            \Kp[6] , \Kp[7] , \PID_CONTROLLER.err[14] , \PID_CONTROLLER.err[15] , 
            \deadband[5] , \PID_CONTROLLER.err[21] , \PID_CONTROLLER.err[22] , 
            \motor_state[17] , \motor_state[16] , \motor_state[15] , \motor_state[14] , 
            \motor_state[13] , \Ki[1] , \PID_CONTROLLER.err[0] , \motor_state[12] , 
            \Ki[0] , \motor_state[11] , \motor_state[10] , \Ki[2] , 
            \motor_state[9] , \Ki[3] , \motor_state[8] , \Ki[4] , \motor_state[7] , 
            \PWMLimit[2] , \motor_state[6] , \motor_state[5] , \motor_state[4] , 
            \Ki[5] , \motor_state[3] , \pwm_23__N_2951[7] , \Ki[6] , 
            \motor_state[2] , \motor_state[1] , \Ki[7] , \pwm_23__N_2951[5] , 
            \motor_state[0] , \pwm_23__N_2951[4] , \deadband[6] , \PID_CONTROLLER.err_prev[31] , 
            \deadband[7] , \PID_CONTROLLER.err_prev[23] , \PID_CONTROLLER.err_prev[22] , 
            \PID_CONTROLLER.err_prev[21] , \PID_CONTROLLER.err_prev[20] , 
            \PWMLimit[3] , \deadband[8] , \PID_CONTROLLER.err_prev[19] , 
            \PID_CONTROLLER.err_prev[18] , \PID_CONTROLLER.err_prev[17] , 
            \PID_CONTROLLER.err_prev[16] , \PID_CONTROLLER.err_prev[15] , 
            \PID_CONTROLLER.err_prev[14] , \PID_CONTROLLER.err_prev[13] , 
            \PID_CONTROLLER.err_prev[12] , \PID_CONTROLLER.err_prev[11] , 
            \PID_CONTROLLER.err_prev[10] , \PID_CONTROLLER.err_prev[9] , 
            \deadband[9] , \PID_CONTROLLER.err_prev[8] , \PID_CONTROLLER.err_prev[7] , 
            \PID_CONTROLLER.err_prev[6] , \PID_CONTROLLER.err_prev[5] , 
            \PID_CONTROLLER.err_prev[4] , \PID_CONTROLLER.err_prev[3] , 
            \PID_CONTROLLER.err_prev[2] , \PID_CONTROLLER.err_prev[1] , 
            \PID_CONTROLLER.err_prev[0] , n22, n21, n24, n20, n23, 
            n19, \PID_CONTROLLER.err[10] , \PID_CONTROLLER.err[11] , IntegralLimit, 
            n17, n48196, n18, n868, n869, n870, n871, n872, 
            n873, n874, n875, n46539, \PID_CONTROLLER.err[9] , \PID_CONTROLLER.err[8] , 
            \PID_CONTROLLER.err[7] , \PID_CONTROLLER.err[6] , \PID_CONTROLLER.err[5] , 
            \PID_CONTROLLER.err[4] , \PID_CONTROLLER.err[3] , \PID_CONTROLLER.err[2] , 
            \PID_CONTROLLER.err[1] , \pwm_count[8] , \pwm_count[7] , \pwm_count[6] , 
            \pwm_count[5] , \pwm_count[4] , \pwm_count[3] , \pwm_count[2] , 
            \pwm_count[1] , n23966, n23965, n23964, n23963, n23962, 
            n23961, n23960, n23959, n23958, n23957, n23956, n23955, 
            n23954, n23953, n23952, n23951, n23950, n23949, n23948, 
            n23947, n23946, n23945, n23944, n23943, \PID_CONTROLLER.result[4] , 
            \PID_CONTROLLER.result[5] , \PID_CONTROLLER.result[7] , PIN_6_c_0, 
            PIN_5_c_1, PIN_4_c_2, PIN_3_c_3, PIN_2_c_4, \PID_CONTROLLER.err[12] , 
            \PID_CONTROLLER.err[13] , \PID_CONTROLLER.err[16] , \PID_CONTROLLER.err[17] , 
            \PID_CONTROLLER.err[18] , \PID_CONTROLLER.err[19] , \PID_CONTROLLER.err[20] , 
            hall3, PIN_1_c_5, n413, n415, n23812, n416, n421, 
            n470, n469, n468, pwm_23__N_2948, n28170, \PWMLimit[4] , 
            n387, n28227, \PWMLimit[5] , n465, n1, \PWMLimit[7] , 
            n463, n462, n461, n460, n459, n458, n457, n456, 
            n455, \PWMLimit[9] , n9, n15, \deadband[2] , \deadband[0] , 
            \deadband[1] , \PWMLimit[6] , n11, n9_adj_10, n15_adj_11, 
            \PWMLimit[8] , n11_adj_12, n9_adj_13, n15_adj_14, n11_adj_15, 
            n9_adj_16, n15_adj_17, n471, \PWMLimit[0] , \PWMLimit[1] , 
            hall2, hall1, n29, n30, n48193, n46604, n46565, n46567, 
            n46573, n46571, n46569, n44066, n4) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input VCC_net;
    output \PID_CONTROLLER.err[31] ;
    input \Kd[1] ;
    input \Kd[0] ;
    input \Kd[2] ;
    input \Kd[3] ;
    input \deadband[3] ;
    input \Kd[4] ;
    input \Kd[5] ;
    input \Kd[6] ;
    input \motor_state[23] ;
    input \deadband[4] ;
    input \Kd[7] ;
    input \motor_state[22] ;
    input [23:0]setpoint;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \Kp[1] ;
    output \PID_CONTROLLER.err[23] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \motor_state[19] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \motor_state[18] ;
    input \Kp[5] ;
    input n24454;
    output [23:0]pwm;
    input clk32MHz;
    input n24451;
    input n24450;
    input n24449;
    input n24448;
    input n24447;
    input n41480;
    input n24444;
    input n24443;
    input n24442;
    input n24441;
    input n24440;
    input n24439;
    input n24438;
    input n24437;
    input n24436;
    input n24434;
    input n24431;
    input n24430;
    input n24426;
    input \Kp[6] ;
    input \Kp[7] ;
    output \PID_CONTROLLER.err[14] ;
    output \PID_CONTROLLER.err[15] ;
    input \deadband[5] ;
    output \PID_CONTROLLER.err[21] ;
    output \PID_CONTROLLER.err[22] ;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input \Ki[1] ;
    output \PID_CONTROLLER.err[0] ;
    input \motor_state[12] ;
    input \Ki[0] ;
    input \motor_state[11] ;
    input \motor_state[10] ;
    input \Ki[2] ;
    input \motor_state[9] ;
    input \Ki[3] ;
    input \motor_state[8] ;
    input \Ki[4] ;
    input \motor_state[7] ;
    input \PWMLimit[2] ;
    input \motor_state[6] ;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input \Ki[5] ;
    input \motor_state[3] ;
    output \pwm_23__N_2951[7] ;
    input \Ki[6] ;
    input \motor_state[2] ;
    input \motor_state[1] ;
    input \Ki[7] ;
    output \pwm_23__N_2951[5] ;
    input \motor_state[0] ;
    output \pwm_23__N_2951[4] ;
    input \deadband[6] ;
    output \PID_CONTROLLER.err_prev[31] ;
    input \deadband[7] ;
    output \PID_CONTROLLER.err_prev[23] ;
    output \PID_CONTROLLER.err_prev[22] ;
    output \PID_CONTROLLER.err_prev[21] ;
    output \PID_CONTROLLER.err_prev[20] ;
    input \PWMLimit[3] ;
    input \deadband[8] ;
    output \PID_CONTROLLER.err_prev[19] ;
    output \PID_CONTROLLER.err_prev[18] ;
    output \PID_CONTROLLER.err_prev[17] ;
    output \PID_CONTROLLER.err_prev[16] ;
    output \PID_CONTROLLER.err_prev[15] ;
    output \PID_CONTROLLER.err_prev[14] ;
    output \PID_CONTROLLER.err_prev[13] ;
    output \PID_CONTROLLER.err_prev[12] ;
    output \PID_CONTROLLER.err_prev[11] ;
    output \PID_CONTROLLER.err_prev[10] ;
    output \PID_CONTROLLER.err_prev[9] ;
    input \deadband[9] ;
    output \PID_CONTROLLER.err_prev[8] ;
    output \PID_CONTROLLER.err_prev[7] ;
    output \PID_CONTROLLER.err_prev[6] ;
    output \PID_CONTROLLER.err_prev[5] ;
    output \PID_CONTROLLER.err_prev[4] ;
    output \PID_CONTROLLER.err_prev[3] ;
    output \PID_CONTROLLER.err_prev[2] ;
    output \PID_CONTROLLER.err_prev[1] ;
    output \PID_CONTROLLER.err_prev[0] ;
    output n22;
    output n21;
    output n24;
    output n20;
    output n23;
    output n19;
    output \PID_CONTROLLER.err[10] ;
    output \PID_CONTROLLER.err[11] ;
    input [23:0]IntegralLimit;
    output n17;
    input n48196;
    output n18;
    output n868;
    output n869;
    output n870;
    output n871;
    output n872;
    output n873;
    output n874;
    output n875;
    output n46539;
    output \PID_CONTROLLER.err[9] ;
    output \PID_CONTROLLER.err[8] ;
    output \PID_CONTROLLER.err[7] ;
    output \PID_CONTROLLER.err[6] ;
    output \PID_CONTROLLER.err[5] ;
    output \PID_CONTROLLER.err[4] ;
    output \PID_CONTROLLER.err[3] ;
    output \PID_CONTROLLER.err[2] ;
    output \PID_CONTROLLER.err[1] ;
    output \pwm_count[8] ;
    output \pwm_count[7] ;
    output \pwm_count[6] ;
    output \pwm_count[5] ;
    output \pwm_count[4] ;
    output \pwm_count[3] ;
    output \pwm_count[2] ;
    output \pwm_count[1] ;
    input n23966;
    input n23965;
    input n23964;
    input n23963;
    input n23962;
    input n23961;
    input n23960;
    input n23959;
    input n23958;
    input n23957;
    input n23956;
    input n23955;
    input n23954;
    input n23953;
    input n23952;
    input n23951;
    input n23950;
    input n23949;
    input n23948;
    input n23947;
    input n23946;
    input n23945;
    input n23944;
    input n23943;
    output \PID_CONTROLLER.result[4] ;
    output \PID_CONTROLLER.result[5] ;
    output \PID_CONTROLLER.result[7] ;
    output PIN_6_c_0;
    output PIN_5_c_1;
    output PIN_4_c_2;
    output PIN_3_c_3;
    output PIN_2_c_4;
    output \PID_CONTROLLER.err[12] ;
    output \PID_CONTROLLER.err[13] ;
    output \PID_CONTROLLER.err[16] ;
    output \PID_CONTROLLER.err[17] ;
    output \PID_CONTROLLER.err[18] ;
    output \PID_CONTROLLER.err[19] ;
    output \PID_CONTROLLER.err[20] ;
    input hall3;
    output PIN_1_c_5;
    output n413;
    output n415;
    input n23812;
    output n416;
    output n421;
    output n470;
    output n469;
    output n468;
    output pwm_23__N_2948;
    input n28170;
    input \PWMLimit[4] ;
    output n387;
    input n28227;
    input \PWMLimit[5] ;
    output n465;
    input n1;
    input \PWMLimit[7] ;
    output n463;
    output n462;
    output n461;
    output n460;
    output n459;
    output n458;
    output n457;
    output n456;
    output n455;
    input \PWMLimit[9] ;
    input n9;
    input n15;
    input \deadband[2] ;
    input \deadband[0] ;
    input \deadband[1] ;
    input \PWMLimit[6] ;
    input n11;
    input n9_adj_10;
    input n15_adj_11;
    input \PWMLimit[8] ;
    input n11_adj_12;
    input n9_adj_13;
    input n15_adj_14;
    input n11_adj_15;
    input n9_adj_16;
    input n15_adj_17;
    output n471;
    input \PWMLimit[0] ;
    input \PWMLimit[1] ;
    input hall2;
    input hall1;
    input n29;
    input n30;
    input n48193;
    output n46604;
    output n46565;
    output n46567;
    output n46573;
    output n46571;
    output n46569;
    output n44066;
    output n4;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [18:0]n8257;
    wire [17:0]n8278;
    
    wire n425, n37911, n37912, n37445;
    wire [6:0]Kd_delay_counter;   // verilog/motorControl.v(20[13:29])
    
    wire n37446;
    wire [6:0]n57;
    
    wire n37444;
    wire [22:0]n1800;
    wire [22:0]n1801;
    
    wire n38284, n328, n37910, n37443, n231, n37909, n37442, n38285, 
        n41, n134, n38283;
    wire [19:0]n8235;
    
    wire n37908, n37907, n37906;
    wire [31:0]n58;
    wire [31:0]n61;
    
    wire n36567, n36568, n36566, n37905, n524, n38282, n37904, 
        n451, n38281, n37903, n37902, n378, n38280, n305, n38279, 
        n37901, n37900, n36565, n37899, n232, n38278, n37898, 
        n159, n38277, n37897, n37896;
    wire [23:0]n63;
    wire [23:0]n64;
    
    wire n36564, n45, n36563;
    wire [9:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(26[22:30])
    
    wire n713, n37895, n616, n37894;
    wire [31:0]n66;
    
    wire n519, n37893, n17_c, n86, n422, n37892, n325, n37891;
    wire [22:0]n1799;
    
    wire n38275, n228, n37890;
    wire [31:0]n67;
    
    wire n116, n1695, n38_adj_3370, n131, n36900;
    wire [21:0]n13113;
    
    wire n36901;
    wire [22:0]n12579;
    
    wire n36899, n38274;
    wire [20:0]n8212;
    
    wire n37889, n37888, n37887, n37886, n38273, n23_c, n37885, 
        n38272, n37884, n37883, n38271, n36898, n38270, n37882, 
        n37881, n37880, n38269, n36897, n37879, n38268, n37878, 
        n36896, n37877, n37876, n38267, n710, n37875, n43, n36562, 
        n613, n37874, n516, n37873, n36895, n36894, n419_adj_3371, 
        n37872, n38266, n38265, n322, n37871, n36893, n225, n37870, 
        n38264, n36892, n35, n128, n38263, n41_adj_3372, n36561;
    wire [21:0]n8188;
    
    wire n37869, n36891, n38262, n37868, n213, n36890, n38261, 
        n37867, n36889, n38260, n37866, n704, n36888, n521, n38259, 
        n37865, n607, n36887, n448, n38258, n37864, n510, n36886, 
        n375, n38257, n37863, n413_c, n36885, n302, n38256, n37862, 
        n316, n36884, n229, n38255, n37861, n219, n36883, n156, 
        n38254, n37860, n29_c, n122, n310, n14, n83, n37859;
    wire [10:0]n16318;
    wire [9:0]n16424;
    
    wire n36882;
    wire [22:0]n1798;
    
    wire n38252, n37858, n1691, n36881, n38251, n37857, n36880, 
        n38250;
    wire [31:0]n69;
    
    wire n37856, n407, n36879, n38249, n37855, n740, n36878, n38248, 
        n707, n37854, n643, n36877, n38247, n610, n37853, n546, 
        n36876, n38246, n513, n37852, n449_adj_3374, n36875, n38245, 
        n416_c, n37851, n352, n36874, n38244, n319, n37850, n255, 
        n36873, n38243, n222, n37849, n65, n158, n38242, n32_adj_3375, 
        n125;
    wire [20:0]n13598;
    
    wire n36872, n36871, n38241;
    wire [22:0]n8163;
    
    wire n37848, n37847, n36870, n504, n38240, n37846, n36869, 
        n38239, n37845, n36868, n39_adj_3376, n36560, n38238, n37844, 
        n36867, n38237, n37843, n36866, n518, n38236, n37842, 
        n36865, n445, n38235, n37841, n36864, n37_adj_3378, n36559, 
        n372, n38234, n37840, n36863, n601_adj_3380, n299, n38233, 
        n37839, n36862, n226, n38232, n37838, n36861, n153, n38231, 
        n37837;
    wire [24:0]\PID_CONTROLLER.err_31__N_2816 ;
    wire [24:0]n70;
    
    wire n36670, n35_adj_3382, n36558, n36860, n11_c, n80, n37836, 
        n36669, n33_adj_3383, n36557, n36859;
    wire [22:0]n1797;
    
    wire n38229, n37835, n1687, n698, n38228, n37834, n36858, 
        n38227, n37833, n707_adj_3385, n36857, n38226, n704_adj_3386, 
        n37832, n31_adj_3387, n36556, n610_adj_3388, n36856, n38225, 
        n607_adj_3389, n37831, n36668, n29_adj_3391, n36555, n513_adj_3393, 
        n36855, n38224, n510_adj_3394, n37830, n416_adj_3395, n36854, 
        n38223, n413_adj_3396, n37829, n319_adj_3397, n36853, n38222, 
        n316_adj_3398, n37828, n27, n36554, n222_adj_3399, n36852, 
        n38221, n219_adj_3400, n37827, n36667, n25, n36553, n32_adj_3402, 
        n125_adj_3403, n38220, n29_adj_3404, n122_adj_3405;
    wire [19:0]n14039;
    
    wire n36851, n38219;
    wire [23:0]n8137;
    
    wire n37826, n37825, n36850, n38218, n37824, n36849, n36666, 
        n23_adj_3407, n36552, n38217, n37823, n36848, n21_c, n36551, 
        n167, n86_adj_3409, n38216, n37822, n36847, n264, n38215, 
        n37821, n36846, n38214, n36845, n19_c, n36550, n37820, 
        n36665, n17_adj_3411, n36549, n515, n38213, n36844, n37819, 
        n15_adj_3414, n36548, n442, n38212, n37818, n36843, n361, 
        n369, n38211, n37817, n36842, n296, n38210, n36841, n13_adj_3415, 
        n36547, n37816, n458_c, n36664, n11_adj_3418, n36546, n223, 
        n38209, n36840, n37815, n555, n41482, n24435, n24433, 
        n24432, n652, n749, n140, n47, n237, n334, n431, n528_adj_3419, 
        n625, n722, n9_adj_3420, n36545, n150, n38208, n161, n68, 
        n37814, n8_adj_3422, n77, n37813, n37812, n37811, n37810, 
        n36839;
    wire [22:0]n1796;
    
    wire n38206, n36838, n36663, n1683, n701, n37809, n710_adj_3424, 
        n36837, n36662;
    wire [33:0]n282;
    
    wire n38205, n613_adj_3426, n36836, n36661, n604, n37808, n516_adj_3428, 
        n36835, n36660, n7_adj_3430, n36544, n36659;
    wire [31:0]\PID_CONTROLLER.result_31__N_2994 ;
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(25[23:29])
    
    wire n38204, n74, n507, n37807, n419_adj_3432, n36834, n36658, 
        n5_adj_3434, n36543, n322_adj_3436, n36833, n3_adj_3437, n36542, 
        n38203, n410, n37806, n5_adj_3439, n38202, n36657, n225_adj_3442, 
        n36832, n313, n37805, n38201, n36656, n147, n35_adj_3445, 
        n128_adj_3446, n36655, n220, n216, n37804;
    wire [31:0]pwm_23__N_2951;
    
    wire n36541, n36654, n36540, n293, n26_adj_3450, n119;
    wire [24:0]n8110;
    
    wire n37803, n37802, n37801, n37800, n37799;
    wire [8:0]n16509;
    
    wire n36831, n36830, n38200, n36829, n36653, n37798, n743, 
        n36828, n36652, n38199, n36651, n646, n36827, n36539, 
        n37797, n36650, n366, n38198, n549, n36826, n37796, n36649, 
        n36538, n439, n38197, n37795, n452_adj_3461, n36825, n36648, 
        n38196, n37794, n355, n36824, n36537, n36647, n37793, 
        n512, n38195, n38194, n258, n36823, n38193, n38192, n38191, 
        n38190, n38189, n38188, n38187, n38186, n38185;
    wire [16:0]n15118;
    wire [15:0]n15403;
    
    wire n38184, n38183, n37792, n36536;
    wire [18:0]n14438;
    
    wire n36822, n38182, n38181, n38180, n38179, n38178, n38177, 
        n38176, n38175, n38174, n38173, n38172, n38171, n38170, 
        n38169;
    wire [7:0]n16575;
    wire [6:0]n16624;
    
    wire n38168, n38167, n38166, n37791, n38165, n37790, n38164, 
        n36821, n38163, n37789, n38162, n37788;
    wire [14:0]n15644;
    
    wire n38161, n37787, n38160, n36820, n37786, n38159, n37785, 
        n36535, n37784, n38158, n37783, n37782, n36534, n38157, 
        n37781, n38156, n37780, n38155, n38154;
    wire [25:0]n8082;
    
    wire n37779, n37778, n36819, n37777, n36646, n38153, n37776, 
        n37775, n725, n38152, n628, n38151, n531, n38150, n434, 
        n38149, n337, n38148, n240, n38147, n50, n143;
    wire [5:0]n16633;
    
    wire n43817, n658, n38146;
    wire [4:0]n16641;
    
    wire n558, n38145, n37774, n37773, n37772, n37771, n37770, 
        n37769, n37768, n37767, n464, n38144, n37766, n37765;
    wire [2:0]n16654;
    
    wire n370_adj_3471, n38143, n37764, n37763, n37762, n36645, 
        n36533, n276, n38142, n36532, n46507, n28960, n182, n36644, 
        n37761;
    wire [13:0]n15854;
    
    wire n38141, n695, n37760, n598_adj_3477, n37759, n38140, n501, 
        n37758, n36643, n36818, n38139, n404, n37757, n307_adj_3479, 
        n37756, n210, n37755, n20_adj_3480, n113, n38138;
    wire [26:0]n8053;
    
    wire n37754, n37753, n37752, n38137, n37751, n19326, n881_adj_3481, 
        n16802, n17_adj_3482, n43915, n37750, n38136, n37749, n37748, 
        n36642, n37747, n36641, n38135, n37746;
    wire [8:0]n7069;
    wire [22:0]n1804;
    
    wire n1711, n38418, n38134, n36640;
    wire [22:0]n1803;
    
    wire n1707, n38417, n728, n38133, n37745, n36639, n37744, 
        n631, n38132, n534, n38131, n37743, n37742, n36638, n37741, 
        n37740, n36637;
    wire [22:0]n1802;
    
    wire n1703, n38416, n437, n38130, n36636, n36635, n37739, 
        n1699, n38415, n340, n38129, n37738, n36634, n37737, n243, 
        n38128, n37736, n53_adj_3492, n146, n36817, n37735, n692, 
        n37734, n36633, n595_adj_3495, n37733, n498, n37732, n36632, 
        n38414, n752, n38127, n38413, n38126, n36631, n401, n37731, 
        n36816, n38125, n304_adj_3498, n37730, n207, n37729, n36630, 
        n38412, n17_adj_3500, n110, n38124;
    wire [27:0]n8023;
    
    wire n37728, n37727, n38123, n37726, n37725, n37724, n38411, 
        n37723, n38122, n37722, n37721, n37720, n37719, n37718;
    wire [20:0]n8476;
    wire [19:0]n9331;
    
    wire n38410, n37717, n38409, n37716, n37715, n38408, n37714, 
        n37713, n38407, n36815, n37712, n36814, n36813, n36629;
    wire [12:0]n16035;
    
    wire n38121, n37711, n38406, n36812, n36628, n38120, n36811, 
        n38119, n37710, n36810, n38405, n37709, n713_adj_3503, n36809, 
        n36627, n38118, n37708, n616_adj_3505, n36808, n36626, n38404, 
        n38117, n519_adj_3507, n36807, n689, n37707, n36625, n38116, 
        n422_adj_3509, n36806, n36624, n38403, n592_adj_3511, n37706, 
        n325_adj_3512, n36805, n38115, n36623, n495, n37705, n228_adj_3514, 
        n36804, n36622, n731, n38114, n38_adj_3517, n131_adj_3518, 
        PHASES_5__N_3046, n36621;
    wire [23:0]n852;
    wire [23:0]n73;
    
    wire n36620, n398, n37704, n38402, n634, n38113, n301_adj_3522, 
        n37703, n204, n37702;
    wire [17:0]n14797;
    
    wire n36803, n36619, n537, n38112, n36802, n440, n38111, n14_adj_3525, 
        n107;
    wire [28:0]n7992;
    
    wire n37701, n36618, n38401, n37700, n36801, n36617, n343, 
        n38110, n37699, n36616, n37698, n246, n38109, n36615, 
        n38400, n37697, n56, n149, n37696, n36800, n37695;
    wire [11:0]n16189;
    
    wire n38108, n38107, n37694, n36799, n38399, n38106, n37693, 
        n37692, n36798, n37691, n38398, n37690, n38105, n36614, 
        n38397, n37689, n38104, n36797, n37688;
    wire [8:0]n75;
    wire [8:0]pwm_count;   // verilog/motorControl.v(55[13:22])
    
    wire n38103, n36613, n734, n38102, n37687, n545, n38396, n637, 
        n38101, n37686, n36796, n540, n38100, n37685, n472, n38395, 
        n36795, n37684, n37683, n443_adj_3536, n38099, n36612, n37682, 
        n346, n38098, n36794, n36611, n399, n38394, n37681;
    wire [0:0]n5790;
    wire [29:0]n6546;
    
    wire n37192;
    wire [55:0]n76;
    
    wire n37191, n249, n38097, n36793, n37680, n37190, n686, n37679, 
        n37189, n36792, n59, n152, n37188, n589_adj_3541, n37678, 
        n37187, n38096, n492, n37677, n716, n36791, n326, n38393, 
        n37186, n38095, n36610, n395, n37676, n37185, n619, n36790, 
        n38094, n298_adj_3545, n37675, n37184, n522_adj_3547, n36789, 
        n253, n38392, n201, n37674, n37183, n37182, n11_adj_3548, 
        n104, n38093, n37181, n37180, n37179, n425_adj_3549, n36788, 
        n36609;
    wire [0:0]n7065;
    wire [29:0]n7960;
    
    wire n37673, n37178, n38092;
    wire [55:0]n191;
    
    wire n37672, n37177, n737, n38091, n180_adj_3552, n38391, n37176, 
        n37671, n328_adj_3553, n36787, n37175, n640, n38090, n37174, 
        n37670, n35_adj_3556, n107_adj_3557, n37173, n231_adj_3558, 
        n36786, n543, n38089, n446_adj_3559, n38088, n37172, n37669, 
        n349, n38087, n37171, n41_adj_3563, n134_adj_3564, n36608, 
        n37170;
    wire [21:0]n8452;
    
    wire n38390, n38389, n252, n38086, n37668, n37169, n62, n155, 
        n37667, n38085, n680, n37168, n36785, n583, n37167, n37666, 
        n38388, n38084, n486, n37166, n389, n37165, n37665, n38083, 
        n292, n37164, n36784, n38082, n195, n37163, n37664, n5_adj_3578, 
        n98, n38081, n746, n36783, n38387, n37663, n38080, n649, 
        n36782, n36607, n37662, n38079, n552, n36781, n37661, 
        n36606, n37660, n38078, n37659, n38386, n36605, n38077, 
        n37658, n455_adj_3588, n36780;
    wire [28:0]n7764;
    
    wire n37155, n37154, n37657, n37656, n38076, n37153, n37152, 
        n37655, n36604, n358, n36779, n37151, n38385, n38075, 
        n37654, n37150, n36603, n37149, n38074, n37653, n37148, 
        n37652, n37147, n261, n36778, n38384, n38073, n36602, 
        n37146, n37651, n37145, n38383, n38072, n37650, n71, n164, 
        n38071, n37144, n680_adj_3597, n37649, n37143, n583_adj_3598, 
        n37648, n37142, n36601, n37141, n36600, n38382, n38070, 
        n486_adj_3601, n37647, n389_adj_3603, n37646, n38069, n38381, 
        n37140, n292_adj_3604, n37645, n38380, n38068, n195_adj_3605, 
        n37644, n37139, n5_adj_3607, n98_adj_3608, n37138, n36599;
    wire [18:0]n10122;
    
    wire n37643, n37137, n38067, n37642, n37136, n37641, n28668, 
        n38066, n38379, n38065, n37640, n37135, n37134, n37639, 
        n37133, n38378, n683, n37132, n37638, n586, n37131, n37637, 
        n489, n37130;
    wire [6:0]n8443;
    wire [5:0]n9323;
    
    wire n752_adj_3611, n38064, n37636, n655, n38063, n392, n37129, 
        n295_adj_3612, n37128, n37635, n558_adj_3613, n38062, n37634, 
        n198, n37127, n8_adj_3614, n101;
    wire [27:0]n9129;
    
    wire n37126, n37633, n38377, n461_c, n38061, n37125, n37632, 
        n37631;
    wire [31:0]n79;
    
    wire n36772, n37124, n36771, n37630, n37123, n38376, n37122, 
        n364, n38060, n37121, n36770, n37629, n37120, n267, n38059, 
        n37119, n36769, n38375, n37628, n37118, n86_adj_3617, n170_adj_3618, 
        n37627, n37117;
    wire [7:0]n8433;
    
    wire n38058, n37626, n37116, n36768, n749_adj_3619, n38057, 
        n37115, n37625, n37114, n36767, n37113, n536, n38374, 
        n652_adj_3621, n38056, n44226, n658_adj_3622, n37624, n37112;
    wire [4:0]n10115;
    
    wire n564, n37623, n555_adj_3623, n38055;
    wire [3:0]n10850;
    
    wire n464_adj_3624, n37622, n37111, n37110, n36766, n463_c, 
        n38373, n458_adj_3626, n38054, n370_adj_3627, n37621, n37109, 
        n361_adj_3628, n38053, n37108, n276_adj_3629, n37620, n37107, 
        n36765, n37106, n264_adj_3630, n38052, n182_adj_3631, n390, 
        n38372, n37105, n686_adj_3632, n37104, n74_adj_3633, n167_adj_3634, 
        n36764;
    wire [17:0]n10856;
    
    wire n37619, n589_adj_3635, n37103, n37618, n492_adj_3636, n37102, 
        n36763;
    wire [8:0]n8422;
    
    wire n38051, n37617, n395_adj_3637, n37101, n38050, n37616, 
        n36762, n298_adj_3638, n37100, n201_adj_3639, n37099, n11_adj_3640, 
        n104_adj_3641, n317, n38371, n37615, n37614, n36761, n746_adj_3642, 
        n38049, n244_adj_3644, n38370, n37613;
    wire [13:0]n13260;
    wire [12:0]n13738;
    
    wire n37098, n37097, n37096, n37612, n37611, n649_adj_3645, 
        n38048, n552_adj_3646, n38047, n37095, n37610, n37609, n37608, 
        n37094, n37093, n37607, n37092, n455_adj_3647, n38046, n37091, 
        n36760, n171_adj_3649, n38369, n358_adj_3650, n38045, n37606, 
        n37605, n37604, n37090, n261_adj_3651, n38044, n37603, n37089, 
        n98_adj_3652, n37088, n37602, n71_adj_3653, n164_adj_3654, 
        n37087;
    wire [16:0]n11535;
    
    wire n37601, n37086, n37600, n38367;
    wire [9:0]n8410;
    
    wire n38043, n37599, n36759, n38042, n37598;
    wire [26:0]n9933;
    
    wire n37085, n37084, n37597, n37083, n38041, n37596, n37082, 
        n38366, n37081, n743_adj_3655, n38040, n37595, n37080, n36758, 
        n37079, n646_adj_3656, n38039, n37594, n37078, n36757, n38365, 
        n37077, n549_adj_3657, n38038, n37593, n37076, n36756, n37075, 
        n452_adj_3658, n38037, n37592, n37074, n36755, n38364, n37591, 
        n37073, n355_adj_3659, n38036, n37590, n37072, n37071, n37589, 
        n37070, n38363, n258_adj_3660, n38035, n37588;
    wire [9:0]n82;
    
    wire n55_adj_3661, n37069, n37587, n37068, n38362, n68_adj_3662, 
        n161_adj_3663, n37586;
    wire [10:0]n8397;
    
    wire n38034, n37067, n37585, n37066, n38033, n37065, n38361, 
        n689_adj_3664, n37064;
    wire [15:0]n12161;
    
    wire n37584, n36754, n37583, n592_adj_3665, n37063, n38032, 
        n37582, n495_adj_3666, n37062, n38031, n37581, n398_adj_3667, 
        n37061, n301_adj_3668, n37060, n37580, n204_adj_3669, n37059, 
        n740_adj_3670, n38030, n37579, n14_adj_3671, n107_adj_3672, 
        n36753, n37578;
    wire [11:0]n14172;
    
    wire n37058, n38360, n37057, n37056, n37577, n36752, n37055, 
        n643_adj_3673, n38029, n38359, n37576, n37054, n36751, n37575, 
        n37053, n546_adj_3674, n38028, n37574, n37052, n36750, n449_adj_3675, 
        n38027, n38358, n37573, n37572, n37051, n352_adj_3676, n38026, 
        n37571, n36749, n37570, n37050, n255_adj_3677, n38025, n36748, 
        n37569, n38357, n65_adj_3678, n158_adj_3679, n37049, n37048, 
        n37047;
    wire [14:0]n12736;
    
    wire n37568;
    wire [11:0]n8383;
    
    wire n38024, n37567;
    wire [25:0]n10675;
    
    wire n37046, n36747, n37045, n36746, n38356, n37566, n36745, 
        n38023, n37044, n37565, n37043, n37042, n38022, n37564, 
        n37041, n36744, n38355, n38021, n37563, n37040, n37039, 
        n37562, n37038, n38020, n37037, n37561, n37036, n37560, 
        n737_adj_3680, n38019, n37559, n37035, n36743, n38354, n640_adj_3681, 
        n38018, n37558, n37034, n37033, n37032, n543_adj_3682, n38017, 
        n37557, n37031, n37030, n37029, n37556, n36742, n37555, 
        n446_adj_3683, n38016, n38353, n37028, n37554, n349_adj_3685, 
        n38015, n37027, n252_adj_3686, n38014, n692_adj_3687, n37026, 
        n595_adj_3688, n37025, n38352, n498_adj_3690, n37024, n533, 
        n38351, n62_adj_3692, n155_adj_3693, n401_adj_3694, n37023;
    wire [12:0]n8368;
    
    wire n38013, n38012, n304_adj_3695, n37022, n207_adj_3696, n37021, 
        n17_adj_3697, n110_adj_3698, n36741, n36740;
    wire [10:0]n14564;
    
    wire n37020, n36739, n37019, n37018, n460_c, n38350, n38011, 
        n37017, n38010, n37016, n37015, n37014, n38009, n37013, 
        n387_c, n38349, n38008, n37012, n37011, n734_adj_3700, n38007, 
        n37010, n36738;
    wire [24:0]n11362;
    
    wire n37009, n637_adj_3701, n38006, n314_adj_3703, n38348, n241_adj_3705, 
        n38347, n37008, n168_adj_3707, n38346, n36737, n540_adj_3708, 
        n38005, n443_adj_3709, n38004, n36736, n26_adj_3710, n95, 
        n346_adj_3711, n38003, n37007, n37006, n38344, n249_adj_3712, 
        n38002, n37005, n36735, n37004, n37003, n36734, n37002, 
        n59_adj_3713, n152_adj_3714, n37001, n36733, n37000, n36732, 
        n36999, n38343, n36998, n36731, n36997;
    wire [13:0]n8352;
    
    wire n38001, n38000, n36996, n36995, n719, n36730, n36994, 
        n622, n36729, n36993, n38342, n36992, n525_adj_3715, n36728, 
        n36991, n37999, n695_adj_3716, n36990, n598_adj_3717, n36989, 
        n37998, n428, n36727, n501_adj_3718, n36988, n38341, n404_adj_3719, 
        n36987, n37997, n307_adj_3720, n36986, n331, n36726, n210_adj_3721, 
        n36985, n37996, n20_adj_3722, n113_adj_3723, n234_adj_3724, 
        n36725, n38340;
    wire [9:0]n14916;
    
    wire n36984, n36983, n37995, n36982, n44, n137_adj_3725, n731_adj_3726, 
        n37994, n36981, n38339, n36980, n36979, n634_adj_3727, n37993, 
        n36978, n36977, n36724, n36976, n36723, n36975, n36722, 
        n36721, n537_adj_3728, n37992;
    wire [23:0]n11996;
    
    wire n36974, n36973, n38338, n38337, n36720, n38336, n440_adj_3729, 
        n37991, n36972, n343_adj_3730, n37990, n36971, n246_adj_3731, 
        n37989, n36970, n38335, n36969, n36968, n36967, n56_adj_3732, 
        n149_adj_3733, n36966, n36719, n36718, n36965;
    wire [14:0]n8335;
    
    wire n37988, n36964, n36717, n38334, n36716, n37987, n37986, 
        n36963, n37985, n37507, n36962, n37506, n36715, n36961, 
        n38333, n38332, n36960, n37505, n37984, n36959, n36714, 
        n37504, n37983, n38331, n37503, n36958, n37982, n37502, 
        n37981, n37501, n36957, n37500, n36713, n37499, n38330, 
        n698_adj_3737, n36956, n728_adj_3738, n37980, n38329, n631_adj_3740, 
        n37979, n37498, n601_adj_3741, n36955, n37497, n36712, n504_adj_3743, 
        n36954, n37496, n407_adj_3745, n36953, n530, n38328, n36711, 
        n310_adj_3747, n36952, n37495, n36710, n37494, n213_adj_3750, 
        n36951, n37493, n534_adj_3752, n37978, n23_adj_3753, n116_adj_3754, 
        n36709, n37492;
    wire [8:0]n15230;
    
    wire n36950, n437_adj_3756, n37977, n36949, n36948, n37491, 
        n36947, n340_adj_3758, n37976, n36946, n36708, n457_c, n38327, 
        n243_adj_3760, n37975, n37490, n36945, n36707, n36944, n37489, 
        n37488, n36943, n53_adj_3761, n146_adj_3762, n37487, n36942, 
        n37486, n36706, n384, n38326;
    wire [15:0]n8317;
    
    wire n37974, n37973, n37485, n37484, n37483, n36705, n37482, 
        n37972, n37481, n311_adj_3764, n38325, n37480;
    wire [5:0]PHASES_5__N_2779;
    
    wire n23562, n23622, n15_adj_3765, n23630, n42681, n36704, n37971, 
        n36935, n36934, n36703, n37479, n238_adj_3767, n38324, n36933, 
        n36932, n37970, n37478, n36702, n36931, n36930, n36701, 
        n165_adj_3769, n38323, n37969, n37477, n36929, n37476, n36928, 
        n37968, n36700, n6_adj_3771, n36574, n36927, n37475, n36926, 
        n37967, n37474, n36925, n36699, n36573, n36924, n36698, 
        n36923, n36697, n37966, n23_adj_3772, n92, n37473, n36922, 
        n38321, n38320, n725_adj_3773, n37965, n37472, n36921, n36920, 
        n628_adj_3774, n37964, n36919;
    wire [5:0]PHASES_5__N_3039;
    
    wire n43441, n934, n22379, n37471, n36572, n37470, n19954, 
        n19616, n38319, n37469, n701_adj_3776, n36918, n36696, n531_adj_3777, 
        n37963, n37468, n604_adj_3778, n36917, n42680, n683_adj_3779, 
        n37467, n507_adj_3780, n36916, n434_adj_3781, n37962, n38318, 
        n410_adj_3782, n36915, n36695, n337_adj_3783, n37961, n586_adj_3784, 
        n37466, n313_adj_3785, n36914, n489_adj_3786, n37465, n240_adj_3787, 
        n37960, n216_adj_3788, n36913, n50_adj_3790, n143_adj_3791, 
        n36694, n392_adj_3792, n37464, n26_adj_3793, n119_adj_3794, 
        n38317;
    wire [16:0]n8298;
    
    wire n37959, n295_adj_3797, n37463, n36912, n36571, n583_adj_3800, 
        n36911, n37958, n198_adj_3801, n37462, n510_adj_3802, n36910, 
        n38316, n37957, n8_adj_3803, n101_adj_3804, n437_adj_3805, 
        n36909, n37461, n364_adj_3806, n36908, n37460, n291, n36907, 
        n37459, n36570, n218_adj_3808, n36906, n38315, n145_adj_3809, 
        n36905, n38314, n37956, n37458, n38313, n37955, n37457, 
        n37954, n72, n36569, n37456, n37455, n36904, n36903, n37454, 
        n36902, n37953, n37453, n38312, n37452, n37952, n37951, 
        n38311, n37950, n38310, n38309, n37451, n722_adj_3813, n37949, 
        n38308, n37450, n625_adj_3814, n37948, n37449, n528_adj_3815, 
        n37947, n38307, n37448, n431_adj_3816, n37946, n334_adj_3817, 
        n37945, n38306, n237_adj_3818, n37944, n47_adj_3819, n140_adj_3820, 
        n527, n38305, n37943, n37942, n454, n38304, n37941, n37447, 
        n37940, n381, n38303, n37939, n37938, n308_adj_3821, n38302, 
        n37937, n37936, n235_adj_3822, n38301, n37935, n162, n38300, 
        n20_adj_3823, n89, n38298, n38297, n37934, n38296, n37933, 
        n719_adj_3824, n37932, n38295, n622_adj_3825, n37931, n525_adj_3826, 
        n37930, n38294, n428_adj_3827, n37929, n331_adj_3828, n37928, 
        n38293, n234_adj_3829, n37927, n44_adj_3830, n137_adj_3831, 
        n38292, n37926, n37925, n38291, n37924, n37923, n38290, 
        n37922, n37921, n38289, n37920, n37919, n38288, n37918, 
        n37917, n38287, n37916, n37915, n38286, n716_adj_3832, n37914, 
        n619_adj_3833, n37913, n522_adj_3834, n46606, n13_adj_3842, 
        n7_adj_3843, n11_adj_3844, n13_adj_3845, n17_adj_3846, n47725, 
        n47719, n47733, n47705, n47685, n30_adj_3849, n47743, n48037, 
        n47729, n48283, n47105, n48021, n48437, n48584, n6_adj_3850, 
        n48169, n47661, n24_adj_3851, n47063, n49657, n8_adj_3852, 
        n48385, n47466, n4_adj_3853, n48167, n47093, n49635, n10_adj_3854, 
        n48503, n47468, n48604, n48605, n47067, n48534, n47474, 
        n48600, n50_adj_3855, n19_adj_3856, n17_adj_3857, n7_adj_3858, 
        n13_adj_3859, n4_adj_3860, n48159, n48160, n46986, n47623, 
        n6_adj_3863, n8_adj_3864, n47478, n48187, n18_adj_3866, n44105, 
        n43893, n26_adj_3867, n44113, n43892, n34_adj_3868, n62_adj_3869, 
        n49_adj_3870, n42736, n42695, n44333, n56_adj_3871, n44118, 
        n42629, n20_adj_3872, n16_adj_3873, n10_adj_3874, n12_adj_3875, 
        n14_adj_3876, n13_adj_3877, n18_adj_3878, n5_adj_3879, n47028, 
        n8_adj_3882, n6_adj_3883, n16_adj_3884, n46504, n4_adj_3885, 
        n48163, n48164, n24_adj_3886, n22_adj_3887, n23_adj_3888, 
        n21_adj_3889, n47018, n47016, n48465, n47476, n44367, n48598, 
        n47655, n56_adj_3891, n60, pwm_23__N_2950, n48183, n17_adj_3892, 
        n42627, n14_adj_3893, n15_adj_3894, n6_adj_3895, n13_adj_3896, 
        n7_adj_3897, n19_adj_3898, n18_adj_3899, n24_adj_3900, n5_adj_3901, 
        n46955, n4_adj_3904, n48157, n48158, n10_adj_3905, n22_adj_3906, 
        n12_adj_3907, n16_adj_3908, n26_adj_3909, n46613, n25_adj_3910, 
        n6_adj_3911, n48349, n48350, n46947, n47486, n48140, n20_adj_3913, 
        n48191, n46608, n43470, n878, n43468, n46609, n43907, 
        n42708, n880, n43507, n46611, n20463, n4_adj_3914, n902_adj_3915, 
        n20_adj_3918, n26_adj_3919, n24_adj_3920, n28_adj_3921, n23_adj_3922, 
        n46593, n12_adj_3923, n4_adj_3924, n6_adj_3925, n8_adj_3926, 
        n8_adj_3927, n4_adj_3928, n36197, n38421, n7_adj_3929, n6_adj_3930, 
        n8_adj_3931, n8_adj_3932, n36328, n8_adj_3933, n18_adj_3934, 
        n24_adj_3935, n22_adj_3936, n26_adj_3937, n44028, n11_adj_3938, 
        n9_adj_3939, n17_adj_3940, n47835, n47831, n47169, n49860, 
        n47845, n47815, n47216, n49848, n10_adj_3941, n30_adj_3942, 
        n5_adj_3943, n47855, n47851, n47258, n48085, n48461, n47821, 
        n48297, n48532, n48622, n6_adj_3944, n47403, n24_adj_3945, 
        n48177, n47185, n49813, n47923, n47452, n4_adj_3946, n48171, 
        n48172, n8_adj_3947, n47155, n6_adj_3948, n16_adj_3949, n47159, 
        n48253, n47462, n48509, n4_adj_3950, n48175, n47220, n48487, 
        n47454, n48602, n48603, n47783, n48387, n47460, n48510, 
        n48507, n36343, n7_adj_3951, n20375;
    
    SB_LUT4 add_3095_5_lut (.I0(GND_net), .I1(n8278[2]), .I2(n425), .I3(n37911), 
            .O(n8257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_5 (.CI(n37911), .I0(n8278[2]), .I1(n425), .CO(n37912));
    SB_CARRY Kd_delay_counter_1047_add_4_6 (.CI(n37445), .I0(GND_net), .I1(Kd_delay_counter[4]), 
            .CO(n37446));
    SB_LUT4 Kd_delay_counter_1047_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[3]), .I3(n37444), .O(n57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1047_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1047_add_4_5 (.CI(n37444), .I0(GND_net), .I1(Kd_delay_counter[3]), 
            .CO(n37445));
    SB_LUT4 mult_14_add_1215_10_lut (.I0(GND_net), .I1(n1801[7]), .I2(GND_net), 
            .I3(n38284), .O(n1800[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_4_lut (.I0(GND_net), .I1(n8278[1]), .I2(n328), .I3(n37910), 
            .O(n8257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_4 (.CI(n37910), .I0(n8278[1]), .I1(n328), .CO(n37911));
    SB_LUT4 Kd_delay_counter_1047_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[2]), .I3(n37443), .O(n57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1047_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_3_lut (.I0(GND_net), .I1(n8278[0]), .I2(n231), .I3(n37909), 
            .O(n8257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1047_add_4_4 (.CI(n37443), .I0(GND_net), .I1(Kd_delay_counter[2]), 
            .CO(n37444));
    SB_LUT4 Kd_delay_counter_1047_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[1]), .I3(n37442), .O(n57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1047_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_10 (.CI(n38284), .I0(n1801[7]), .I1(GND_net), 
            .CO(n38285));
    SB_CARRY add_3095_3 (.CI(n37909), .I0(n8278[0]), .I1(n231), .CO(n37910));
    SB_LUT4 add_3095_2_lut (.I0(GND_net), .I1(n41), .I2(n134), .I3(GND_net), 
            .O(n8257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1047_add_4_3 (.CI(n37442), .I0(GND_net), .I1(Kd_delay_counter[1]), 
            .CO(n37443));
    SB_LUT4 Kd_delay_counter_1047_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[0]), .I3(VCC_net), .O(n57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1047_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_9_lut (.I0(GND_net), .I1(n1801[6]), .I2(GND_net), 
            .I3(n38283), .O(n1800[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_2 (.CI(GND_net), .I0(n41), .I1(n134), .CO(n37909));
    SB_LUT4 add_3094_21_lut (.I0(GND_net), .I1(n8257[18]), .I2(GND_net), 
            .I3(n37908), .O(n8235[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_20_lut (.I0(GND_net), .I1(n8257[17]), .I2(GND_net), 
            .I3(n37907), .O(n8235[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_20 (.CI(n37907), .I0(n8257[17]), .I1(GND_net), .CO(n37908));
    SB_CARRY Kd_delay_counter_1047_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(Kd_delay_counter[0]), .CO(n37442));
    SB_LUT4 add_3094_19_lut (.I0(GND_net), .I1(n8257[16]), .I2(GND_net), 
            .I3(n37906), .O(n8235[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_19 (.CI(n37906), .I0(n8257[16]), .I1(GND_net), .CO(n37907));
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n61[3]), 
            .I3(n36567), .O(n58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_5 (.CI(n36567), .I0(GND_net), .I1(n61[3]), 
            .CO(n36568));
    SB_CARRY mult_14_add_1215_9 (.CI(n38283), .I0(n1801[6]), .I1(GND_net), 
            .CO(n38284));
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n61[2]), 
            .I3(n36566), .O(n58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_18_lut (.I0(GND_net), .I1(n8257[15]), .I2(GND_net), 
            .I3(n37905), .O(n8235[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_8_lut (.I0(GND_net), .I1(n1801[5]), .I2(n524), 
            .I3(n38282), .O(n1800[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_18 (.CI(n37905), .I0(n8257[15]), .I1(GND_net), .CO(n37906));
    SB_CARRY mult_14_add_1215_8 (.CI(n38282), .I0(n1801[5]), .I1(n524), 
            .CO(n38283));
    SB_LUT4 add_3094_17_lut (.I0(GND_net), .I1(n8257[14]), .I2(GND_net), 
            .I3(n37904), .O(n8235[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_4 (.CI(n36566), .I0(GND_net), .I1(n61[2]), 
            .CO(n36567));
    SB_CARRY add_3094_17 (.CI(n37904), .I0(n8257[14]), .I1(GND_net), .CO(n37905));
    SB_LUT4 mult_14_add_1215_7_lut (.I0(GND_net), .I1(n1801[4]), .I2(n451), 
            .I3(n38281), .O(n1800[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_16_lut (.I0(GND_net), .I1(n8257[13]), .I2(GND_net), 
            .I3(n37903), .O(n8235[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_16 (.CI(n37903), .I0(n8257[13]), .I1(GND_net), .CO(n37904));
    SB_CARRY mult_14_add_1215_7 (.CI(n38281), .I0(n1801[4]), .I1(n451), 
            .CO(n38282));
    SB_LUT4 add_3094_15_lut (.I0(GND_net), .I1(n8257[12]), .I2(GND_net), 
            .I3(n37902), .O(n8235[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_6_lut (.I0(GND_net), .I1(n1801[3]), .I2(n378), 
            .I3(n38280), .O(n1800[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_15 (.CI(n37902), .I0(n8257[12]), .I1(GND_net), .CO(n37903));
    SB_CARRY mult_14_add_1215_6 (.CI(n38280), .I0(n1801[3]), .I1(n378), 
            .CO(n38281));
    SB_LUT4 mult_14_add_1215_5_lut (.I0(GND_net), .I1(n1801[2]), .I2(n305), 
            .I3(n38279), .O(n1800[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_14_lut (.I0(GND_net), .I1(n8257[11]), .I2(GND_net), 
            .I3(n37901), .O(n8235[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_14 (.CI(n37901), .I0(n8257[11]), .I1(GND_net), .CO(n37902));
    SB_LUT4 add_3094_13_lut (.I0(GND_net), .I1(n8257[10]), .I2(GND_net), 
            .I3(n37900), .O(n8235[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_13 (.CI(n37900), .I0(n8257[10]), .I1(GND_net), .CO(n37901));
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n61[1]), 
            .I3(n36565), .O(n58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_12_lut (.I0(GND_net), .I1(n8257[9]), .I2(GND_net), 
            .I3(n37899), .O(n8235[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_3 (.CI(n36565), .I0(GND_net), .I1(n61[1]), 
            .CO(n36566));
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n61[0]), 
            .I3(VCC_net), .O(n58[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_12 (.CI(n37899), .I0(n8257[9]), .I1(GND_net), .CO(n37900));
    SB_CARRY mult_14_add_1215_5 (.CI(n38279), .I0(n1801[2]), .I1(n305), 
            .CO(n38280));
    SB_LUT4 mult_14_add_1215_4_lut (.I0(GND_net), .I1(n1801[1]), .I2(n232), 
            .I3(n38278), .O(n1800[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n61[0]), 
            .CO(n36565));
    SB_LUT4 add_3094_11_lut (.I0(GND_net), .I1(n8257[8]), .I2(GND_net), 
            .I3(n37898), .O(n8235[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_4 (.CI(n38278), .I0(n1801[1]), .I1(n232), 
            .CO(n38279));
    SB_CARRY add_3094_11 (.CI(n37898), .I0(n8257[8]), .I1(GND_net), .CO(n37899));
    SB_LUT4 mult_14_add_1215_3_lut (.I0(GND_net), .I1(n1801[0]), .I2(n159), 
            .I3(n38277), .O(n1800[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_10_lut (.I0(GND_net), .I1(n8257[7]), .I2(GND_net), 
            .I3(n37897), .O(n8235[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_10 (.CI(n37897), .I0(n8257[7]), .I1(GND_net), .CO(n37898));
    SB_LUT4 add_3094_9_lut (.I0(GND_net), .I1(n8257[6]), .I2(GND_net), 
            .I3(n37896), .O(n8235[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n64[23]), 
            .I3(n36564), .O(n63[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_9 (.CI(n37896), .I0(n8257[6]), .I1(GND_net), .CO(n37897));
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[22]), .I3(n36563), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3094_8_lut (.I0(GND_net), .I1(n8257[5]), .I2(n713), .I3(n37895), 
            .O(n8235[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_8 (.CI(n37895), .I0(n8257[5]), .I1(n713), .CO(n37896));
    SB_LUT4 add_3094_7_lut (.I0(GND_net), .I1(n8257[4]), .I2(n616), .I3(n37894), 
            .O(n8235[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_7 (.CI(n37894), .I0(n8257[4]), .I1(n616), .CO(n37895));
    SB_CARRY mult_14_add_1215_3 (.CI(n38277), .I0(n1801[0]), .I1(n159), 
            .CO(n38278));
    SB_LUT4 sub_11_inv_0_i32_1_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[26]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3094_6_lut (.I0(GND_net), .I1(n8257[3]), .I2(n519), .I3(n37893), 
            .O(n8235[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_2_lut (.I0(GND_net), .I1(n17_c), .I2(n86), 
            .I3(GND_net), .O(n1800[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_6 (.CI(n37893), .I0(n8257[3]), .I1(n519), .CO(n37894));
    SB_LUT4 add_3094_5_lut (.I0(GND_net), .I1(n8257[2]), .I2(n422), .I3(n37892), 
            .O(n8235[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_5 (.CI(n37892), .I0(n8257[2]), .I1(n422), .CO(n37893));
    SB_CARRY mult_14_add_1215_2 (.CI(GND_net), .I0(n17_c), .I1(n86), .CO(n38277));
    SB_LUT4 add_3094_4_lut (.I0(GND_net), .I1(n8257[1]), .I2(n325), .I3(n37891), 
            .O(n8235[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_4 (.CI(n37891), .I0(n8257[1]), .I1(n325), .CO(n37892));
    SB_LUT4 mult_14_add_1214_24_lut (.I0(GND_net), .I1(n1800[21]), .I2(GND_net), 
            .I3(n38275), .O(n1799[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_3_lut (.I0(GND_net), .I1(n8257[0]), .I2(n228), .I3(n37890), 
            .O(n8235[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_3 (.CI(n37890), .I0(n8257[0]), .I1(n228), .CO(n37891));
    SB_LUT4 mult_12_i79_2_lut (.I0(\Kd[1] ), .I1(n67[6]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i79_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1214_24 (.CI(n38275), .I0(n1800[21]), .I1(GND_net), 
            .CO(n1695));
    SB_LUT4 add_3094_2_lut (.I0(GND_net), .I1(n38_adj_3370), .I2(n131), 
            .I3(GND_net), .O(n8235[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_2 (.CI(GND_net), .I0(n38_adj_3370), .I1(n131), .CO(n37890));
    SB_CARRY add_3276_20 (.CI(n36900), .I0(n13113[17]), .I1(GND_net), 
            .CO(n36901));
    SB_LUT4 add_3276_19_lut (.I0(GND_net), .I1(n13113[16]), .I2(GND_net), 
            .I3(n36899), .O(n12579[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_23_lut (.I0(GND_net), .I1(n1800[20]), .I2(GND_net), 
            .I3(n38274), .O(n1799[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_22_lut (.I0(GND_net), .I1(n8235[19]), .I2(GND_net), 
            .I3(n37889), .O(n8212[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_21_lut (.I0(GND_net), .I1(n8235[18]), .I2(GND_net), 
            .I3(n37888), .O(n8212[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_21 (.CI(n37888), .I0(n8235[18]), .I1(GND_net), .CO(n37889));
    SB_LUT4 add_3093_20_lut (.I0(GND_net), .I1(n8235[17]), .I2(GND_net), 
            .I3(n37887), .O(n8212[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_20 (.CI(n37887), .I0(n8235[17]), .I1(GND_net), .CO(n37888));
    SB_CARRY mult_14_add_1214_23 (.CI(n38274), .I0(n1800[20]), .I1(GND_net), 
            .CO(n38275));
    SB_LUT4 add_3093_19_lut (.I0(GND_net), .I1(n8235[16]), .I2(GND_net), 
            .I3(n37886), .O(n8212[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_22_lut (.I0(GND_net), .I1(n1800[19]), .I2(GND_net), 
            .I3(n38273), .O(n1799[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_19 (.CI(n37886), .I0(n8235[16]), .I1(GND_net), .CO(n37887));
    SB_CARRY mult_14_add_1214_22 (.CI(n38273), .I0(n1800[19]), .I1(GND_net), 
            .CO(n38274));
    SB_LUT4 mult_12_i16_2_lut (.I0(\Kd[0] ), .I1(n67[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_c));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3093_18_lut (.I0(GND_net), .I1(n8235[15]), .I2(GND_net), 
            .I3(n37885), .O(n8212[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_19 (.CI(n36899), .I0(n13113[16]), .I1(GND_net), 
            .CO(n36900));
    SB_LUT4 mult_14_add_1214_21_lut (.I0(GND_net), .I1(n1800[18]), .I2(GND_net), 
            .I3(n38272), .O(n1799[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_18 (.CI(n37885), .I0(n8235[15]), .I1(GND_net), .CO(n37886));
    SB_LUT4 add_3093_17_lut (.I0(GND_net), .I1(n8235[14]), .I2(GND_net), 
            .I3(n37884), .O(n8212[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n36563), .I0(GND_net), .I1(n64[22]), 
            .CO(n36564));
    SB_CARRY add_3093_17 (.CI(n37884), .I0(n8235[14]), .I1(GND_net), .CO(n37885));
    SB_CARRY mult_14_add_1214_21 (.CI(n38272), .I0(n1800[18]), .I1(GND_net), 
            .CO(n38273));
    SB_LUT4 add_3093_16_lut (.I0(GND_net), .I1(n8235[13]), .I2(GND_net), 
            .I3(n37883), .O(n8212[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_20_lut (.I0(GND_net), .I1(n1800[17]), .I2(GND_net), 
            .I3(n38271), .O(n1799[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_16 (.CI(n37883), .I0(n8235[13]), .I1(GND_net), .CO(n37884));
    SB_LUT4 add_3276_18_lut (.I0(GND_net), .I1(n13113[15]), .I2(GND_net), 
            .I3(n36898), .O(n12579[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_20 (.CI(n38271), .I0(n1800[17]), .I1(GND_net), 
            .CO(n38272));
    SB_LUT4 mult_14_add_1214_19_lut (.I0(GND_net), .I1(n1800[16]), .I2(GND_net), 
            .I3(n38270), .O(n1799[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_15_lut (.I0(GND_net), .I1(n8235[12]), .I2(GND_net), 
            .I3(n37882), .O(n8212[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_19 (.CI(n38270), .I0(n1800[16]), .I1(GND_net), 
            .CO(n38271));
    SB_CARRY add_3093_15 (.CI(n37882), .I0(n8235[12]), .I1(GND_net), .CO(n37883));
    SB_LUT4 add_3093_14_lut (.I0(GND_net), .I1(n8235[11]), .I2(GND_net), 
            .I3(n37881), .O(n8212[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_18 (.CI(n36898), .I0(n13113[15]), .I1(GND_net), 
            .CO(n36899));
    SB_CARRY add_3093_14 (.CI(n37881), .I0(n8235[11]), .I1(GND_net), .CO(n37882));
    SB_LUT4 add_3093_13_lut (.I0(GND_net), .I1(n8235[10]), .I2(GND_net), 
            .I3(n37880), .O(n8212[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_13 (.CI(n37880), .I0(n8235[10]), .I1(GND_net), .CO(n37881));
    SB_LUT4 mult_14_add_1214_18_lut (.I0(GND_net), .I1(n1800[15]), .I2(GND_net), 
            .I3(n38269), .O(n1799[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_17_lut (.I0(GND_net), .I1(n13113[14]), .I2(GND_net), 
            .I3(n36897), .O(n12579[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_18 (.CI(n38269), .I0(n1800[15]), .I1(GND_net), 
            .CO(n38270));
    SB_LUT4 add_3093_12_lut (.I0(GND_net), .I1(n8235[9]), .I2(GND_net), 
            .I3(n37879), .O(n8212[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_12 (.CI(n37879), .I0(n8235[9]), .I1(GND_net), .CO(n37880));
    SB_CARRY add_3276_17 (.CI(n36897), .I0(n13113[14]), .I1(GND_net), 
            .CO(n36898));
    SB_LUT4 mult_14_add_1214_17_lut (.I0(GND_net), .I1(n1800[14]), .I2(GND_net), 
            .I3(n38268), .O(n1799[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_11_lut (.I0(GND_net), .I1(n8235[8]), .I2(GND_net), 
            .I3(n37878), .O(n8212[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_16_lut (.I0(GND_net), .I1(n13113[13]), .I2(GND_net), 
            .I3(n36896), .O(n12579[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_17 (.CI(n38268), .I0(n1800[14]), .I1(GND_net), 
            .CO(n38269));
    SB_CARRY add_3093_11 (.CI(n37878), .I0(n8235[8]), .I1(GND_net), .CO(n37879));
    SB_CARRY add_3276_16 (.CI(n36896), .I0(n13113[13]), .I1(GND_net), 
            .CO(n36897));
    SB_LUT4 add_3093_10_lut (.I0(GND_net), .I1(n8235[7]), .I2(GND_net), 
            .I3(n37877), .O(n8212[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_10 (.CI(n37877), .I0(n8235[7]), .I1(GND_net), .CO(n37878));
    SB_LUT4 add_3093_9_lut (.I0(GND_net), .I1(n8235[6]), .I2(GND_net), 
            .I3(n37876), .O(n8212[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_9 (.CI(n37876), .I0(n8235[6]), .I1(GND_net), .CO(n37877));
    SB_LUT4 mult_14_add_1214_16_lut (.I0(GND_net), .I1(n1800[13]), .I2(GND_net), 
            .I3(n38267), .O(n1799[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_8_lut (.I0(GND_net), .I1(n8235[5]), .I2(n710), .I3(n37875), 
            .O(n8212[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_8 (.CI(n37875), .I0(n8235[5]), .I1(n710), .CO(n37876));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[21]), .I3(n36562), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3093_7_lut (.I0(GND_net), .I1(n8235[4]), .I2(n613), .I3(n37874), 
            .O(n8212[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_16 (.CI(n38267), .I0(n1800[13]), .I1(GND_net), 
            .CO(n38268));
    SB_CARRY add_3093_7 (.CI(n37874), .I0(n8235[4]), .I1(n613), .CO(n37875));
    SB_LUT4 add_3093_6_lut (.I0(GND_net), .I1(n8235[3]), .I2(n516), .I3(n37873), 
            .O(n8212[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_6 (.CI(n37873), .I0(n8235[3]), .I1(n516), .CO(n37874));
    SB_LUT4 add_3276_15_lut (.I0(GND_net), .I1(n13113[12]), .I2(GND_net), 
            .I3(n36895), .O(n12579[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_15 (.CI(n36895), .I0(n13113[12]), .I1(GND_net), 
            .CO(n36896));
    SB_LUT4 add_3276_14_lut (.I0(GND_net), .I1(n13113[11]), .I2(GND_net), 
            .I3(n36894), .O(n12579[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_5_lut (.I0(GND_net), .I1(n8235[2]), .I2(n419_adj_3371), 
            .I3(n37872), .O(n8212[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_15_lut (.I0(GND_net), .I1(n1800[12]), .I2(GND_net), 
            .I3(n38266), .O(n1799[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_15 (.CI(n38266), .I0(n1800[12]), .I1(GND_net), 
            .CO(n38267));
    SB_CARRY add_3093_5 (.CI(n37872), .I0(n8235[2]), .I1(n419_adj_3371), 
            .CO(n37873));
    SB_LUT4 mult_14_add_1214_14_lut (.I0(GND_net), .I1(n1800[11]), .I2(GND_net), 
            .I3(n38265), .O(n1799[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_4_lut (.I0(GND_net), .I1(n8235[1]), .I2(n322), .I3(n37871), 
            .O(n8212[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_14 (.CI(n36894), .I0(n13113[11]), .I1(GND_net), 
            .CO(n36895));
    SB_CARRY add_3093_4 (.CI(n37871), .I0(n8235[1]), .I1(n322), .CO(n37872));
    SB_LUT4 add_3276_13_lut (.I0(GND_net), .I1(n13113[10]), .I2(GND_net), 
            .I3(n36893), .O(n12579[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_14 (.CI(n38265), .I0(n1800[11]), .I1(GND_net), 
            .CO(n38266));
    SB_LUT4 add_3093_3_lut (.I0(GND_net), .I1(n8235[0]), .I2(n225), .I3(n37870), 
            .O(n8212[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_13_lut (.I0(GND_net), .I1(n1800[10]), .I2(GND_net), 
            .I3(n38264), .O(n1799[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_3 (.CI(n37870), .I0(n8235[0]), .I1(n225), .CO(n37871));
    SB_CARRY add_3276_13 (.CI(n36893), .I0(n13113[10]), .I1(GND_net), 
            .CO(n36894));
    SB_LUT4 add_3276_12_lut (.I0(GND_net), .I1(n13113[9]), .I2(GND_net), 
            .I3(n36892), .O(n12579[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_13 (.CI(n38264), .I0(n1800[10]), .I1(GND_net), 
            .CO(n38265));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n36562), .I0(GND_net), .I1(n64[21]), 
            .CO(n36563));
    SB_LUT4 add_3093_2_lut (.I0(GND_net), .I1(n35), .I2(n128), .I3(GND_net), 
            .O(n8212[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_12_lut (.I0(GND_net), .I1(n1800[9]), .I2(GND_net), 
            .I3(n38263), .O(n1799[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[20]), .I3(n36561), .O(n41_adj_3372)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_14_add_1214_12 (.CI(n38263), .I0(n1800[9]), .I1(GND_net), 
            .CO(n38264));
    SB_CARRY add_3093_2 (.CI(GND_net), .I0(n35), .I1(n128), .CO(n37870));
    SB_CARRY add_3276_12 (.CI(n36892), .I0(n13113[9]), .I1(GND_net), .CO(n36893));
    SB_CARRY unary_minus_5_add_3_22 (.CI(n36561), .I0(GND_net), .I1(n64[20]), 
            .CO(n36562));
    SB_LUT4 add_3092_23_lut (.I0(GND_net), .I1(n8212[20]), .I2(GND_net), 
            .I3(n37869), .O(n8188[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_11_lut (.I0(GND_net), .I1(n13113[8]), .I2(GND_net), 
            .I3(n36891), .O(n12579[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_11_lut (.I0(GND_net), .I1(n1800[8]), .I2(GND_net), 
            .I3(n38262), .O(n1799[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_22_lut (.I0(GND_net), .I1(n8212[19]), .I2(GND_net), 
            .I3(n37868), .O(n8188[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i144_2_lut (.I0(\Kd[2] ), .I1(n67[6]), .I2(GND_net), 
            .I3(GND_net), .O(n213));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i144_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1214_11 (.CI(n38262), .I0(n1800[8]), .I1(GND_net), 
            .CO(n38263));
    SB_CARRY add_3092_22 (.CI(n37868), .I0(n8212[19]), .I1(GND_net), .CO(n37869));
    SB_CARRY add_3276_11 (.CI(n36891), .I0(n13113[8]), .I1(GND_net), .CO(n36892));
    SB_LUT4 add_3276_10_lut (.I0(GND_net), .I1(n13113[7]), .I2(GND_net), 
            .I3(n36890), .O(n12579[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_10_lut (.I0(GND_net), .I1(n1800[7]), .I2(GND_net), 
            .I3(n38261), .O(n1799[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_21_lut (.I0(GND_net), .I1(n8212[18]), .I2(GND_net), 
            .I3(n37867), .O(n8188[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_10 (.CI(n38261), .I0(n1800[7]), .I1(GND_net), 
            .CO(n38262));
    SB_CARRY add_3092_21 (.CI(n37867), .I0(n8212[18]), .I1(GND_net), .CO(n37868));
    SB_CARRY add_3276_10 (.CI(n36890), .I0(n13113[7]), .I1(GND_net), .CO(n36891));
    SB_LUT4 add_3276_9_lut (.I0(GND_net), .I1(n13113[6]), .I2(GND_net), 
            .I3(n36889), .O(n12579[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_9_lut (.I0(GND_net), .I1(n1800[6]), .I2(GND_net), 
            .I3(n38260), .O(n1799[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_20_lut (.I0(GND_net), .I1(n8212[17]), .I2(GND_net), 
            .I3(n37866), .O(n8188[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_9 (.CI(n38260), .I0(n1800[6]), .I1(GND_net), 
            .CO(n38261));
    SB_CARRY add_3092_20 (.CI(n37866), .I0(n8212[17]), .I1(GND_net), .CO(n37867));
    SB_CARRY add_3276_9 (.CI(n36889), .I0(n13113[6]), .I1(GND_net), .CO(n36890));
    SB_LUT4 add_3276_8_lut (.I0(GND_net), .I1(n13113[5]), .I2(n704), .I3(n36888), 
            .O(n12579[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_8_lut (.I0(GND_net), .I1(n1800[5]), .I2(n521), 
            .I3(n38259), .O(n1799[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_19_lut (.I0(GND_net), .I1(n8212[16]), .I2(GND_net), 
            .I3(n37865), .O(n8188[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_8 (.CI(n38259), .I0(n1800[5]), .I1(n521), 
            .CO(n38260));
    SB_CARRY add_3092_19 (.CI(n37865), .I0(n8212[16]), .I1(GND_net), .CO(n37866));
    SB_CARRY add_3276_8 (.CI(n36888), .I0(n13113[5]), .I1(n704), .CO(n36889));
    SB_LUT4 add_3276_7_lut (.I0(GND_net), .I1(n13113[4]), .I2(n607), .I3(n36887), 
            .O(n12579[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_7_lut (.I0(GND_net), .I1(n1800[4]), .I2(n448), 
            .I3(n38258), .O(n1799[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_18_lut (.I0(GND_net), .I1(n8212[15]), .I2(GND_net), 
            .I3(n37864), .O(n8188[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_7 (.CI(n38258), .I0(n1800[4]), .I1(n448), 
            .CO(n38259));
    SB_CARRY add_3092_18 (.CI(n37864), .I0(n8212[15]), .I1(GND_net), .CO(n37865));
    SB_CARRY add_3276_7 (.CI(n36887), .I0(n13113[4]), .I1(n607), .CO(n36888));
    SB_LUT4 add_3276_6_lut (.I0(GND_net), .I1(n13113[3]), .I2(n510), .I3(n36886), 
            .O(n12579[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_6_lut (.I0(GND_net), .I1(n1800[3]), .I2(n375), 
            .I3(n38257), .O(n1799[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_17_lut (.I0(GND_net), .I1(n8212[14]), .I2(GND_net), 
            .I3(n37863), .O(n8188[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_6 (.CI(n38257), .I0(n1800[3]), .I1(n375), 
            .CO(n38258));
    SB_CARRY add_3092_17 (.CI(n37863), .I0(n8212[14]), .I1(GND_net), .CO(n37864));
    SB_CARRY add_3276_6 (.CI(n36886), .I0(n13113[3]), .I1(n510), .CO(n36887));
    SB_LUT4 add_3276_5_lut (.I0(GND_net), .I1(n13113[2]), .I2(n413_c), 
            .I3(n36885), .O(n12579[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_5_lut (.I0(GND_net), .I1(n1800[2]), .I2(n302), 
            .I3(n38256), .O(n1799[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_16_lut (.I0(GND_net), .I1(n8212[13]), .I2(GND_net), 
            .I3(n37862), .O(n8188[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_5 (.CI(n38256), .I0(n1800[2]), .I1(n302), 
            .CO(n38257));
    SB_CARRY add_3092_16 (.CI(n37862), .I0(n8212[13]), .I1(GND_net), .CO(n37863));
    SB_CARRY add_3276_5 (.CI(n36885), .I0(n13113[2]), .I1(n413_c), .CO(n36886));
    SB_LUT4 add_3276_4_lut (.I0(GND_net), .I1(n13113[1]), .I2(n316), .I3(n36884), 
            .O(n12579[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_4_lut (.I0(GND_net), .I1(n1800[1]), .I2(n229), 
            .I3(n38255), .O(n1799[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_15_lut (.I0(GND_net), .I1(n8212[12]), .I2(GND_net), 
            .I3(n37861), .O(n8188[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_4 (.CI(n38255), .I0(n1800[1]), .I1(n229), 
            .CO(n38256));
    SB_CARRY add_3092_15 (.CI(n37861), .I0(n8212[12]), .I1(GND_net), .CO(n37862));
    SB_CARRY add_3276_4 (.CI(n36884), .I0(n13113[1]), .I1(n316), .CO(n36885));
    SB_LUT4 add_3276_3_lut (.I0(GND_net), .I1(n13113[0]), .I2(n219), .I3(n36883), 
            .O(n12579[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_3_lut (.I0(GND_net), .I1(n1800[0]), .I2(n156), 
            .I3(n38254), .O(n1799[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_14_lut (.I0(GND_net), .I1(n8212[11]), .I2(GND_net), 
            .I3(n37860), .O(n8188[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_3 (.CI(n38254), .I0(n1800[0]), .I1(n156), 
            .CO(n38255));
    SB_CARRY add_3092_14 (.CI(n37860), .I0(n8212[11]), .I1(GND_net), .CO(n37861));
    SB_CARRY add_3276_3 (.CI(n36883), .I0(n13113[0]), .I1(n219), .CO(n36884));
    SB_LUT4 add_3276_2_lut (.I0(GND_net), .I1(n29_c), .I2(n122), .I3(GND_net), 
            .O(n12579[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i209_2_lut (.I0(\Kd[3] ), .I1(n67[6]), .I2(GND_net), 
            .I3(GND_net), .O(n310));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_2_lut (.I0(GND_net), .I1(n14), .I2(n83), 
            .I3(GND_net), .O(n1799[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_13_lut (.I0(GND_net), .I1(n8212[10]), .I2(GND_net), 
            .I3(n37859), .O(n8188[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n38254));
    SB_CARRY add_3092_13 (.CI(n37859), .I0(n8212[10]), .I1(GND_net), .CO(n37860));
    SB_CARRY add_3276_2 (.CI(GND_net), .I0(n29_c), .I1(n122), .CO(n36883));
    SB_LUT4 add_3482_12_lut (.I0(GND_net), .I1(n16424[9]), .I2(GND_net), 
            .I3(n36882), .O(n16318[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_24_lut (.I0(GND_net), .I1(n1799[21]), .I2(GND_net), 
            .I3(n38252), .O(n1798[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_12_lut (.I0(GND_net), .I1(n8212[9]), .I2(GND_net), 
            .I3(n37858), .O(n8188[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_24 (.CI(n38252), .I0(n1799[21]), .I1(GND_net), 
            .CO(n1691));
    SB_CARRY add_3092_12 (.CI(n37858), .I0(n8212[9]), .I1(GND_net), .CO(n37859));
    SB_LUT4 add_3482_11_lut (.I0(GND_net), .I1(n16424[8]), .I2(GND_net), 
            .I3(n36881), .O(n16318[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_11 (.CI(n36881), .I0(n16424[8]), .I1(GND_net), .CO(n36882));
    SB_LUT4 mult_14_add_1213_23_lut (.I0(GND_net), .I1(n1799[20]), .I2(GND_net), 
            .I3(n38251), .O(n1798[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_11_lut (.I0(GND_net), .I1(n8212[8]), .I2(GND_net), 
            .I3(n37857), .O(n8188[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_23 (.CI(n38251), .I0(n1799[20]), .I1(GND_net), 
            .CO(n38252));
    SB_CARRY add_3092_11 (.CI(n37857), .I0(n8212[8]), .I1(GND_net), .CO(n37858));
    SB_LUT4 add_3482_10_lut (.I0(GND_net), .I1(n16424[7]), .I2(GND_net), 
            .I3(n36880), .O(n16318[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_10 (.CI(n36880), .I0(n16424[7]), .I1(GND_net), .CO(n36881));
    SB_LUT4 mult_14_add_1213_22_lut (.I0(GND_net), .I1(n1799[19]), .I2(GND_net), 
            .I3(n38250), .O(n1798[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i4_1_lut (.I0(\deadband[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[3]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3092_10_lut (.I0(GND_net), .I1(n8212[7]), .I2(GND_net), 
            .I3(n37856), .O(n8188[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i274_2_lut (.I0(\Kd[4] ), .I1(n67[6]), .I2(GND_net), 
            .I3(GND_net), .O(n407));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i274_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1213_22 (.CI(n38250), .I0(n1799[19]), .I1(GND_net), 
            .CO(n38251));
    SB_CARRY add_3092_10 (.CI(n37856), .I0(n8212[7]), .I1(GND_net), .CO(n37857));
    SB_LUT4 add_3482_9_lut (.I0(GND_net), .I1(n16424[6]), .I2(GND_net), 
            .I3(n36879), .O(n16318[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_9 (.CI(n36879), .I0(n16424[6]), .I1(GND_net), .CO(n36880));
    SB_LUT4 mult_14_add_1213_21_lut (.I0(GND_net), .I1(n1799[18]), .I2(GND_net), 
            .I3(n38249), .O(n1798[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_9_lut (.I0(GND_net), .I1(n8212[6]), .I2(GND_net), 
            .I3(n37855), .O(n8188[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_21 (.CI(n38249), .I0(n1799[18]), .I1(GND_net), 
            .CO(n38250));
    SB_CARRY add_3092_9 (.CI(n37855), .I0(n8212[6]), .I1(GND_net), .CO(n37856));
    SB_LUT4 add_3482_8_lut (.I0(GND_net), .I1(n16424[5]), .I2(n740), .I3(n36878), 
            .O(n16318[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_8 (.CI(n36878), .I0(n16424[5]), .I1(n740), .CO(n36879));
    SB_LUT4 mult_14_add_1213_20_lut (.I0(GND_net), .I1(n1799[17]), .I2(GND_net), 
            .I3(n38248), .O(n1798[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_8_lut (.I0(GND_net), .I1(n8212[5]), .I2(n707), .I3(n37854), 
            .O(n8188[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_20 (.CI(n38248), .I0(n1799[17]), .I1(GND_net), 
            .CO(n38249));
    SB_CARRY add_3092_8 (.CI(n37854), .I0(n8212[5]), .I1(n707), .CO(n37855));
    SB_LUT4 add_3482_7_lut (.I0(GND_net), .I1(n16424[4]), .I2(n643), .I3(n36877), 
            .O(n16318[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_7 (.CI(n36877), .I0(n16424[4]), .I1(n643), .CO(n36878));
    SB_LUT4 mult_14_add_1213_19_lut (.I0(GND_net), .I1(n1799[16]), .I2(GND_net), 
            .I3(n38247), .O(n1798[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_7_lut (.I0(GND_net), .I1(n8212[4]), .I2(n610), .I3(n37853), 
            .O(n8188[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_19 (.CI(n38247), .I0(n1799[16]), .I1(GND_net), 
            .CO(n38248));
    SB_CARRY add_3092_7 (.CI(n37853), .I0(n8212[4]), .I1(n610), .CO(n37854));
    SB_LUT4 add_3482_6_lut (.I0(GND_net), .I1(n16424[3]), .I2(n546), .I3(n36876), 
            .O(n16318[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_6 (.CI(n36876), .I0(n16424[3]), .I1(n546), .CO(n36877));
    SB_LUT4 mult_14_add_1213_18_lut (.I0(GND_net), .I1(n1799[15]), .I2(GND_net), 
            .I3(n38246), .O(n1798[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_6_lut (.I0(GND_net), .I1(n8212[3]), .I2(n513), .I3(n37852), 
            .O(n8188[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_18 (.CI(n38246), .I0(n1799[15]), .I1(GND_net), 
            .CO(n38247));
    SB_CARRY add_3092_6 (.CI(n37852), .I0(n8212[3]), .I1(n513), .CO(n37853));
    SB_LUT4 add_3482_5_lut (.I0(GND_net), .I1(n16424[2]), .I2(n449_adj_3374), 
            .I3(n36875), .O(n16318[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_5 (.CI(n36875), .I0(n16424[2]), .I1(n449_adj_3374), 
            .CO(n36876));
    SB_LUT4 mult_14_add_1213_17_lut (.I0(GND_net), .I1(n1799[14]), .I2(GND_net), 
            .I3(n38245), .O(n1798[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_5_lut (.I0(GND_net), .I1(n8212[2]), .I2(n416_c), 
            .I3(n37851), .O(n8188[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_17 (.CI(n38245), .I0(n1799[14]), .I1(GND_net), 
            .CO(n38246));
    SB_CARRY add_3092_5 (.CI(n37851), .I0(n8212[2]), .I1(n416_c), .CO(n37852));
    SB_LUT4 add_3482_4_lut (.I0(GND_net), .I1(n16424[1]), .I2(n352), .I3(n36874), 
            .O(n16318[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_4 (.CI(n36874), .I0(n16424[1]), .I1(n352), .CO(n36875));
    SB_LUT4 mult_14_add_1213_16_lut (.I0(GND_net), .I1(n1799[13]), .I2(GND_net), 
            .I3(n38244), .O(n1798[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_4_lut (.I0(GND_net), .I1(n8212[1]), .I2(n319), .I3(n37850), 
            .O(n8188[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_16 (.CI(n38244), .I0(n1799[13]), .I1(GND_net), 
            .CO(n38245));
    SB_CARRY add_3092_4 (.CI(n37850), .I0(n8212[1]), .I1(n319), .CO(n37851));
    SB_LUT4 add_3482_3_lut (.I0(GND_net), .I1(n16424[0]), .I2(n255), .I3(n36873), 
            .O(n16318[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_3 (.CI(n36873), .I0(n16424[0]), .I1(n255), .CO(n36874));
    SB_LUT4 mult_14_add_1213_15_lut (.I0(GND_net), .I1(n1799[12]), .I2(GND_net), 
            .I3(n38243), .O(n1798[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_3_lut (.I0(GND_net), .I1(n8212[0]), .I2(n222), .I3(n37849), 
            .O(n8188[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_15 (.CI(n38243), .I0(n1799[12]), .I1(GND_net), 
            .CO(n38244));
    SB_CARRY add_3092_3 (.CI(n37849), .I0(n8212[0]), .I1(n222), .CO(n37850));
    SB_LUT4 add_3482_2_lut (.I0(GND_net), .I1(n65), .I2(n158), .I3(GND_net), 
            .O(n16318[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_2 (.CI(GND_net), .I0(n65), .I1(n158), .CO(n36873));
    SB_LUT4 mult_14_add_1213_14_lut (.I0(GND_net), .I1(n1799[11]), .I2(GND_net), 
            .I3(n38242), .O(n1798[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_2_lut (.I0(GND_net), .I1(n32_adj_3375), .I2(n125), 
            .I3(GND_net), .O(n8188[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_14 (.CI(n38242), .I0(n1799[11]), .I1(GND_net), 
            .CO(n38243));
    SB_CARRY add_3092_2 (.CI(GND_net), .I0(n32_adj_3375), .I1(n125), .CO(n37849));
    SB_LUT4 add_3300_23_lut (.I0(GND_net), .I1(n13598[20]), .I2(GND_net), 
            .I3(n36872), .O(n13113[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3300_22_lut (.I0(GND_net), .I1(n13598[19]), .I2(GND_net), 
            .I3(n36871), .O(n13113[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_13_lut (.I0(GND_net), .I1(n1799[10]), .I2(GND_net), 
            .I3(n38241), .O(n1798[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_24_lut (.I0(GND_net), .I1(n8188[21]), .I2(GND_net), 
            .I3(n37848), .O(n8163[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_13 (.CI(n38241), .I0(n1799[10]), .I1(GND_net), 
            .CO(n38242));
    SB_LUT4 add_3091_23_lut (.I0(GND_net), .I1(n8188[20]), .I2(GND_net), 
            .I3(n37847), .O(n8163[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_22 (.CI(n36871), .I0(n13598[19]), .I1(GND_net), 
            .CO(n36872));
    SB_LUT4 add_3300_21_lut (.I0(GND_net), .I1(n13598[18]), .I2(GND_net), 
            .I3(n36870), .O(n13113[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i339_2_lut (.I0(\Kd[5] ), .I1(n67[6]), .I2(GND_net), 
            .I3(GND_net), .O(n504));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i339_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1213_12_lut (.I0(GND_net), .I1(n1799[9]), .I2(GND_net), 
            .I3(n38240), .O(n1798[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_23 (.CI(n37847), .I0(n8188[20]), .I1(GND_net), .CO(n37848));
    SB_CARRY mult_14_add_1213_12 (.CI(n38240), .I0(n1799[9]), .I1(GND_net), 
            .CO(n38241));
    SB_LUT4 add_3091_22_lut (.I0(GND_net), .I1(n8188[19]), .I2(GND_net), 
            .I3(n37846), .O(n8163[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_21 (.CI(n36870), .I0(n13598[18]), .I1(GND_net), 
            .CO(n36871));
    SB_LUT4 add_3300_20_lut (.I0(GND_net), .I1(n13598[17]), .I2(GND_net), 
            .I3(n36869), .O(n13113[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_11_lut (.I0(GND_net), .I1(n1799[8]), .I2(GND_net), 
            .I3(n38239), .O(n1798[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_22 (.CI(n37846), .I0(n8188[19]), .I1(GND_net), .CO(n37847));
    SB_CARRY mult_14_add_1213_11 (.CI(n38239), .I0(n1799[8]), .I1(GND_net), 
            .CO(n38240));
    SB_LUT4 add_3091_21_lut (.I0(GND_net), .I1(n8188[18]), .I2(GND_net), 
            .I3(n37845), .O(n8163[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_20 (.CI(n36869), .I0(n13598[17]), .I1(GND_net), 
            .CO(n36870));
    SB_LUT4 add_3300_19_lut (.I0(GND_net), .I1(n13598[16]), .I2(GND_net), 
            .I3(n36868), .O(n13113[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[19]), .I3(n36560), .O(n39_adj_3376)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1213_10_lut (.I0(GND_net), .I1(n1799[7]), .I2(GND_net), 
            .I3(n38238), .O(n1798[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_21 (.CI(n37845), .I0(n8188[18]), .I1(GND_net), .CO(n37846));
    SB_CARRY mult_14_add_1213_10 (.CI(n38238), .I0(n1799[7]), .I1(GND_net), 
            .CO(n38239));
    SB_LUT4 add_3091_20_lut (.I0(GND_net), .I1(n8188[17]), .I2(GND_net), 
            .I3(n37844), .O(n8163[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_19 (.CI(n36868), .I0(n13598[16]), .I1(GND_net), 
            .CO(n36869));
    SB_LUT4 add_3300_18_lut (.I0(GND_net), .I1(n13598[15]), .I2(GND_net), 
            .I3(n36867), .O(n13113[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n36560), .I0(GND_net), .I1(n64[19]), 
            .CO(n36561));
    SB_LUT4 mult_14_add_1213_9_lut (.I0(GND_net), .I1(n1799[6]), .I2(GND_net), 
            .I3(n38237), .O(n1798[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_20 (.CI(n37844), .I0(n8188[17]), .I1(GND_net), .CO(n37845));
    SB_CARRY mult_14_add_1213_9 (.CI(n38237), .I0(n1799[6]), .I1(GND_net), 
            .CO(n38238));
    SB_LUT4 add_3091_19_lut (.I0(GND_net), .I1(n8188[16]), .I2(GND_net), 
            .I3(n37843), .O(n8163[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_18 (.CI(n36867), .I0(n13598[15]), .I1(GND_net), 
            .CO(n36868));
    SB_LUT4 add_3300_17_lut (.I0(GND_net), .I1(n13598[14]), .I2(GND_net), 
            .I3(n36866), .O(n13113[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_8_lut (.I0(GND_net), .I1(n1799[5]), .I2(n518), 
            .I3(n38236), .O(n1798[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_19 (.CI(n37843), .I0(n8188[16]), .I1(GND_net), .CO(n37844));
    SB_CARRY mult_14_add_1213_8 (.CI(n38236), .I0(n1799[5]), .I1(n518), 
            .CO(n38237));
    SB_LUT4 add_3091_18_lut (.I0(GND_net), .I1(n8188[15]), .I2(GND_net), 
            .I3(n37842), .O(n8163[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_17 (.CI(n36866), .I0(n13598[14]), .I1(GND_net), 
            .CO(n36867));
    SB_LUT4 add_3300_16_lut (.I0(GND_net), .I1(n13598[13]), .I2(GND_net), 
            .I3(n36865), .O(n13113[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_7_lut (.I0(GND_net), .I1(n1799[4]), .I2(n445), 
            .I3(n38235), .O(n1798[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_18 (.CI(n37842), .I0(n8188[15]), .I1(GND_net), .CO(n37843));
    SB_CARRY mult_14_add_1213_7 (.CI(n38235), .I0(n1799[4]), .I1(n445), 
            .CO(n38236));
    SB_LUT4 add_3091_17_lut (.I0(GND_net), .I1(n8188[14]), .I2(GND_net), 
            .I3(n37841), .O(n8163[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_16 (.CI(n36865), .I0(n13598[13]), .I1(GND_net), 
            .CO(n36866));
    SB_LUT4 add_3300_15_lut (.I0(GND_net), .I1(n13598[12]), .I2(GND_net), 
            .I3(n36864), .O(n13113[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[18]), .I3(n36559), .O(n37_adj_3378)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1213_6_lut (.I0(GND_net), .I1(n1799[3]), .I2(n372), 
            .I3(n38234), .O(n1798[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_17 (.CI(n37841), .I0(n8188[14]), .I1(GND_net), .CO(n37842));
    SB_CARRY mult_14_add_1213_6 (.CI(n38234), .I0(n1799[3]), .I1(n372), 
            .CO(n38235));
    SB_LUT4 add_3091_16_lut (.I0(GND_net), .I1(n8188[13]), .I2(GND_net), 
            .I3(n37840), .O(n8163[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_15 (.CI(n36864), .I0(n13598[12]), .I1(GND_net), 
            .CO(n36865));
    SB_LUT4 add_3300_14_lut (.I0(GND_net), .I1(n13598[11]), .I2(GND_net), 
            .I3(n36863), .O(n13113[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n36559), .I0(GND_net), .I1(n64[18]), 
            .CO(n36560));
    SB_LUT4 mult_12_i404_2_lut (.I0(\Kd[6] ), .I1(n67[6]), .I2(GND_net), 
            .I3(GND_net), .O(n601_adj_3380));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1213_5_lut (.I0(GND_net), .I1(n1799[2]), .I2(n299), 
            .I3(n38233), .O(n1798[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_16 (.CI(n37840), .I0(n8188[13]), .I1(GND_net), .CO(n37841));
    SB_CARRY mult_14_add_1213_5 (.CI(n38233), .I0(n1799[2]), .I1(n299), 
            .CO(n38234));
    SB_LUT4 add_3091_15_lut (.I0(GND_net), .I1(n8188[12]), .I2(GND_net), 
            .I3(n37839), .O(n8163[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_14 (.CI(n36863), .I0(n13598[11]), .I1(GND_net), 
            .CO(n36864));
    SB_LUT4 add_3300_13_lut (.I0(GND_net), .I1(n13598[10]), .I2(GND_net), 
            .I3(n36862), .O(n13113[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_4_lut (.I0(GND_net), .I1(n1799[1]), .I2(n226), 
            .I3(n38232), .O(n1798[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_15 (.CI(n37839), .I0(n8188[12]), .I1(GND_net), .CO(n37840));
    SB_CARRY mult_14_add_1213_4 (.CI(n38232), .I0(n1799[1]), .I1(n226), 
            .CO(n38233));
    SB_LUT4 add_3091_14_lut (.I0(GND_net), .I1(n8188[11]), .I2(GND_net), 
            .I3(n37838), .O(n8163[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_13 (.CI(n36862), .I0(n13598[10]), .I1(GND_net), 
            .CO(n36863));
    SB_LUT4 add_3300_12_lut (.I0(GND_net), .I1(n13598[9]), .I2(GND_net), 
            .I3(n36861), .O(n13113[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_3_lut (.I0(GND_net), .I1(n1799[0]), .I2(n153), 
            .I3(n38231), .O(n1798[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_14 (.CI(n37838), .I0(n8188[11]), .I1(GND_net), .CO(n37839));
    SB_CARRY mult_14_add_1213_3 (.CI(n38231), .I0(n1799[0]), .I1(n153), 
            .CO(n38232));
    SB_LUT4 add_3091_13_lut (.I0(GND_net), .I1(n8188[10]), .I2(GND_net), 
            .I3(n37837), .O(n8163[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_12 (.CI(n36861), .I0(n13598[9]), .I1(GND_net), .CO(n36862));
    SB_LUT4 state_23__I_0_add_2_26_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n70[23]), .I3(n36670), .O(\PID_CONTROLLER.err_31__N_2816 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[17]), .I3(n36558), .O(n35_adj_3382)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3300_11_lut (.I0(GND_net), .I1(n13598[8]), .I2(GND_net), 
            .I3(n36860), .O(n13113[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n36558), .I0(GND_net), .I1(n64[17]), 
            .CO(n36559));
    SB_LUT4 mult_14_add_1213_2_lut (.I0(GND_net), .I1(n11_c), .I2(n80), 
            .I3(GND_net), .O(n1798[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_13 (.CI(n37837), .I0(n8188[10]), .I1(GND_net), .CO(n37838));
    SB_CARRY mult_14_add_1213_2 (.CI(GND_net), .I0(n11_c), .I1(n80), .CO(n38231));
    SB_LUT4 add_3091_12_lut (.I0(GND_net), .I1(n8188[9]), .I2(GND_net), 
            .I3(n37836), .O(n8163[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_11 (.CI(n36860), .I0(n13598[8]), .I1(GND_net), .CO(n36861));
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n70[23]), .I3(n36669), .O(\PID_CONTROLLER.err_31__N_2816 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[16]), .I3(n36557), .O(n33_adj_3383)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3300_10_lut (.I0(GND_net), .I1(n13598[7]), .I2(GND_net), 
            .I3(n36859), .O(n13113[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n36557), .I0(GND_net), .I1(n64[16]), 
            .CO(n36558));
    SB_LUT4 unary_minus_17_inv_0_i5_1_lut (.I0(\deadband[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[4]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_add_1212_24_lut (.I0(GND_net), .I1(n1798[21]), .I2(GND_net), 
            .I3(n38229), .O(n1797[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_12 (.CI(n37836), .I0(n8188[9]), .I1(GND_net), .CO(n37837));
    SB_LUT4 add_3091_11_lut (.I0(GND_net), .I1(n8188[8]), .I2(GND_net), 
            .I3(n37835), .O(n8163[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_24 (.CI(n38229), .I0(n1798[21]), .I1(GND_net), 
            .CO(n1687));
    SB_CARRY add_3091_11 (.CI(n37835), .I0(n8188[8]), .I1(GND_net), .CO(n37836));
    SB_LUT4 mult_12_i469_2_lut (.I0(\Kd[7] ), .I1(n67[6]), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1212_23_lut (.I0(GND_net), .I1(n1798[20]), .I2(GND_net), 
            .I3(n38228), .O(n1797[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_10_lut (.I0(GND_net), .I1(n8188[7]), .I2(GND_net), 
            .I3(n37834), .O(n8163[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_10 (.CI(n36859), .I0(n13598[7]), .I1(GND_net), .CO(n36860));
    SB_LUT4 add_3300_9_lut (.I0(GND_net), .I1(n13598[6]), .I2(GND_net), 
            .I3(n36858), .O(n13113[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_23 (.CI(n38228), .I0(n1798[20]), .I1(GND_net), 
            .CO(n38229));
    SB_CARRY add_3091_10 (.CI(n37834), .I0(n8188[7]), .I1(GND_net), .CO(n37835));
    SB_LUT4 mult_14_add_1212_22_lut (.I0(GND_net), .I1(n1798[19]), .I2(GND_net), 
            .I3(n38227), .O(n1797[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_9_lut (.I0(GND_net), .I1(n8188[6]), .I2(GND_net), 
            .I3(n37833), .O(n8163[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_9 (.CI(n36858), .I0(n13598[6]), .I1(GND_net), .CO(n36859));
    SB_LUT4 add_3300_8_lut (.I0(GND_net), .I1(n13598[5]), .I2(n707_adj_3385), 
            .I3(n36857), .O(n13113[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_22 (.CI(n38227), .I0(n1798[19]), .I1(GND_net), 
            .CO(n38228));
    SB_CARRY add_3091_9 (.CI(n37833), .I0(n8188[6]), .I1(GND_net), .CO(n37834));
    SB_LUT4 mult_14_add_1212_21_lut (.I0(GND_net), .I1(n1798[18]), .I2(GND_net), 
            .I3(n38226), .O(n1797[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_8_lut (.I0(GND_net), .I1(n8188[5]), .I2(n704_adj_3386), 
            .I3(n37832), .O(n8163[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_8 (.CI(n36857), .I0(n13598[5]), .I1(n707_adj_3385), 
            .CO(n36858));
    SB_CARRY state_23__I_0_add_2_25 (.CI(n36669), .I0(\motor_state[23] ), 
            .I1(n70[23]), .CO(n36670));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[15]), .I3(n36556), .O(n31_adj_3387)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3300_7_lut (.I0(GND_net), .I1(n13598[4]), .I2(n610_adj_3388), 
            .I3(n36856), .O(n13113[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n36556), .I0(GND_net), .I1(n64[15]), 
            .CO(n36557));
    SB_CARRY mult_14_add_1212_21 (.CI(n38226), .I0(n1798[18]), .I1(GND_net), 
            .CO(n38227));
    SB_CARRY add_3091_8 (.CI(n37832), .I0(n8188[5]), .I1(n704_adj_3386), 
            .CO(n37833));
    SB_LUT4 mult_14_add_1212_20_lut (.I0(GND_net), .I1(n1798[17]), .I2(GND_net), 
            .I3(n38225), .O(n1797[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_7_lut (.I0(GND_net), .I1(n8188[4]), .I2(n607_adj_3389), 
            .I3(n37831), .O(n8163[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_7 (.CI(n36856), .I0(n13598[4]), .I1(n610_adj_3388), 
            .CO(n36857));
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(\motor_state[22] ), 
            .I2(n70[22]), .I3(n36668), .O(\PID_CONTROLLER.err_31__N_2816 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[14]), .I3(n36555), .O(n29_adj_3391)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3300_6_lut (.I0(GND_net), .I1(n13598[3]), .I2(n513_adj_3393), 
            .I3(n36855), .O(n13113[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n36555), .I0(GND_net), .I1(n64[14]), 
            .CO(n36556));
    SB_CARRY mult_14_add_1212_20 (.CI(n38225), .I0(n1798[17]), .I1(GND_net), 
            .CO(n38226));
    SB_CARRY add_3091_7 (.CI(n37831), .I0(n8188[4]), .I1(n607_adj_3389), 
            .CO(n37832));
    SB_LUT4 mult_14_add_1212_19_lut (.I0(GND_net), .I1(n1798[16]), .I2(GND_net), 
            .I3(n38224), .O(n1797[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_6_lut (.I0(GND_net), .I1(n8188[3]), .I2(n510_adj_3394), 
            .I3(n37830), .O(n8163[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_6 (.CI(n36855), .I0(n13598[3]), .I1(n513_adj_3393), 
            .CO(n36856));
    SB_LUT4 add_3300_5_lut (.I0(GND_net), .I1(n13598[2]), .I2(n416_adj_3395), 
            .I3(n36854), .O(n13113[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[0]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_14_add_1212_19 (.CI(n38224), .I0(n1798[16]), .I1(GND_net), 
            .CO(n38225));
    SB_CARRY add_3091_6 (.CI(n37830), .I0(n8188[3]), .I1(n510_adj_3394), 
            .CO(n37831));
    SB_LUT4 mult_14_add_1212_18_lut (.I0(GND_net), .I1(n1798[15]), .I2(GND_net), 
            .I3(n38223), .O(n1797[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_5_lut (.I0(GND_net), .I1(n8188[2]), .I2(n413_adj_3396), 
            .I3(n37829), .O(n8163[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_5 (.CI(n36854), .I0(n13598[2]), .I1(n416_adj_3395), 
            .CO(n36855));
    SB_LUT4 add_3300_4_lut (.I0(GND_net), .I1(n13598[1]), .I2(n319_adj_3397), 
            .I3(n36853), .O(n13113[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_18 (.CI(n38223), .I0(n1798[15]), .I1(GND_net), 
            .CO(n38224));
    SB_CARRY add_3091_5 (.CI(n37829), .I0(n8188[2]), .I1(n413_adj_3396), 
            .CO(n37830));
    SB_LUT4 mult_14_add_1212_17_lut (.I0(GND_net), .I1(n1798[14]), .I2(GND_net), 
            .I3(n38222), .O(n1797[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_4_lut (.I0(GND_net), .I1(n8188[1]), .I2(n316_adj_3398), 
            .I3(n37828), .O(n8163[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_4 (.CI(n36853), .I0(n13598[1]), .I1(n319_adj_3397), 
            .CO(n36854));
    SB_CARRY state_23__I_0_add_2_24 (.CI(n36668), .I0(\motor_state[22] ), 
            .I1(n70[22]), .CO(n36669));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[13]), .I3(n36554), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3300_3_lut (.I0(GND_net), .I1(n13598[0]), .I2(n222_adj_3399), 
            .I3(n36852), .O(n13113[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n36554), .I0(GND_net), .I1(n64[13]), 
            .CO(n36555));
    SB_CARRY mult_14_add_1212_17 (.CI(n38222), .I0(n1798[14]), .I1(GND_net), 
            .CO(n38223));
    SB_CARRY add_3091_4 (.CI(n37828), .I0(n8188[1]), .I1(n316_adj_3398), 
            .CO(n37829));
    SB_LUT4 mult_14_add_1212_16_lut (.I0(GND_net), .I1(n1798[13]), .I2(GND_net), 
            .I3(n38221), .O(n1797[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_3_lut (.I0(GND_net), .I1(n8188[0]), .I2(n219_adj_3400), 
            .I3(n37827), .O(n8163[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_3 (.CI(n36852), .I0(n13598[0]), .I1(n222_adj_3399), 
            .CO(n36853));
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(\motor_state[21] ), 
            .I2(n70[21]), .I3(n36667), .O(\PID_CONTROLLER.err_31__N_2816 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[12]), .I3(n36553), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3300_2_lut (.I0(GND_net), .I1(n32_adj_3402), .I2(n125_adj_3403), 
            .I3(GND_net), .O(n13113[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n36667), .I0(\motor_state[21] ), 
            .I1(n70[21]), .CO(n36668));
    SB_CARRY unary_minus_5_add_3_14 (.CI(n36553), .I0(GND_net), .I1(n64[12]), 
            .CO(n36554));
    SB_CARRY mult_14_add_1212_16 (.CI(n38221), .I0(n1798[13]), .I1(GND_net), 
            .CO(n38222));
    SB_CARRY add_3091_3 (.CI(n37827), .I0(n8188[0]), .I1(n219_adj_3400), 
            .CO(n37828));
    SB_LUT4 mult_14_add_1212_15_lut (.I0(GND_net), .I1(n1798[12]), .I2(GND_net), 
            .I3(n38220), .O(n1797[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_2_lut (.I0(GND_net), .I1(n29_adj_3404), .I2(n122_adj_3405), 
            .I3(GND_net), .O(n8163[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_15 (.CI(n38220), .I0(n1798[12]), .I1(GND_net), 
            .CO(n38221));
    SB_CARRY add_3091_2 (.CI(GND_net), .I0(n29_adj_3404), .I1(n122_adj_3405), 
            .CO(n37827));
    SB_CARRY add_3300_2 (.CI(GND_net), .I0(n32_adj_3402), .I1(n125_adj_3403), 
            .CO(n36852));
    SB_LUT4 add_3322_22_lut (.I0(GND_net), .I1(n14039[19]), .I2(GND_net), 
            .I3(n36851), .O(n13598[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_14_lut (.I0(GND_net), .I1(n1798[11]), .I2(GND_net), 
            .I3(n38219), .O(n1797[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_25_lut (.I0(GND_net), .I1(n8163[22]), .I2(GND_net), 
            .I3(n37826), .O(n8137[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_14 (.CI(n38219), .I0(n1798[11]), .I1(GND_net), 
            .CO(n38220));
    SB_LUT4 add_3090_24_lut (.I0(GND_net), .I1(n8163[21]), .I2(GND_net), 
            .I3(n37825), .O(n8137[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_21_lut (.I0(GND_net), .I1(n14039[18]), .I2(GND_net), 
            .I3(n36850), .O(n13598[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_21 (.CI(n36850), .I0(n14039[18]), .I1(GND_net), 
            .CO(n36851));
    SB_LUT4 mult_14_add_1212_13_lut (.I0(GND_net), .I1(n1798[10]), .I2(GND_net), 
            .I3(n38218), .O(n1797[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_24 (.CI(n37825), .I0(n8163[21]), .I1(GND_net), .CO(n37826));
    SB_CARRY mult_14_add_1212_13 (.CI(n38218), .I0(n1798[10]), .I1(GND_net), 
            .CO(n38219));
    SB_LUT4 add_3090_23_lut (.I0(GND_net), .I1(n8163[20]), .I2(GND_net), 
            .I3(n37824), .O(n8137[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_20_lut (.I0(GND_net), .I1(n14039[17]), .I2(GND_net), 
            .I3(n36849), .O(n13598[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(\motor_state[20] ), 
            .I2(n70[20]), .I3(n36666), .O(\PID_CONTROLLER.err_31__N_2816 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[11]), .I3(n36552), .O(n23_adj_3407)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3322_20 (.CI(n36849), .I0(n14039[17]), .I1(GND_net), 
            .CO(n36850));
    SB_CARRY unary_minus_5_add_3_13 (.CI(n36552), .I0(GND_net), .I1(n64[11]), 
            .CO(n36553));
    SB_LUT4 mult_14_add_1212_12_lut (.I0(GND_net), .I1(n1798[9]), .I2(GND_net), 
            .I3(n38217), .O(n1797[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_23 (.CI(n37824), .I0(n8163[20]), .I1(GND_net), .CO(n37825));
    SB_CARRY mult_14_add_1212_12 (.CI(n38217), .I0(n1798[9]), .I1(GND_net), 
            .CO(n38218));
    SB_LUT4 add_3090_22_lut (.I0(GND_net), .I1(n8163[19]), .I2(GND_net), 
            .I3(n37823), .O(n8137[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_19_lut (.I0(GND_net), .I1(n14039[16]), .I2(GND_net), 
            .I3(n36848), .O(n13598[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n36666), .I0(\motor_state[20] ), 
            .I1(n70[20]), .CO(n36667));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[10]), .I3(n36551), .O(n21_c)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3322_19 (.CI(n36848), .I0(n14039[16]), .I1(GND_net), 
            .CO(n36849));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n36551), .I0(GND_net), .I1(n64[10]), 
            .CO(n36552));
    SB_LUT4 mult_10_i113_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n167));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i50_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_3409));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i50_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1212_11_lut (.I0(GND_net), .I1(n1798[8]), .I2(GND_net), 
            .I3(n38216), .O(n1797[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_22 (.CI(n37823), .I0(n8163[19]), .I1(GND_net), .CO(n37824));
    SB_CARRY mult_14_add_1212_11 (.CI(n38216), .I0(n1798[8]), .I1(GND_net), 
            .CO(n38217));
    SB_LUT4 add_3090_21_lut (.I0(GND_net), .I1(n8163[18]), .I2(GND_net), 
            .I3(n37822), .O(n8137[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_18_lut (.I0(GND_net), .I1(n14039[15]), .I2(GND_net), 
            .I3(n36847), .O(n13598[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_18 (.CI(n36847), .I0(n14039[15]), .I1(GND_net), 
            .CO(n36848));
    SB_LUT4 mult_10_i178_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n264));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1212_10_lut (.I0(GND_net), .I1(n1798[7]), .I2(GND_net), 
            .I3(n38215), .O(n1797[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_21 (.CI(n37822), .I0(n8163[18]), .I1(GND_net), .CO(n37823));
    SB_CARRY mult_14_add_1212_10 (.CI(n38215), .I0(n1798[7]), .I1(GND_net), 
            .CO(n38216));
    SB_LUT4 add_3090_20_lut (.I0(GND_net), .I1(n8163[17]), .I2(GND_net), 
            .I3(n37821), .O(n8137[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_17_lut (.I0(GND_net), .I1(n14039[14]), .I2(GND_net), 
            .I3(n36846), .O(n13598[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_17 (.CI(n36846), .I0(n14039[14]), .I1(GND_net), 
            .CO(n36847));
    SB_LUT4 mult_14_add_1212_9_lut (.I0(GND_net), .I1(n1798[6]), .I2(GND_net), 
            .I3(n38214), .O(n1797[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_20 (.CI(n37821), .I0(n8163[17]), .I1(GND_net), .CO(n37822));
    SB_LUT4 add_3322_16_lut (.I0(GND_net), .I1(n14039[13]), .I2(GND_net), 
            .I3(n36845), .O(n13598[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n64[9]), .I3(n36550), .O(n19_c)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_14_add_1212_9 (.CI(n38214), .I0(n1798[6]), .I1(GND_net), 
            .CO(n38215));
    SB_LUT4 add_3090_19_lut (.I0(GND_net), .I1(n8163[16]), .I2(GND_net), 
            .I3(n37820), .O(n8137[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_16 (.CI(n36845), .I0(n14039[13]), .I1(GND_net), 
            .CO(n36846));
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(\motor_state[19] ), 
            .I2(n70[19]), .I3(n36665), .O(\PID_CONTROLLER.err_31__N_2816 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n36550), .I0(GND_net), .I1(n64[9]), 
            .CO(n36551));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n64[8]), .I3(n36549), .O(n17_adj_3411)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1212_8_lut (.I0(GND_net), .I1(n1798[5]), .I2(n515), 
            .I3(n38213), .O(n1797[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_19 (.CI(n37820), .I0(n8163[16]), .I1(GND_net), .CO(n37821));
    SB_LUT4 add_3322_15_lut (.I0(GND_net), .I1(n14039[12]), .I2(GND_net), 
            .I3(n36844), .O(n13598[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n36549), .I0(GND_net), .I1(n64[8]), 
            .CO(n36550));
    SB_CARRY mult_14_add_1212_8 (.CI(n38213), .I0(n1798[5]), .I1(n515), 
            .CO(n38214));
    SB_LUT4 add_3090_18_lut (.I0(GND_net), .I1(n8163[15]), .I2(GND_net), 
            .I3(n37819), .O(n8137[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_15 (.CI(n36844), .I0(n14039[12]), .I1(GND_net), 
            .CO(n36845));
    SB_CARRY state_23__I_0_add_2_21 (.CI(n36665), .I0(\motor_state[19] ), 
            .I1(n70[19]), .CO(n36666));
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n64[7]), .I3(n36548), .O(n15_adj_3414)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n36548), .I0(GND_net), .I1(n64[7]), 
            .CO(n36549));
    SB_LUT4 mult_14_add_1212_7_lut (.I0(GND_net), .I1(n1798[4]), .I2(n442), 
            .I3(n38212), .O(n1797[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_18 (.CI(n37819), .I0(n8163[15]), .I1(GND_net), .CO(n37820));
    SB_CARRY mult_14_add_1212_7 (.CI(n38212), .I0(n1798[4]), .I1(n442), 
            .CO(n38213));
    SB_LUT4 add_3090_17_lut (.I0(GND_net), .I1(n8163[14]), .I2(GND_net), 
            .I3(n37818), .O(n8137[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_14_lut (.I0(GND_net), .I1(n14039[11]), .I2(GND_net), 
            .I3(n36843), .O(n13598[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_14 (.CI(n36843), .I0(n14039[11]), .I1(GND_net), 
            .CO(n36844));
    SB_LUT4 mult_10_i243_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n361));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1212_6_lut (.I0(GND_net), .I1(n1798[3]), .I2(n369), 
            .I3(n38211), .O(n1797[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_17 (.CI(n37818), .I0(n8163[14]), .I1(GND_net), .CO(n37819));
    SB_CARRY mult_14_add_1212_6 (.CI(n38211), .I0(n1798[3]), .I1(n369), 
            .CO(n38212));
    SB_LUT4 add_3090_16_lut (.I0(GND_net), .I1(n8163[13]), .I2(GND_net), 
            .I3(n37817), .O(n8137[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_13_lut (.I0(GND_net), .I1(n14039[10]), .I2(GND_net), 
            .I3(n36842), .O(n13598[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_13 (.CI(n36842), .I0(n14039[10]), .I1(GND_net), 
            .CO(n36843));
    SB_LUT4 mult_14_add_1212_5_lut (.I0(GND_net), .I1(n1798[2]), .I2(n296), 
            .I3(n38210), .O(n1797[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_16 (.CI(n37817), .I0(n8163[13]), .I1(GND_net), .CO(n37818));
    SB_LUT4 add_3322_12_lut (.I0(GND_net), .I1(n14039[9]), .I2(GND_net), 
            .I3(n36841), .O(n13598[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n64[6]), .I3(n36547), .O(n13_adj_3415)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_14_add_1212_5 (.CI(n38210), .I0(n1798[2]), .I1(n296), 
            .CO(n38211));
    SB_LUT4 add_3090_15_lut (.I0(GND_net), .I1(n8163[12]), .I2(GND_net), 
            .I3(n37816), .O(n8137[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n458_c));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3322_12 (.CI(n36841), .I0(n14039[9]), .I1(GND_net), .CO(n36842));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(\motor_state[18] ), 
            .I2(n70[18]), .I3(n36664), .O(\PID_CONTROLLER.err_31__N_2816 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n36547), .I0(GND_net), .I1(n64[6]), 
            .CO(n36548));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n64[5]), .I3(n36546), .O(n11_adj_3418)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1212_4_lut (.I0(GND_net), .I1(n1798[1]), .I2(n223), 
            .I3(n38209), .O(n1797[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_15 (.CI(n37816), .I0(n8163[12]), .I1(GND_net), .CO(n37817));
    SB_LUT4 add_3322_11_lut (.I0(GND_net), .I1(n14039[8]), .I2(GND_net), 
            .I3(n36840), .O(n13598[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n36546), .I0(GND_net), .I1(n64[5]), 
            .CO(n36547));
    SB_CARRY mult_14_add_1212_4 (.CI(n38209), .I0(n1798[1]), .I1(n223), 
            .CO(n38210));
    SB_LUT4 add_3090_14_lut (.I0(GND_net), .I1(n8163[11]), .I2(GND_net), 
            .I3(n37815), .O(n8137[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_11 (.CI(n36840), .I0(n14039[8]), .I1(GND_net), .CO(n36841));
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n555));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_DFF pwm__i0 (.Q(pwm[0]), .C(clk32MHz), .D(n24454));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i23 (.Q(pwm[23]), .C(clk32MHz), .D(n24451));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i22 (.Q(pwm[22]), .C(clk32MHz), .D(n24450));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i21 (.Q(pwm[21]), .C(clk32MHz), .D(n24449));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i20 (.Q(pwm[20]), .C(clk32MHz), .D(n24448));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i19 (.Q(pwm[19]), .C(clk32MHz), .D(n24447));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i18 (.Q(pwm[18]), .C(clk32MHz), .D(n41482));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i17 (.Q(pwm[17]), .C(clk32MHz), .D(n41480));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i16 (.Q(pwm[16]), .C(clk32MHz), .D(n24444));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i15 (.Q(pwm[15]), .C(clk32MHz), .D(n24443));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i14 (.Q(pwm[14]), .C(clk32MHz), .D(n24442));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i13 (.Q(pwm[13]), .C(clk32MHz), .D(n24441));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i12 (.Q(pwm[12]), .C(clk32MHz), .D(n24440));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i11 (.Q(pwm[11]), .C(clk32MHz), .D(n24439));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i10 (.Q(pwm[10]), .C(clk32MHz), .D(n24438));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i9 (.Q(pwm[9]), .C(clk32MHz), .D(n24437));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i8 (.Q(pwm[8]), .C(clk32MHz), .D(n24436));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i7 (.Q(pwm[7]), .C(clk32MHz), .D(n24435));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i6 (.Q(pwm[6]), .C(clk32MHz), .D(n24434));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i5 (.Q(pwm[5]), .C(clk32MHz), .D(n24433));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i4 (.Q(pwm[4]), .C(clk32MHz), .D(n24432));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i3 (.Q(pwm[3]), .C(clk32MHz), .D(n24431));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i2 (.Q(pwm[2]), .C(clk32MHz), .D(n24430));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i1 (.Q(pwm[1]), .C(clk32MHz), .D(n24426));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 mult_10_i438_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n652));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i503_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i95_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n140));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i160_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n237));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i225_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n334));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i290_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n431));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i290_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n36664), .I0(\motor_state[18] ), 
            .I1(n70[18]), .CO(n36665));
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n528_adj_3419));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n625));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i485_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n722));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n64[4]), .I3(n36545), .O(n9_adj_3420)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1212_3_lut (.I0(GND_net), .I1(n1798[0]), .I2(n150), 
            .I3(n38208), .O(n1797[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i6_1_lut (.I0(\deadband[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[5]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i109_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i46_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n68));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i46_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3090_14 (.CI(n37815), .I0(n8163[11]), .I1(GND_net), .CO(n37816));
    SB_CARRY mult_14_add_1212_3 (.CI(n38208), .I0(n1798[0]), .I1(n150), 
            .CO(n38209));
    SB_LUT4 add_3090_13_lut (.I0(GND_net), .I1(n8163[10]), .I2(GND_net), 
            .I3(n37814), .O(n8137[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_13 (.CI(n37814), .I0(n8163[10]), .I1(GND_net), .CO(n37815));
    SB_LUT4 mult_14_add_1212_2_lut (.I0(GND_net), .I1(n8_adj_3422), .I2(n77), 
            .I3(GND_net), .O(n1797[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_12_lut (.I0(GND_net), .I1(n8163[9]), .I2(GND_net), 
            .I3(n37813), .O(n8137[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_12 (.CI(n37813), .I0(n8163[9]), .I1(GND_net), .CO(n37814));
    SB_LUT4 add_3090_11_lut (.I0(GND_net), .I1(n8163[8]), .I2(GND_net), 
            .I3(n37812), .O(n8137[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_11 (.CI(n37812), .I0(n8163[8]), .I1(GND_net), .CO(n37813));
    SB_LUT4 add_3090_10_lut (.I0(GND_net), .I1(n8163[7]), .I2(GND_net), 
            .I3(n37811), .O(n8137[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_10 (.CI(n37811), .I0(n8163[7]), .I1(GND_net), .CO(n37812));
    SB_CARRY mult_14_add_1212_2 (.CI(GND_net), .I0(n8_adj_3422), .I1(n77), 
            .CO(n38208));
    SB_LUT4 add_3090_9_lut (.I0(GND_net), .I1(n8163[6]), .I2(GND_net), 
            .I3(n37810), .O(n8137[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_10_lut (.I0(GND_net), .I1(n14039[7]), .I2(GND_net), 
            .I3(n36839), .O(n13598[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_10 (.CI(n36839), .I0(n14039[7]), .I1(GND_net), .CO(n36840));
    SB_LUT4 mult_14_add_1211_24_lut (.I0(GND_net), .I1(n1797[21]), .I2(GND_net), 
            .I3(n38206), .O(n1796[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_9 (.CI(n37810), .I0(n8163[6]), .I1(GND_net), .CO(n37811));
    SB_LUT4 add_3322_9_lut (.I0(GND_net), .I1(n14039[6]), .I2(GND_net), 
            .I3(n36838), .O(n13598[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(\motor_state[17] ), 
            .I2(n70[17]), .I3(n36663), .O(\PID_CONTROLLER.err_31__N_2816 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_9 (.CI(n36838), .I0(n14039[6]), .I1(GND_net), .CO(n36839));
    SB_CARRY state_23__I_0_add_2_19 (.CI(n36663), .I0(\motor_state[17] ), 
            .I1(n70[17]), .CO(n36664));
    SB_CARRY mult_14_add_1211_24 (.CI(n38206), .I0(n1797[21]), .I1(GND_net), 
            .CO(n1683));
    SB_LUT4 add_3090_8_lut (.I0(GND_net), .I1(n8163[5]), .I2(n701), .I3(n37809), 
            .O(n8137[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_8_lut (.I0(GND_net), .I1(n14039[5]), .I2(n710_adj_3424), 
            .I3(n36837), .O(n13598[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(\motor_state[16] ), 
            .I2(n70[16]), .I3(n36662), .O(\PID_CONTROLLER.err_31__N_2816 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_8 (.CI(n36837), .I0(n14039[5]), .I1(n710_adj_3424), 
            .CO(n36838));
    SB_CARRY state_23__I_0_add_2_18 (.CI(n36662), .I0(\motor_state[16] ), 
            .I1(n70[16]), .CO(n36663));
    SB_LUT4 mult_14_add_1211_23_lut (.I0(GND_net), .I1(n1797[20]), .I2(GND_net), 
            .I3(n38205), .O(n282[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_8 (.CI(n37809), .I0(n8163[5]), .I1(n701), .CO(n37810));
    SB_LUT4 add_3322_7_lut (.I0(GND_net), .I1(n14039[4]), .I2(n613_adj_3426), 
            .I3(n36836), .O(n13598[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(\motor_state[15] ), 
            .I2(n70[15]), .I3(n36661), .O(\PID_CONTROLLER.err_31__N_2816 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n36545), .I0(GND_net), .I1(n64[4]), 
            .CO(n36546));
    SB_CARRY state_23__I_0_add_2_17 (.CI(n36661), .I0(\motor_state[15] ), 
            .I1(n70[15]), .CO(n36662));
    SB_CARRY add_3322_7 (.CI(n36836), .I0(n14039[4]), .I1(n613_adj_3426), 
            .CO(n36837));
    SB_LUT4 add_3090_7_lut (.I0(GND_net), .I1(n8163[4]), .I2(n604), .I3(n37808), 
            .O(n8137[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_6_lut (.I0(GND_net), .I1(n14039[3]), .I2(n516_adj_3428), 
            .I3(n36835), .O(n13598[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(\motor_state[14] ), 
            .I2(n70[14]), .I3(n36660), .O(\PID_CONTROLLER.err_31__N_2816 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n64[3]), .I3(n36544), .O(n7_adj_3430)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n36660), .I0(\motor_state[14] ), 
            .I1(n70[14]), .CO(n36661));
    SB_CARRY mult_14_add_1211_23 (.CI(n38205), .I0(n1797[20]), .I1(GND_net), 
            .CO(n38206));
    SB_CARRY add_3090_7 (.CI(n37808), .I0(n8163[4]), .I1(n604), .CO(n37809));
    SB_CARRY add_3322_6 (.CI(n36835), .I0(n14039[3]), .I1(n516_adj_3428), 
            .CO(n36836));
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(\motor_state[13] ), 
            .I2(n70[13]), .I3(n36659), .O(\PID_CONTROLLER.err_31__N_2816 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.result_i0  (.Q(\PID_CONTROLLER.result [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [0]));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 mult_14_add_1211_22_lut (.I0(GND_net), .I1(n1797[19]), .I2(GND_net), 
            .I3(n38204), .O(n282[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n36659), .I0(\motor_state[13] ), 
            .I1(n70[13]), .CO(n36660));
    SB_LUT4 mult_14_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3090_6_lut (.I0(GND_net), .I1(n8163[3]), .I2(n507), .I3(n37807), 
            .O(n8137[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err[0] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [0]));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3322_5_lut (.I0(GND_net), .I1(n14039[2]), .I2(n419_adj_3432), 
            .I3(n36834), .O(n13598[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_22 (.CI(n38204), .I0(n1797[19]), .I1(GND_net), 
            .CO(n38205));
    SB_CARRY add_3090_6 (.CI(n37807), .I0(n8163[3]), .I1(n507), .CO(n37808));
    SB_CARRY add_3322_5 (.CI(n36834), .I0(n14039[2]), .I1(n419_adj_3432), 
            .CO(n36835));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(\motor_state[12] ), 
            .I2(n70[12]), .I3(n36658), .O(\PID_CONTROLLER.err_31__N_2816 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n36544), .I0(GND_net), .I1(n64[3]), 
            .CO(n36545));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n64[2]), .I3(n36543), .O(n5_adj_3434)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3322_4_lut (.I0(GND_net), .I1(n14039[1]), .I2(n322_adj_3436), 
            .I3(n36833), .O(n13598[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n36658), .I0(\motor_state[12] ), 
            .I1(n70[12]), .CO(n36659));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n36543), .I0(GND_net), .I1(n64[2]), 
            .CO(n36544));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n64[1]), .I3(n36542), .O(n3_adj_3437)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1211_21_lut (.I0(GND_net), .I1(n1797[18]), .I2(GND_net), 
            .I3(n38203), .O(n282[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_21 (.CI(n38203), .I0(n1797[18]), .I1(GND_net), 
            .CO(n38204));
    SB_LUT4 add_3090_5_lut (.I0(GND_net), .I1(n8163[2]), .I2(n410), .I3(n37806), 
            .O(n8137[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3439));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i4_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3322_4 (.CI(n36833), .I0(n14039[1]), .I1(n322_adj_3436), 
            .CO(n36834));
    SB_LUT4 mult_14_add_1211_20_lut (.I0(GND_net), .I1(n1797[17]), .I2(GND_net), 
            .I3(n38202), .O(n282[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(\motor_state[11] ), 
            .I2(n70[11]), .I3(n36657), .O(\PID_CONTROLLER.err_31__N_2816 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_3_lut (.I0(GND_net), .I1(n14039[0]), .I2(n225_adj_3442), 
            .I3(n36832), .O(n13598[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_5 (.CI(n37806), .I0(n8163[2]), .I1(n410), .CO(n37807));
    SB_CARRY state_23__I_0_add_2_13 (.CI(n36657), .I0(\motor_state[11] ), 
            .I1(n70[11]), .CO(n36658));
    SB_CARRY mult_14_add_1211_20 (.CI(n38202), .I0(n1797[17]), .I1(GND_net), 
            .CO(n38203));
    SB_LUT4 add_3090_4_lut (.I0(GND_net), .I1(n8163[1]), .I2(n313), .I3(n37805), 
            .O(n8137[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_19_lut (.I0(GND_net), .I1(n1797[16]), .I2(GND_net), 
            .I3(n38201), .O(n282[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_3 (.CI(n36832), .I0(n14039[0]), .I1(n225_adj_3442), 
            .CO(n36833));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(\motor_state[10] ), 
            .I2(n70[10]), .I3(n36656), .O(\PID_CONTROLLER.err_31__N_2816 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n36542), .I0(GND_net), .I1(n64[1]), 
            .CO(n36543));
    SB_LUT4 mult_14_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n64[0]), 
            .I3(VCC_net), .O(n63[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_2_lut (.I0(GND_net), .I1(n35_adj_3445), .I2(n128_adj_3446), 
            .I3(GND_net), .O(n13598[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_12 (.CI(n36656), .I0(\motor_state[10] ), 
            .I1(n70[10]), .CO(n36657));
    SB_CARRY add_3322_2 (.CI(GND_net), .I0(n35_adj_3445), .I1(n128_adj_3446), 
            .CO(n36832));
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(\motor_state[9] ), 
            .I2(n70[9]), .I3(n36655), .O(\PID_CONTROLLER.err_31__N_2816 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n64[0]), 
            .CO(n36542));
    SB_LUT4 mult_14_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i149_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3090_4 (.CI(n37805), .I0(n8163[1]), .I1(n313), .CO(n37806));
    SB_LUT4 add_3090_3_lut (.I0(GND_net), .I1(n8163[0]), .I2(n216), .I3(n37804), 
            .O(n8137[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_3 (.CI(n37804), .I0(n8163[0]), .I1(n216), .CO(n37805));
    SB_CARRY state_23__I_0_add_2_11 (.CI(n36655), .I0(\motor_state[9] ), 
            .I1(n70[9]), .CO(n36656));
    SB_LUT4 unary_minus_17_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n69[31]), 
            .I3(n36541), .O(pwm_23__N_2951[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(\motor_state[8] ), 
            .I2(n70[8]), .I3(n36654), .O(\PID_CONTROLLER.err_31__N_2816 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n69[31]), 
            .I3(n36540), .O(pwm_23__N_2951[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3090_2_lut (.I0(GND_net), .I1(n26_adj_3450), .I2(n119), 
            .I3(GND_net), .O(n8137[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_2 (.CI(GND_net), .I0(n26_adj_3450), .I1(n119), .CO(n37804));
    SB_LUT4 add_3089_26_lut (.I0(GND_net), .I1(n8137[23]), .I2(GND_net), 
            .I3(n37803), .O(n8110[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_25_lut (.I0(GND_net), .I1(n8137[22]), .I2(GND_net), 
            .I3(n37802), .O(n8110[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_25 (.CI(n37802), .I0(n8137[22]), .I1(GND_net), .CO(n37803));
    SB_LUT4 add_3089_24_lut (.I0(GND_net), .I1(n8137[21]), .I2(GND_net), 
            .I3(n37801), .O(n8110[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_24 (.CI(n37801), .I0(n8137[21]), .I1(GND_net), .CO(n37802));
    SB_LUT4 add_3089_23_lut (.I0(GND_net), .I1(n8137[20]), .I2(GND_net), 
            .I3(n37800), .O(n8110[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_23 (.CI(n37800), .I0(n8137[20]), .I1(GND_net), .CO(n37801));
    SB_CARRY mult_14_add_1211_19 (.CI(n38201), .I0(n1797[16]), .I1(GND_net), 
            .CO(n38202));
    SB_LUT4 add_3089_22_lut (.I0(GND_net), .I1(n8137[19]), .I2(GND_net), 
            .I3(n37799), .O(n8110[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_11_lut (.I0(GND_net), .I1(n16509[8]), .I2(GND_net), 
            .I3(n36831), .O(n16424[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_10_lut (.I0(GND_net), .I1(n16509[7]), .I2(GND_net), 
            .I3(n36830), .O(n16424[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_18_lut (.I0(GND_net), .I1(n1797[15]), .I2(GND_net), 
            .I3(n38200), .O(n282[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_22 (.CI(n37799), .I0(n8137[19]), .I1(GND_net), .CO(n37800));
    SB_CARRY add_3492_10 (.CI(n36830), .I0(n16509[7]), .I1(GND_net), .CO(n36831));
    SB_CARRY state_23__I_0_add_2_10 (.CI(n36654), .I0(\motor_state[8] ), 
            .I1(n70[8]), .CO(n36655));
    SB_LUT4 add_3492_9_lut (.I0(GND_net), .I1(n16509[6]), .I2(GND_net), 
            .I3(n36829), .O(n16424[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(\motor_state[7] ), 
            .I2(n70[7]), .I3(n36653), .O(\PID_CONTROLLER.err_31__N_2816 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_18 (.CI(n38200), .I0(n1797[15]), .I1(GND_net), 
            .CO(n38201));
    SB_LUT4 unary_minus_21_inv_0_i3_1_lut (.I0(\PWMLimit[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[2]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3089_21_lut (.I0(GND_net), .I1(n8137[18]), .I2(GND_net), 
            .I3(n37798), .O(n8110[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_9 (.CI(n36829), .I0(n16509[6]), .I1(GND_net), .CO(n36830));
    SB_CARRY state_23__I_0_add_2_9 (.CI(n36653), .I0(\motor_state[7] ), 
            .I1(n70[7]), .CO(n36654));
    SB_LUT4 add_3492_8_lut (.I0(GND_net), .I1(n16509[5]), .I2(n743), .I3(n36828), 
            .O(n16424[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(\motor_state[6] ), 
            .I2(n70[6]), .I3(n36652), .O(\PID_CONTROLLER.err_31__N_2816 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_17_lut (.I0(GND_net), .I1(n1797[14]), .I2(GND_net), 
            .I3(n38199), .O(n282[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_21 (.CI(n37798), .I0(n8137[18]), .I1(GND_net), .CO(n37799));
    SB_CARRY add_3492_8 (.CI(n36828), .I0(n16509[5]), .I1(n743), .CO(n36829));
    SB_CARRY state_23__I_0_add_2_8 (.CI(n36652), .I0(\motor_state[6] ), 
            .I1(n70[6]), .CO(n36653));
    SB_CARRY unary_minus_17_add_3_11 (.CI(n36540), .I0(GND_net), .I1(n69[31]), 
            .CO(n36541));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(\motor_state[5] ), 
            .I2(n70[5]), .I3(n36651), .O(\PID_CONTROLLER.err_31__N_2816 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_7_lut (.I0(GND_net), .I1(n16509[4]), .I2(n646), .I3(n36827), 
            .O(n16424[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n36651), .I0(\motor_state[5] ), 
            .I1(n70[5]), .CO(n36652));
    SB_LUT4 unary_minus_17_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n69[8]), 
            .I3(n36539), .O(pwm_23__N_2951[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_20_lut (.I0(GND_net), .I1(n8137[17]), .I2(GND_net), 
            .I3(n37797), .O(n8110[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(\motor_state[4] ), 
            .I2(n70[4]), .I3(n36650), .O(\PID_CONTROLLER.err_31__N_2816 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i247_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1211_17 (.CI(n38199), .I0(n1797[14]), .I1(GND_net), 
            .CO(n38200));
    SB_CARRY unary_minus_17_add_3_10 (.CI(n36539), .I0(GND_net), .I1(n69[8]), 
            .CO(n36540));
    SB_CARRY add_3089_20 (.CI(n37797), .I0(n8137[17]), .I1(GND_net), .CO(n37798));
    SB_CARRY add_3492_7 (.CI(n36827), .I0(n16509[4]), .I1(n646), .CO(n36828));
    SB_LUT4 mult_14_add_1211_16_lut (.I0(GND_net), .I1(n1797[13]), .I2(GND_net), 
            .I3(n38198), .O(n282[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_6_lut (.I0(GND_net), .I1(n16509[3]), .I2(n549), .I3(n36826), 
            .O(n16424[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_16 (.CI(n38198), .I0(n1797[13]), .I1(GND_net), 
            .CO(n38199));
    SB_CARRY state_23__I_0_add_2_6 (.CI(n36650), .I0(\motor_state[4] ), 
            .I1(n70[4]), .CO(n36651));
    SB_LUT4 add_3089_19_lut (.I0(GND_net), .I1(n8137[16]), .I2(GND_net), 
            .I3(n37796), .O(n8110[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_6 (.CI(n36826), .I0(n16509[3]), .I1(n549), .CO(n36827));
    SB_CARRY add_3089_19 (.CI(n37796), .I0(n8137[16]), .I1(GND_net), .CO(n37797));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(\motor_state[3] ), 
            .I2(n70[3]), .I3(n36649), .O(\PID_CONTROLLER.err_31__N_2816 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n69[7]), 
            .I3(n36538), .O(\pwm_23__N_2951[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1211_15_lut (.I0(GND_net), .I1(n1797[12]), .I2(GND_net), 
            .I3(n38197), .O(n282[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_15 (.CI(n38197), .I0(n1797[12]), .I1(GND_net), 
            .CO(n38198));
    SB_LUT4 add_3089_18_lut (.I0(GND_net), .I1(n8137[15]), .I2(GND_net), 
            .I3(n37795), .O(n8110[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_5_lut (.I0(GND_net), .I1(n16509[2]), .I2(n452_adj_3461), 
            .I3(n36825), .O(n16424[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n36649), .I0(\motor_state[3] ), 
            .I1(n70[3]), .CO(n36650));
    SB_CARRY add_3492_5 (.CI(n36825), .I0(n16509[2]), .I1(n452_adj_3461), 
            .CO(n36826));
    SB_CARRY add_3089_18 (.CI(n37795), .I0(n8137[15]), .I1(GND_net), .CO(n37796));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(\motor_state[2] ), 
            .I2(n70[2]), .I3(n36648), .O(\PID_CONTROLLER.err_31__N_2816 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_14_lut (.I0(GND_net), .I1(n1797[11]), .I2(GND_net), 
            .I3(n38196), .O(n282[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_14 (.CI(n38196), .I0(n1797[11]), .I1(GND_net), 
            .CO(n38197));
    SB_LUT4 add_3089_17_lut (.I0(GND_net), .I1(n8137[14]), .I2(GND_net), 
            .I3(n37794), .O(n8110[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_4_lut (.I0(GND_net), .I1(n16509[1]), .I2(n355), .I3(n36824), 
            .O(n16424[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_4 (.CI(n36648), .I0(\motor_state[2] ), 
            .I1(n70[2]), .CO(n36649));
    SB_CARRY unary_minus_17_add_3_9 (.CI(n36538), .I0(GND_net), .I1(n69[7]), 
            .CO(n36539));
    SB_CARRY add_3089_17 (.CI(n37794), .I0(n8137[14]), .I1(GND_net), .CO(n37795));
    SB_LUT4 unary_minus_17_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n69[6]), 
            .I3(n36537), .O(pwm_23__N_2951[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(\motor_state[1] ), 
            .I2(n70[1]), .I3(n36647), .O(\PID_CONTROLLER.err_31__N_2816 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_16_lut (.I0(GND_net), .I1(n8137[13]), .I2(GND_net), 
            .I3(n37793), .O(n8110[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_4 (.CI(n36824), .I0(n16509[1]), .I1(n355), .CO(n36825));
    SB_CARRY state_23__I_0_add_2_3 (.CI(n36647), .I0(\motor_state[1] ), 
            .I1(n70[1]), .CO(n36648));
    SB_LUT4 mult_14_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1211_13_lut (.I0(GND_net), .I1(n1797[10]), .I2(GND_net), 
            .I3(n38195), .O(n282[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_13 (.CI(n38195), .I0(n1797[10]), .I1(GND_net), 
            .CO(n38196));
    SB_LUT4 mult_14_add_1211_12_lut (.I0(GND_net), .I1(n1797[9]), .I2(GND_net), 
            .I3(n38194), .O(n282[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_3_lut (.I0(GND_net), .I1(n16509[0]), .I2(n258), .I3(n36823), 
            .O(n16424[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_12 (.CI(n38194), .I0(n1797[9]), .I1(GND_net), 
            .CO(n38195));
    SB_LUT4 mult_14_add_1211_11_lut (.I0(GND_net), .I1(n1797[8]), .I2(GND_net), 
            .I3(n38193), .O(n282[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_11 (.CI(n38193), .I0(n1797[8]), .I1(GND_net), 
            .CO(n38194));
    SB_LUT4 mult_14_add_1211_10_lut (.I0(GND_net), .I1(n1797[7]), .I2(GND_net), 
            .I3(n38192), .O(n282[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_10 (.CI(n38192), .I0(n1797[7]), .I1(GND_net), 
            .CO(n38193));
    SB_LUT4 mult_14_add_1211_9_lut (.I0(GND_net), .I1(n1797[6]), .I2(GND_net), 
            .I3(n38191), .O(n282[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_9 (.CI(n38191), .I0(n1797[6]), .I1(GND_net), 
            .CO(n38192));
    SB_LUT4 mult_10_i174_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n258));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1211_8_lut (.I0(GND_net), .I1(n1797[5]), .I2(n512), 
            .I3(n38190), .O(n282[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_8 (.CI(n38190), .I0(n1797[5]), .I1(n512), 
            .CO(n38191));
    SB_LUT4 mult_14_add_1211_7_lut (.I0(GND_net), .I1(n1797[4]), .I2(n439), 
            .I3(n38189), .O(n282[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_7 (.CI(n38189), .I0(n1797[4]), .I1(n439), 
            .CO(n38190));
    SB_LUT4 mult_14_add_1211_6_lut (.I0(GND_net), .I1(n1797[3]), .I2(n366), 
            .I3(n38188), .O(n282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_6 (.CI(n38188), .I0(n1797[3]), .I1(n366), 
            .CO(n38189));
    SB_LUT4 mult_14_add_1211_5_lut (.I0(GND_net), .I1(n1797[2]), .I2(n293), 
            .I3(n38187), .O(n282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_16 (.CI(n37793), .I0(n8137[13]), .I1(GND_net), .CO(n37794));
    SB_CARRY mult_14_add_1211_5 (.CI(n38187), .I0(n1797[2]), .I1(n293), 
            .CO(n38188));
    SB_LUT4 mult_14_add_1211_4_lut (.I0(GND_net), .I1(n1797[1]), .I2(n220), 
            .I3(n38186), .O(n282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_4 (.CI(n38186), .I0(n1797[1]), .I1(n220), 
            .CO(n38187));
    SB_LUT4 mult_14_add_1211_3_lut (.I0(GND_net), .I1(n1797[0]), .I2(n147), 
            .I3(n38185), .O(n282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_3 (.CI(n38185), .I0(n1797[0]), .I1(n147), 
            .CO(n38186));
    SB_LUT4 mult_14_add_1211_2_lut (.I0(GND_net), .I1(n5_adj_3439), .I2(n74), 
            .I3(GND_net), .O(n282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_2 (.CI(GND_net), .I0(n5_adj_3439), .I1(n74), 
            .CO(n38185));
    SB_LUT4 add_3400_18_lut (.I0(GND_net), .I1(n15403[15]), .I2(GND_net), 
            .I3(n38184), .O(n15118[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_17_lut (.I0(GND_net), .I1(n15403[14]), .I2(GND_net), 
            .I3(n38183), .O(n15118[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_3 (.CI(n36823), .I0(n16509[0]), .I1(n258), .CO(n36824));
    SB_CARRY unary_minus_17_add_3_8 (.CI(n36537), .I0(GND_net), .I1(n69[6]), 
            .CO(n36538));
    SB_LUT4 add_3089_15_lut (.I0(GND_net), .I1(n8137[12]), .I2(GND_net), 
            .I3(n37792), .O(n8110[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_2_lut (.I0(GND_net), .I1(n68), .I2(n161), .I3(GND_net), 
            .O(n16424[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n69[5]), 
            .I3(n36536), .O(\pwm_23__N_2951[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_17 (.CI(n38183), .I0(n15403[14]), .I1(GND_net), 
            .CO(n38184));
    SB_CARRY add_3492_2 (.CI(GND_net), .I0(n68), .I1(n161), .CO(n36823));
    SB_CARRY add_3089_15 (.CI(n37792), .I0(n8137[12]), .I1(GND_net), .CO(n37793));
    SB_LUT4 add_3343_21_lut (.I0(GND_net), .I1(n14438[18]), .I2(GND_net), 
            .I3(n36822), .O(n14039[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_16_lut (.I0(GND_net), .I1(n15403[13]), .I2(GND_net), 
            .I3(n38182), .O(n15118[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_16 (.CI(n38182), .I0(n15403[13]), .I1(GND_net), 
            .CO(n38183));
    SB_LUT4 add_3400_15_lut (.I0(GND_net), .I1(n15403[12]), .I2(GND_net), 
            .I3(n38181), .O(n15118[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_7 (.CI(n36536), .I0(GND_net), .I1(n69[5]), 
            .CO(n36537));
    SB_CARRY add_3400_15 (.CI(n38181), .I0(n15403[12]), .I1(GND_net), 
            .CO(n38182));
    SB_LUT4 add_3400_14_lut (.I0(GND_net), .I1(n15403[11]), .I2(GND_net), 
            .I3(n38180), .O(n15118[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_14 (.CI(n38180), .I0(n15403[11]), .I1(GND_net), 
            .CO(n38181));
    SB_LUT4 add_3400_13_lut (.I0(GND_net), .I1(n15403[10]), .I2(GND_net), 
            .I3(n38179), .O(n15118[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_13 (.CI(n38179), .I0(n15403[10]), .I1(GND_net), 
            .CO(n38180));
    SB_LUT4 add_3400_12_lut (.I0(GND_net), .I1(n15403[9]), .I2(GND_net), 
            .I3(n38178), .O(n15118[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_12 (.CI(n38178), .I0(n15403[9]), .I1(GND_net), .CO(n38179));
    SB_LUT4 add_3400_11_lut (.I0(GND_net), .I1(n15403[8]), .I2(GND_net), 
            .I3(n38177), .O(n15118[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_11 (.CI(n38177), .I0(n15403[8]), .I1(GND_net), .CO(n38178));
    SB_LUT4 add_3400_10_lut (.I0(GND_net), .I1(n15403[7]), .I2(GND_net), 
            .I3(n38176), .O(n15118[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_10 (.CI(n38176), .I0(n15403[7]), .I1(GND_net), .CO(n38177));
    SB_LUT4 add_3400_9_lut (.I0(GND_net), .I1(n15403[6]), .I2(GND_net), 
            .I3(n38175), .O(n15118[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_9 (.CI(n38175), .I0(n15403[6]), .I1(GND_net), .CO(n38176));
    SB_LUT4 add_3400_8_lut (.I0(GND_net), .I1(n15403[5]), .I2(n722), .I3(n38174), 
            .O(n15118[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_8 (.CI(n38174), .I0(n15403[5]), .I1(n722), .CO(n38175));
    SB_LUT4 add_3400_7_lut (.I0(GND_net), .I1(n15403[4]), .I2(n625), .I3(n38173), 
            .O(n15118[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_7 (.CI(n38173), .I0(n15403[4]), .I1(n625), .CO(n38174));
    SB_LUT4 add_3400_6_lut (.I0(GND_net), .I1(n15403[3]), .I2(n528_adj_3419), 
            .I3(n38172), .O(n15118[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_6 (.CI(n38172), .I0(n15403[3]), .I1(n528_adj_3419), 
            .CO(n38173));
    SB_LUT4 add_3400_5_lut (.I0(GND_net), .I1(n15403[2]), .I2(n431), .I3(n38171), 
            .O(n15118[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_5 (.CI(n38171), .I0(n15403[2]), .I1(n431), .CO(n38172));
    SB_LUT4 add_3400_4_lut (.I0(GND_net), .I1(n15403[1]), .I2(n334), .I3(n38170), 
            .O(n15118[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_4 (.CI(n38170), .I0(n15403[1]), .I1(n334), .CO(n38171));
    SB_LUT4 add_3400_3_lut (.I0(GND_net), .I1(n15403[0]), .I2(n237), .I3(n38169), 
            .O(n15118[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_3 (.CI(n38169), .I0(n15403[0]), .I1(n237), .CO(n38170));
    SB_LUT4 add_3400_2_lut (.I0(GND_net), .I1(n47), .I2(n140), .I3(GND_net), 
            .O(n15118[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_2 (.CI(GND_net), .I0(n47), .I1(n140), .CO(n38169));
    SB_LUT4 add_3509_9_lut (.I0(GND_net), .I1(n16624[6]), .I2(GND_net), 
            .I3(n38168), .O(n16575[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3509_8_lut (.I0(GND_net), .I1(n16624[5]), .I2(n749), .I3(n38167), 
            .O(n16575[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3509_8 (.CI(n38167), .I0(n16624[5]), .I1(n749), .CO(n38168));
    SB_LUT4 add_3509_7_lut (.I0(GND_net), .I1(n16624[4]), .I2(n652), .I3(n38166), 
            .O(n16575[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3509_7 (.CI(n38166), .I0(n16624[4]), .I1(n652), .CO(n38167));
    SB_LUT4 add_3089_14_lut (.I0(GND_net), .I1(n8137[11]), .I2(GND_net), 
            .I3(n37791), .O(n8110[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3509_6_lut (.I0(GND_net), .I1(n16624[3]), .I2(n555), .I3(n38165), 
            .O(n16575[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_14 (.CI(n37791), .I0(n8137[11]), .I1(GND_net), .CO(n37792));
    SB_LUT4 add_3089_13_lut (.I0(GND_net), .I1(n8137[10]), .I2(GND_net), 
            .I3(n37790), .O(n8110[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3509_6 (.CI(n38165), .I0(n16624[3]), .I1(n555), .CO(n38166));
    SB_LUT4 add_3509_5_lut (.I0(GND_net), .I1(n16624[2]), .I2(n458_c), 
            .I3(n38164), .O(n16575[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_13 (.CI(n37790), .I0(n8137[10]), .I1(GND_net), .CO(n37791));
    SB_CARRY add_3509_5 (.CI(n38164), .I0(n16624[2]), .I1(n458_c), .CO(n38165));
    SB_LUT4 add_3343_20_lut (.I0(GND_net), .I1(n14438[17]), .I2(GND_net), 
            .I3(n36821), .O(n14039[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3509_4_lut (.I0(GND_net), .I1(n16624[1]), .I2(n361), .I3(n38163), 
            .O(n16575[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3509_4 (.CI(n38163), .I0(n16624[1]), .I1(n361), .CO(n38164));
    SB_LUT4 add_3089_12_lut (.I0(GND_net), .I1(n8137[9]), .I2(GND_net), 
            .I3(n37789), .O(n8110[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3509_3_lut (.I0(GND_net), .I1(n16624[0]), .I2(n264), .I3(n38162), 
            .O(n16575[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[1]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3509_3 (.CI(n38162), .I0(n16624[0]), .I1(n264), .CO(n38163));
    SB_CARRY add_3089_12 (.CI(n37789), .I0(n8137[9]), .I1(GND_net), .CO(n37790));
    SB_LUT4 add_3509_2_lut (.I0(GND_net), .I1(n86_adj_3409), .I2(n167), 
            .I3(GND_net), .O(n16575[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_11_lut (.I0(GND_net), .I1(n8137[8]), .I2(GND_net), 
            .I3(n37788), .O(n8110[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3509_2 (.CI(GND_net), .I0(n86_adj_3409), .I1(n167), .CO(n38162));
    SB_CARRY add_3089_11 (.CI(n37788), .I0(n8137[8]), .I1(GND_net), .CO(n37789));
    SB_LUT4 add_3417_17_lut (.I0(GND_net), .I1(n15644[14]), .I2(GND_net), 
            .I3(n38161), .O(n15403[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_10_lut (.I0(GND_net), .I1(n8137[7]), .I2(GND_net), 
            .I3(n37787), .O(n8110[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3417_16_lut (.I0(GND_net), .I1(n15644[13]), .I2(GND_net), 
            .I3(n38160), .O(n15403[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_16 (.CI(n38160), .I0(n15644[13]), .I1(GND_net), 
            .CO(n38161));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(\motor_state[0] ), 
            .I2(n70[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_31__N_2816 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_20 (.CI(n36821), .I0(n14438[17]), .I1(GND_net), 
            .CO(n36822));
    SB_LUT4 add_3343_19_lut (.I0(GND_net), .I1(n14438[16]), .I2(GND_net), 
            .I3(n36820), .O(n14039[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_10 (.CI(n37787), .I0(n8137[7]), .I1(GND_net), .CO(n37788));
    SB_LUT4 add_3089_9_lut (.I0(GND_net), .I1(n8137[6]), .I2(GND_net), 
            .I3(n37786), .O(n8110[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_9 (.CI(n37786), .I0(n8137[6]), .I1(GND_net), .CO(n37787));
    SB_LUT4 add_3417_15_lut (.I0(GND_net), .I1(n15644[12]), .I2(GND_net), 
            .I3(n38159), .O(n15403[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_8_lut (.I0(GND_net), .I1(n8137[5]), .I2(n698), .I3(n37785), 
            .O(n8110[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n69[4]), 
            .I3(n36535), .O(\pwm_23__N_2951[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_8 (.CI(n37785), .I0(n8137[5]), .I1(n698), .CO(n37786));
    SB_CARRY add_3417_15 (.CI(n38159), .I0(n15644[12]), .I1(GND_net), 
            .CO(n38160));
    SB_LUT4 add_3089_7_lut (.I0(GND_net), .I1(n8137[4]), .I2(n601_adj_3380), 
            .I3(n37784), .O(n8110[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3417_14_lut (.I0(GND_net), .I1(n15644[11]), .I2(GND_net), 
            .I3(n38158), .O(n15403[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_7 (.CI(n37784), .I0(n8137[4]), .I1(n601_adj_3380), 
            .CO(n37785));
    SB_CARRY add_3417_14 (.CI(n38158), .I0(n15644[11]), .I1(GND_net), 
            .CO(n38159));
    SB_LUT4 add_3089_6_lut (.I0(GND_net), .I1(n8137[3]), .I2(n504), .I3(n37783), 
            .O(n8110[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(\motor_state[0] ), 
            .I1(n70[0]), .CO(n36647));
    SB_CARRY unary_minus_17_add_3_6 (.CI(n36535), .I0(GND_net), .I1(n69[4]), 
            .CO(n36536));
    SB_CARRY add_3089_6 (.CI(n37783), .I0(n8137[3]), .I1(n504), .CO(n37784));
    SB_LUT4 add_3089_5_lut (.I0(GND_net), .I1(n8137[2]), .I2(n407), .I3(n37782), 
            .O(n8110[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n69[3]), 
            .I3(n36534), .O(pwm_23__N_2951[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3417_13_lut (.I0(GND_net), .I1(n15644[10]), .I2(GND_net), 
            .I3(n38157), .O(n15403[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_5 (.CI(n37782), .I0(n8137[2]), .I1(n407), .CO(n37783));
    SB_CARRY add_3417_13 (.CI(n38157), .I0(n15644[10]), .I1(GND_net), 
            .CO(n38158));
    SB_LUT4 unary_minus_17_inv_0_i7_1_lut (.I0(\deadband[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[6]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3089_4_lut (.I0(GND_net), .I1(n8137[1]), .I2(n310), .I3(n37781), 
            .O(n8110[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_4 (.CI(n37781), .I0(n8137[1]), .I1(n310), .CO(n37782));
    SB_LUT4 add_3417_12_lut (.I0(GND_net), .I1(n15644[9]), .I2(GND_net), 
            .I3(n38156), .O(n15403[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_3_lut (.I0(GND_net), .I1(n8137[0]), .I2(n213), .I3(n37780), 
            .O(n8110[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_5 (.CI(n36534), .I0(GND_net), .I1(n69[3]), 
            .CO(n36535));
    SB_LUT4 mult_10_i239_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n355));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i239_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3417_12 (.CI(n38156), .I0(n15644[9]), .I1(GND_net), .CO(n38157));
    SB_LUT4 add_3417_11_lut (.I0(GND_net), .I1(n15644[8]), .I2(GND_net), 
            .I3(n38155), .O(n15403[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_11 (.CI(n38155), .I0(n15644[8]), .I1(GND_net), .CO(n38156));
    SB_CARRY add_3089_3 (.CI(n37780), .I0(n8137[0]), .I1(n213), .CO(n37781));
    SB_LUT4 add_3417_10_lut (.I0(GND_net), .I1(n15644[7]), .I2(GND_net), 
            .I3(n38154), .O(n15403[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_2_lut (.I0(GND_net), .I1(n23_c), .I2(n116), .I3(GND_net), 
            .O(n8110[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[2]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3089_2 (.CI(GND_net), .I0(n23_c), .I1(n116), .CO(n37780));
    SB_LUT4 add_3088_27_lut (.I0(GND_net), .I1(n8110[24]), .I2(GND_net), 
            .I3(n37779), .O(n8082[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_19 (.CI(n36820), .I0(n14438[16]), .I1(GND_net), 
            .CO(n36821));
    SB_CARRY add_3417_10 (.CI(n38154), .I0(n15644[7]), .I1(GND_net), .CO(n38155));
    SB_LUT4 add_3088_26_lut (.I0(GND_net), .I1(n8110[23]), .I2(GND_net), 
            .I3(n37778), .O(n8082[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_18_lut (.I0(GND_net), .I1(n14438[15]), .I2(GND_net), 
            .I3(n36819), .O(n14039[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_26 (.CI(n37778), .I0(n8110[23]), .I1(GND_net), .CO(n37779));
    SB_LUT4 add_3088_25_lut (.I0(GND_net), .I1(n8110[22]), .I2(GND_net), 
            .I3(n37777), .O(n8082[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_27_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n66[26]), .I3(n36646), .O(n67[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3417_9_lut (.I0(GND_net), .I1(n15644[6]), .I2(GND_net), 
            .I3(n38153), .O(n15403[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_25 (.CI(n37777), .I0(n8110[22]), .I1(GND_net), .CO(n37778));
    SB_CARRY add_3417_9 (.CI(n38153), .I0(n15644[6]), .I1(GND_net), .CO(n38154));
    SB_LUT4 add_3088_24_lut (.I0(GND_net), .I1(n8110[21]), .I2(GND_net), 
            .I3(n37776), .O(n8082[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_24 (.CI(n37776), .I0(n8110[21]), .I1(GND_net), .CO(n37777));
    SB_LUT4 add_3088_23_lut (.I0(GND_net), .I1(n8110[20]), .I2(GND_net), 
            .I3(n37775), .O(n8082[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3417_8_lut (.I0(GND_net), .I1(n15644[5]), .I2(n725), .I3(n38152), 
            .O(n15403[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_23 (.CI(n37775), .I0(n8110[20]), .I1(GND_net), .CO(n37776));
    SB_CARRY add_3417_8 (.CI(n38152), .I0(n15644[5]), .I1(n725), .CO(n38153));
    SB_LUT4 add_3417_7_lut (.I0(GND_net), .I1(n15644[4]), .I2(n628), .I3(n38151), 
            .O(n15403[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_7 (.CI(n38151), .I0(n15644[4]), .I1(n628), .CO(n38152));
    SB_LUT4 add_3417_6_lut (.I0(GND_net), .I1(n15644[3]), .I2(n531), .I3(n38150), 
            .O(n15403[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_6 (.CI(n38150), .I0(n15644[3]), .I1(n531), .CO(n38151));
    SB_LUT4 add_3417_5_lut (.I0(GND_net), .I1(n15644[2]), .I2(n434), .I3(n38149), 
            .O(n15403[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_5 (.CI(n38149), .I0(n15644[2]), .I1(n434), .CO(n38150));
    SB_LUT4 add_3417_4_lut (.I0(GND_net), .I1(n15644[1]), .I2(n337), .I3(n38148), 
            .O(n15403[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_4 (.CI(n38148), .I0(n15644[1]), .I1(n337), .CO(n38149));
    SB_LUT4 add_3417_3_lut (.I0(GND_net), .I1(n15644[0]), .I2(n240), .I3(n38147), 
            .O(n15403[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_3 (.CI(n38147), .I0(n15644[0]), .I1(n240), .CO(n38148));
    SB_LUT4 add_3417_2_lut (.I0(GND_net), .I1(n50), .I2(n143), .I3(GND_net), 
            .O(n15403[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n452_adj_3461));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3417_2 (.CI(GND_net), .I0(n50), .I1(n143), .CO(n38147));
    SB_LUT4 add_3517_7_lut (.I0(GND_net), .I1(n43817), .I2(n658), .I3(n38146), 
            .O(n16633[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3517_6_lut (.I0(GND_net), .I1(n16641[3]), .I2(n558), .I3(n38145), 
            .O(n16633[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_6 (.CI(n38145), .I0(n16641[3]), .I1(n558), .CO(n38146));
    SB_LUT4 add_3088_22_lut (.I0(GND_net), .I1(n8110[19]), .I2(GND_net), 
            .I3(n37774), .O(n8082[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_22 (.CI(n37774), .I0(n8110[19]), .I1(GND_net), .CO(n37775));
    SB_LUT4 add_3088_21_lut (.I0(GND_net), .I1(n8110[18]), .I2(GND_net), 
            .I3(n37773), .O(n8082[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_21 (.CI(n37773), .I0(n8110[18]), .I1(GND_net), .CO(n37774));
    SB_LUT4 add_3088_20_lut (.I0(GND_net), .I1(n8110[17]), .I2(GND_net), 
            .I3(n37772), .O(n8082[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_20 (.CI(n37772), .I0(n8110[17]), .I1(GND_net), .CO(n37773));
    SB_LUT4 unary_minus_17_inv_0_i8_1_lut (.I0(\deadband[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[7]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3088_19_lut (.I0(GND_net), .I1(n8110[16]), .I2(GND_net), 
            .I3(n37771), .O(n8082[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_19 (.CI(n37771), .I0(n8110[16]), .I1(GND_net), .CO(n37772));
    SB_LUT4 add_3088_18_lut (.I0(GND_net), .I1(n8110[15]), .I2(GND_net), 
            .I3(n37770), .O(n8082[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_18 (.CI(n37770), .I0(n8110[15]), .I1(GND_net), .CO(n37771));
    SB_LUT4 add_3088_17_lut (.I0(GND_net), .I1(n8110[14]), .I2(GND_net), 
            .I3(n37769), .O(n8082[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_17 (.CI(n37769), .I0(n8110[14]), .I1(GND_net), .CO(n37770));
    SB_LUT4 add_3088_16_lut (.I0(GND_net), .I1(n8110[13]), .I2(GND_net), 
            .I3(n37768), .O(n8082[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_16 (.CI(n37768), .I0(n8110[13]), .I1(GND_net), .CO(n37769));
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[3]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3088_15_lut (.I0(GND_net), .I1(n8110[12]), .I2(GND_net), 
            .I3(n37767), .O(n8082[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_15 (.CI(n37767), .I0(n8110[12]), .I1(GND_net), .CO(n37768));
    SB_LUT4 add_3517_5_lut (.I0(GND_net), .I1(n16641[2]), .I2(n464), .I3(n38144), 
            .O(n16633[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_14_lut (.I0(GND_net), .I1(n8110[11]), .I2(GND_net), 
            .I3(n37766), .O(n8082[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_14 (.CI(n37766), .I0(n8110[11]), .I1(GND_net), .CO(n37767));
    SB_CARRY add_3517_5 (.CI(n38144), .I0(n16641[2]), .I1(n464), .CO(n38145));
    SB_LUT4 add_3088_13_lut (.I0(GND_net), .I1(n8110[10]), .I2(GND_net), 
            .I3(n37765), .O(n8082[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_13 (.CI(n37765), .I0(n8110[10]), .I1(GND_net), .CO(n37766));
    SB_LUT4 add_3517_4_lut (.I0(GND_net), .I1(n16654[1]), .I2(n370_adj_3471), 
            .I3(n38143), .O(n16633[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_12_lut (.I0(GND_net), .I1(n8110[9]), .I2(GND_net), 
            .I3(n37764), .O(n8082[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_12 (.CI(n37764), .I0(n8110[9]), .I1(GND_net), .CO(n37765));
    SB_CARRY add_3517_4 (.CI(n38143), .I0(n16654[1]), .I1(n370_adj_3471), 
            .CO(n38144));
    SB_LUT4 add_3088_11_lut (.I0(GND_net), .I1(n8110[8]), .I2(GND_net), 
            .I3(n37763), .O(n8082[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_11 (.CI(n37763), .I0(n8110[8]), .I1(GND_net), .CO(n37764));
    SB_LUT4 add_3088_10_lut (.I0(GND_net), .I1(n8110[7]), .I2(GND_net), 
            .I3(n37762), .O(n8082[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_26_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n66[26]), .I3(n36645), .O(n67[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n69[2]), 
            .I3(n36533), .O(pwm_23__N_2951[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3517_3_lut (.I0(GND_net), .I1(n16641[0]), .I2(n276), .I3(n38142), 
            .O(n16633[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_10 (.CI(n37762), .I0(n8110[7]), .I1(GND_net), .CO(n37763));
    SB_CARRY add_3517_3 (.CI(n38142), .I0(n16641[0]), .I1(n276), .CO(n38143));
    SB_CARRY unary_minus_17_add_3_4 (.CI(n36533), .I0(GND_net), .I1(n69[2]), 
            .CO(n36534));
    SB_CARRY sub_11_add_2_26 (.CI(n36645), .I0(\PID_CONTROLLER.err_prev[31] ), 
            .I1(n66[26]), .CO(n36646));
    SB_LUT4 unary_minus_17_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n69[1]), 
            .I3(n36532), .O(pwm_23__N_2951[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_3 (.CI(n36532), .I0(GND_net), .I1(n69[1]), 
            .CO(n36533));
    SB_LUT4 unary_minus_17_add_3_2_lut (.I0(n28960), .I1(GND_net), .I2(n69[0]), 
            .I3(VCC_net), .O(n46507)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3517_2_lut (.I0(GND_net), .I1(n86_adj_3409), .I2(n182), 
            .I3(GND_net), .O(n16633[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[23] ), 
            .I2(n66[23]), .I3(n36644), .O(n67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_9_lut (.I0(GND_net), .I1(n8110[6]), .I2(GND_net), 
            .I3(n37761), .O(n8082[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3517_2 (.CI(GND_net), .I0(n86_adj_3409), .I1(n182), .CO(n38142));
    SB_CARRY unary_minus_17_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n69[0]), 
            .CO(n36532));
    SB_LUT4 add_3432_16_lut (.I0(GND_net), .I1(n15854[13]), .I2(GND_net), 
            .I3(n38141), .O(n15644[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_9 (.CI(n37761), .I0(n8110[6]), .I1(GND_net), .CO(n37762));
    SB_LUT4 add_3088_8_lut (.I0(GND_net), .I1(n8110[5]), .I2(n695), .I3(n37760), 
            .O(n8082[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_8 (.CI(n37760), .I0(n8110[5]), .I1(n695), .CO(n37761));
    SB_CARRY add_3343_18 (.CI(n36819), .I0(n14438[15]), .I1(GND_net), 
            .CO(n36820));
    SB_LUT4 add_3088_7_lut (.I0(GND_net), .I1(n8110[4]), .I2(n598_adj_3477), 
            .I3(n37759), .O(n8082[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_25 (.CI(n36644), .I0(\PID_CONTROLLER.err_prev[23] ), 
            .I1(n66[23]), .CO(n36645));
    SB_LUT4 add_3432_15_lut (.I0(GND_net), .I1(n15854[12]), .I2(GND_net), 
            .I3(n38140), .O(n15644[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_7 (.CI(n37759), .I0(n8110[4]), .I1(n598_adj_3477), 
            .CO(n37760));
    SB_LUT4 add_3088_6_lut (.I0(GND_net), .I1(n8110[3]), .I2(n501), .I3(n37758), 
            .O(n8082[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[22] ), 
            .I2(n66[22]), .I3(n36643), .O(n67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_6 (.CI(n37758), .I0(n8110[3]), .I1(n501), .CO(n37759));
    SB_LUT4 add_3343_17_lut (.I0(GND_net), .I1(n14438[14]), .I2(GND_net), 
            .I3(n36818), .O(n14039[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_17 (.CI(n36818), .I0(n14438[14]), .I1(GND_net), 
            .CO(n36819));
    SB_CARRY add_3432_15 (.CI(n38140), .I0(n15854[12]), .I1(GND_net), 
            .CO(n38141));
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n549));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3432_14_lut (.I0(GND_net), .I1(n15854[11]), .I2(GND_net), 
            .I3(n38139), .O(n15644[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_5_lut (.I0(GND_net), .I1(n8110[2]), .I2(n404), .I3(n37757), 
            .O(n8082[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_5 (.CI(n37757), .I0(n8110[2]), .I1(n404), .CO(n37758));
    SB_LUT4 add_3088_4_lut (.I0(GND_net), .I1(n8110[1]), .I2(n307_adj_3479), 
            .I3(n37756), .O(n8082[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_4 (.CI(n37756), .I0(n8110[1]), .I1(n307_adj_3479), 
            .CO(n37757));
    SB_LUT4 add_3088_3_lut (.I0(GND_net), .I1(n8110[0]), .I2(n210), .I3(n37755), 
            .O(n8082[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_14 (.CI(n38139), .I0(n15854[11]), .I1(GND_net), 
            .CO(n38140));
    SB_CARRY add_3088_3 (.CI(n37755), .I0(n8110[0]), .I1(n210), .CO(n37756));
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[4]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3088_2_lut (.I0(GND_net), .I1(n20_adj_3480), .I2(n113), 
            .I3(GND_net), .O(n8082[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_2 (.CI(GND_net), .I0(n20_adj_3480), .I1(n113), .CO(n37755));
    SB_LUT4 add_3432_13_lut (.I0(GND_net), .I1(n15854[10]), .I2(GND_net), 
            .I3(n38138), .O(n15644[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_28_lut (.I0(GND_net), .I1(n8082[25]), .I2(GND_net), 
            .I3(n37754), .O(n8053[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_27_lut (.I0(GND_net), .I1(n8082[24]), .I2(GND_net), 
            .I3(n37753), .O(n8053[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_27 (.CI(n37753), .I0(n8082[24]), .I1(GND_net), .CO(n37754));
    SB_CARRY add_3432_13 (.CI(n38138), .I0(n15854[10]), .I1(GND_net), 
            .CO(n38139));
    SB_LUT4 add_3087_26_lut (.I0(GND_net), .I1(n8082[23]), .I2(GND_net), 
            .I3(n37752), .O(n8053[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_26 (.CI(n37752), .I0(n8082[23]), .I1(GND_net), .CO(n37753));
    SB_LUT4 add_3432_12_lut (.I0(GND_net), .I1(n15854[9]), .I2(GND_net), 
            .I3(n38137), .O(n15644[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_12 (.CI(n38137), .I0(n15854[9]), .I1(GND_net), .CO(n38138));
    SB_CARRY sub_11_add_2_24 (.CI(n36643), .I0(\PID_CONTROLLER.err_prev[22] ), 
            .I1(n66[22]), .CO(n36644));
    SB_LUT4 add_3087_25_lut (.I0(GND_net), .I1(n8082[22]), .I2(GND_net), 
            .I3(n37751), .O(n8053[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(n19326), .I1(n881_adj_3481), .I2(n16802), 
            .I3(n17_adj_3482), .O(n43915));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3087_25 (.CI(n37751), .I0(n8082[22]), .I1(GND_net), .CO(n37752));
    SB_LUT4 add_3087_24_lut (.I0(GND_net), .I1(n8082[21]), .I2(GND_net), 
            .I3(n37750), .O(n8053[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3432_11_lut (.I0(GND_net), .I1(n15854[8]), .I2(GND_net), 
            .I3(n38136), .O(n15644[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_24 (.CI(n37750), .I0(n8082[21]), .I1(GND_net), .CO(n37751));
    SB_LUT4 add_3087_23_lut (.I0(GND_net), .I1(n8082[20]), .I2(GND_net), 
            .I3(n37749), .O(n8053[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_23 (.CI(n37749), .I0(n8082[20]), .I1(GND_net), .CO(n37750));
    SB_LUT4 add_3087_22_lut (.I0(GND_net), .I1(n8082[19]), .I2(GND_net), 
            .I3(n37748), .O(n8053[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[21] ), 
            .I2(n66[21]), .I3(n36642), .O(n67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_22 (.CI(n37748), .I0(n8082[19]), .I1(GND_net), .CO(n37749));
    SB_CARRY add_3432_11 (.CI(n38136), .I0(n15854[8]), .I1(GND_net), .CO(n38137));
    SB_LUT4 add_3087_21_lut (.I0(GND_net), .I1(n8082[18]), .I2(GND_net), 
            .I3(n37747), .O(n8053[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_23 (.CI(n36642), .I0(\PID_CONTROLLER.err_prev[21] ), 
            .I1(n66[21]), .CO(n36643));
    SB_CARRY add_3087_21 (.CI(n37747), .I0(n8082[18]), .I1(GND_net), .CO(n37748));
    SB_LUT4 sub_11_add_2_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[20] ), 
            .I2(n66[20]), .I3(n36641), .O(n67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i4_1_lut (.I0(\PWMLimit[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[3]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3432_10_lut (.I0(GND_net), .I1(n15854[7]), .I2(GND_net), 
            .I3(n38135), .O(n15644[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_20_lut (.I0(GND_net), .I1(n8082[17]), .I2(GND_net), 
            .I3(n37746), .O(n8053[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3052_10_lut (.I0(GND_net), .I1(n1804[22]), .I2(n1711), 
            .I3(n38418), .O(n7069[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i9_1_lut (.I0(\deadband[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[8]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3432_10 (.CI(n38135), .I0(n15854[7]), .I1(GND_net), .CO(n38136));
    SB_LUT4 add_3432_9_lut (.I0(GND_net), .I1(n15854[6]), .I2(GND_net), 
            .I3(n38134), .O(n15644[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_20 (.CI(n37746), .I0(n8082[17]), .I1(GND_net), .CO(n37747));
    SB_CARRY sub_11_add_2_22 (.CI(n36641), .I0(\PID_CONTROLLER.err_prev[20] ), 
            .I1(n66[20]), .CO(n36642));
    SB_LUT4 sub_11_add_2_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[19] ), 
            .I2(n66[19]), .I3(n36640), .O(n67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3052_9_lut (.I0(GND_net), .I1(n1803[22]), .I2(n1707), 
            .I3(n38417), .O(n7069[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_9 (.CI(n38134), .I0(n15854[6]), .I1(GND_net), .CO(n38135));
    SB_CARRY add_3052_9 (.CI(n38417), .I0(n1803[22]), .I1(n1707), .CO(n38418));
    SB_LUT4 add_3432_8_lut (.I0(GND_net), .I1(n15854[5]), .I2(n728), .I3(n38133), 
            .O(n15644[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_8 (.CI(n38133), .I0(n15854[5]), .I1(n728), .CO(n38134));
    SB_LUT4 add_3087_19_lut (.I0(GND_net), .I1(n8082[16]), .I2(GND_net), 
            .I3(n37745), .O(n8053[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i434_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n646));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i434_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_11_add_2_21 (.CI(n36640), .I0(\PID_CONTROLLER.err_prev[19] ), 
            .I1(n66[19]), .CO(n36641));
    SB_LUT4 sub_11_add_2_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[18] ), 
            .I2(n66[18]), .I3(n36639), .O(n67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_19 (.CI(n37745), .I0(n8082[16]), .I1(GND_net), .CO(n37746));
    SB_LUT4 add_3087_18_lut (.I0(GND_net), .I1(n8082[15]), .I2(GND_net), 
            .I3(n37744), .O(n8053[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[5]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3087_18 (.CI(n37744), .I0(n8082[15]), .I1(GND_net), .CO(n37745));
    SB_CARRY sub_11_add_2_20 (.CI(n36639), .I0(\PID_CONTROLLER.err_prev[18] ), 
            .I1(n66[18]), .CO(n36640));
    SB_LUT4 add_3432_7_lut (.I0(GND_net), .I1(n15854[4]), .I2(n631), .I3(n38132), 
            .O(n15644[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_7 (.CI(n38132), .I0(n15854[4]), .I1(n631), .CO(n38133));
    SB_LUT4 add_3432_6_lut (.I0(GND_net), .I1(n15854[3]), .I2(n534), .I3(n38131), 
            .O(n15644[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[6]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3087_17_lut (.I0(GND_net), .I1(n8082[14]), .I2(GND_net), 
            .I3(n37743), .O(n8053[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_17 (.CI(n37743), .I0(n8082[14]), .I1(GND_net), .CO(n37744));
    SB_LUT4 add_3087_16_lut (.I0(GND_net), .I1(n8082[13]), .I2(GND_net), 
            .I3(n37742), .O(n8053[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[17] ), 
            .I2(n66[17]), .I3(n36638), .O(n67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_6 (.CI(n38131), .I0(n15854[3]), .I1(n534), .CO(n38132));
    SB_CARRY add_3087_16 (.CI(n37742), .I0(n8082[13]), .I1(GND_net), .CO(n37743));
    SB_LUT4 add_3087_15_lut (.I0(GND_net), .I1(n8082[12]), .I2(GND_net), 
            .I3(n37741), .O(n8053[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_19 (.CI(n36638), .I0(\PID_CONTROLLER.err_prev[17] ), 
            .I1(n66[17]), .CO(n36639));
    SB_CARRY add_3087_15 (.CI(n37741), .I0(n8082[12]), .I1(GND_net), .CO(n37742));
    SB_LUT4 add_3087_14_lut (.I0(GND_net), .I1(n8082[11]), .I2(GND_net), 
            .I3(n37740), .O(n8053[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[16] ), 
            .I2(n66[16]), .I3(n36637), .O(n67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_18 (.CI(n36637), .I0(\PID_CONTROLLER.err_prev[16] ), 
            .I1(n66[16]), .CO(n36638));
    SB_LUT4 add_3052_8_lut (.I0(GND_net), .I1(n1802[22]), .I2(n1703), 
            .I3(n38416), .O(n7069[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3432_5_lut (.I0(GND_net), .I1(n15854[2]), .I2(n437), .I3(n38130), 
            .O(n15644[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i499_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[7]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3087_14 (.CI(n37740), .I0(n8082[11]), .I1(GND_net), .CO(n37741));
    SB_LUT4 sub_11_add_2_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[15] ), 
            .I2(n66[15]), .I3(n36636), .O(n67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_17 (.CI(n36636), .I0(\PID_CONTROLLER.err_prev[15] ), 
            .I1(n66[15]), .CO(n36637));
    SB_LUT4 sub_11_add_2_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[14] ), 
            .I2(n66[14]), .I3(n36635), .O(n67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3052_8 (.CI(n38416), .I0(n1802[22]), .I1(n1703), .CO(n38417));
    SB_CARRY add_3432_5 (.CI(n38130), .I0(n15854[2]), .I1(n437), .CO(n38131));
    SB_LUT4 add_3087_13_lut (.I0(GND_net), .I1(n8082[10]), .I2(GND_net), 
            .I3(n37739), .O(n8053[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_13 (.CI(n37739), .I0(n8082[10]), .I1(GND_net), .CO(n37740));
    SB_CARRY sub_11_add_2_16 (.CI(n36635), .I0(\PID_CONTROLLER.err_prev[14] ), 
            .I1(n66[14]), .CO(n36636));
    SB_LUT4 add_3052_7_lut (.I0(GND_net), .I1(n1801[22]), .I2(n1699), 
            .I3(n38415), .O(n7069[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3432_4_lut (.I0(GND_net), .I1(n15854[1]), .I2(n340), .I3(n38129), 
            .O(n15644[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_12_lut (.I0(GND_net), .I1(n8082[9]), .I2(GND_net), 
            .I3(n37738), .O(n8053[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_12 (.CI(n37738), .I0(n8082[9]), .I1(GND_net), .CO(n37739));
    SB_LUT4 sub_11_add_2_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[13] ), 
            .I2(n66[13]), .I3(n36634), .O(n67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_15 (.CI(n36634), .I0(\PID_CONTROLLER.err_prev[13] ), 
            .I1(n66[13]), .CO(n36635));
    SB_LUT4 add_3087_11_lut (.I0(GND_net), .I1(n8082[8]), .I2(GND_net), 
            .I3(n37737), .O(n8053[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_11 (.CI(n37737), .I0(n8082[8]), .I1(GND_net), .CO(n37738));
    SB_CARRY add_3432_4 (.CI(n38129), .I0(n15854[1]), .I1(n340), .CO(n38130));
    SB_LUT4 add_3432_3_lut (.I0(GND_net), .I1(n15854[0]), .I2(n243), .I3(n38128), 
            .O(n15644[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_3 (.CI(n38128), .I0(n15854[0]), .I1(n243), .CO(n38129));
    SB_LUT4 add_3087_10_lut (.I0(GND_net), .I1(n8082[7]), .I2(GND_net), 
            .I3(n37736), .O(n8053[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3432_2_lut (.I0(GND_net), .I1(n53_adj_3492), .I2(n146), 
            .I3(GND_net), .O(n15644[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1047__i0 (.Q(Kd_delay_counter[0]), .C(clk32MHz), 
           .D(n57[0]));   // verilog/motorControl.v(48[27:47])
    SB_CARRY add_3087_10 (.CI(n37736), .I0(n8082[7]), .I1(GND_net), .CO(n37737));
    SB_LUT4 add_3343_16_lut (.I0(GND_net), .I1(n14438[13]), .I2(GND_net), 
            .I3(n36817), .O(n14039[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i81_2_lut (.I0(\Kd[1] ), .I1(n67[7]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3087_9_lut (.I0(GND_net), .I1(n8082[6]), .I2(GND_net), 
            .I3(n37735), .O(n8053[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_9 (.CI(n37735), .I0(n8082[6]), .I1(GND_net), .CO(n37736));
    SB_LUT4 mult_12_i18_2_lut (.I0(\Kd[0] ), .I1(n67[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_3450));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3087_8_lut (.I0(GND_net), .I1(n8082[5]), .I2(n692), .I3(n37734), 
            .O(n8053[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_8 (.CI(n37734), .I0(n8082[5]), .I1(n692), .CO(n37735));
    SB_LUT4 sub_11_add_2_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[12] ), 
            .I2(n66[12]), .I3(n36633), .O(n67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_2 (.CI(GND_net), .I0(n53_adj_3492), .I1(n146), .CO(n38128));
    SB_LUT4 add_3087_7_lut (.I0(GND_net), .I1(n8082[4]), .I2(n595_adj_3495), 
            .I3(n37733), .O(n8053[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_7 (.CI(n37733), .I0(n8082[4]), .I1(n595_adj_3495), 
            .CO(n37734));
    SB_CARRY add_3052_7 (.CI(n38415), .I0(n1801[22]), .I1(n1699), .CO(n38416));
    SB_CARRY sub_11_add_2_14 (.CI(n36633), .I0(\PID_CONTROLLER.err_prev[12] ), 
            .I1(n66[12]), .CO(n36634));
    SB_LUT4 add_3087_6_lut (.I0(GND_net), .I1(n8082[3]), .I2(n498), .I3(n37732), 
            .O(n8053[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[11] ), 
            .I2(n66[11]), .I3(n36632), .O(n67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3052_6_lut (.I0(GND_net), .I1(n1800[22]), .I2(n1695), 
            .I3(n38414), .O(n7069[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3052_6 (.CI(n38414), .I0(n1800[22]), .I1(n1695), .CO(n38415));
    SB_LUT4 add_3516_8_lut (.I0(GND_net), .I1(n16633[5]), .I2(n752), .I3(n38127), 
            .O(n16624[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_6 (.CI(n37732), .I0(n8082[3]), .I1(n498), .CO(n37733));
    SB_CARRY add_3343_16 (.CI(n36817), .I0(n14438[13]), .I1(GND_net), 
            .CO(n36818));
    SB_LUT4 add_3052_5_lut (.I0(GND_net), .I1(n1799[22]), .I2(n1691), 
            .I3(n38413), .O(n7069[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_13 (.CI(n36632), .I0(\PID_CONTROLLER.err_prev[11] ), 
            .I1(n66[11]), .CO(n36633));
    SB_LUT4 add_3516_7_lut (.I0(GND_net), .I1(n16633[4]), .I2(n658), .I3(n38126), 
            .O(n16624[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_7 (.CI(n38126), .I0(n16633[4]), .I1(n658), .CO(n38127));
    SB_LUT4 sub_11_add_2_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[10] ), 
            .I2(n66[10]), .I3(n36631), .O(n67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_5_lut (.I0(GND_net), .I1(n8082[2]), .I2(n401), .I3(n37731), 
            .O(n8053[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_15_lut (.I0(GND_net), .I1(n14438[12]), .I2(GND_net), 
            .I3(n36816), .O(n14039[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3516_6_lut (.I0(GND_net), .I1(n16633[3]), .I2(n558), .I3(n38125), 
            .O(n16624[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[8]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3087_5 (.CI(n37731), .I0(n8082[2]), .I1(n401), .CO(n37732));
    SB_LUT4 add_3087_4_lut (.I0(GND_net), .I1(n8082[1]), .I2(n304_adj_3498), 
            .I3(n37730), .O(n8053[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_4 (.CI(n37730), .I0(n8082[1]), .I1(n304_adj_3498), 
            .CO(n37731));
    SB_CARRY add_3343_15 (.CI(n36816), .I0(n14438[12]), .I1(GND_net), 
            .CO(n36817));
    SB_CARRY sub_11_add_2_12 (.CI(n36631), .I0(\PID_CONTROLLER.err_prev[10] ), 
            .I1(n66[10]), .CO(n36632));
    SB_LUT4 add_3087_3_lut (.I0(GND_net), .I1(n8082[0]), .I2(n207), .I3(n37729), 
            .O(n8053[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[9] ), 
            .I2(n66[9]), .I3(n36630), .O(n67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_6 (.CI(n38125), .I0(n16633[3]), .I1(n558), .CO(n38126));
    SB_CARRY add_3052_5 (.CI(n38413), .I0(n1799[22]), .I1(n1691), .CO(n38414));
    SB_CARRY add_3087_3 (.CI(n37729), .I0(n8082[0]), .I1(n207), .CO(n37730));
    SB_LUT4 add_3052_4_lut (.I0(GND_net), .I1(n1798[22]), .I2(n1687), 
            .I3(n38412), .O(n7069[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_2_lut (.I0(GND_net), .I1(n17_adj_3500), .I2(n110), 
            .I3(GND_net), .O(n8053[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_2 (.CI(GND_net), .I0(n17_adj_3500), .I1(n110), .CO(n37729));
    SB_CARRY add_3052_4 (.CI(n38412), .I0(n1798[22]), .I1(n1687), .CO(n38413));
    SB_LUT4 add_3516_5_lut (.I0(GND_net), .I1(n16633[2]), .I2(n464), .I3(n38124), 
            .O(n16624[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_29_lut (.I0(GND_net), .I1(n8053[26]), .I2(GND_net), 
            .I3(n37728), .O(n8023[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_5 (.CI(n38124), .I0(n16633[2]), .I1(n464), .CO(n38125));
    SB_LUT4 add_3086_28_lut (.I0(GND_net), .I1(n8053[25]), .I2(GND_net), 
            .I3(n37727), .O(n8023[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3516_4_lut (.I0(GND_net), .I1(n16633[1]), .I2(n370_adj_3471), 
            .I3(n38123), .O(n16624[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_28 (.CI(n37727), .I0(n8053[25]), .I1(GND_net), .CO(n37728));
    SB_LUT4 add_3086_27_lut (.I0(GND_net), .I1(n8053[24]), .I2(GND_net), 
            .I3(n37726), .O(n8023[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_27 (.CI(n37726), .I0(n8053[24]), .I1(GND_net), .CO(n37727));
    SB_CARRY sub_11_add_2_11 (.CI(n36630), .I0(\PID_CONTROLLER.err_prev[9] ), 
            .I1(n66[9]), .CO(n36631));
    SB_LUT4 unary_minus_17_inv_0_i32_1_lut (.I0(\deadband[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[31]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3086_26_lut (.I0(GND_net), .I1(n8053[23]), .I2(GND_net), 
            .I3(n37725), .O(n8023[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_26 (.CI(n37725), .I0(n8053[23]), .I1(GND_net), .CO(n37726));
    SB_LUT4 add_3086_25_lut (.I0(GND_net), .I1(n8053[22]), .I2(GND_net), 
            .I3(n37724), .O(n8023[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3052_3_lut (.I0(GND_net), .I1(n1797[22]), .I2(n1683), 
            .I3(n38411), .O(n7069[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_4 (.CI(n38123), .I0(n16633[1]), .I1(n370_adj_3471), 
            .CO(n38124));
    SB_CARRY add_3086_25 (.CI(n37724), .I0(n8053[22]), .I1(GND_net), .CO(n37725));
    SB_LUT4 add_3086_24_lut (.I0(GND_net), .I1(n8053[21]), .I2(GND_net), 
            .I3(n37723), .O(n8023[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_24 (.CI(n37723), .I0(n8053[21]), .I1(GND_net), .CO(n37724));
    SB_LUT4 add_3516_3_lut (.I0(GND_net), .I1(n16633[0]), .I2(n276), .I3(n38122), 
            .O(n16624[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_23_lut (.I0(GND_net), .I1(n8053[20]), .I2(GND_net), 
            .I3(n37722), .O(n8023[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_23 (.CI(n37722), .I0(n8053[20]), .I1(GND_net), .CO(n37723));
    SB_CARRY add_3052_3 (.CI(n38411), .I0(n1797[22]), .I1(n1683), .CO(n38412));
    SB_LUT4 add_3086_22_lut (.I0(GND_net), .I1(n8053[19]), .I2(GND_net), 
            .I3(n37721), .O(n8023[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_22 (.CI(n37721), .I0(n8053[19]), .I1(GND_net), .CO(n37722));
    SB_LUT4 add_3052_2_lut (.I0(GND_net), .I1(n1796[22]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n7069[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_21_lut (.I0(GND_net), .I1(n8053[18]), .I2(GND_net), 
            .I3(n37720), .O(n8023[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_21 (.CI(n37720), .I0(n8053[18]), .I1(GND_net), .CO(n37721));
    SB_CARRY add_3052_2 (.CI(GND_net), .I0(n1796[22]), .I1(\PID_CONTROLLER.integral [9]), 
            .CO(n38411));
    SB_LUT4 add_3086_20_lut (.I0(GND_net), .I1(n8053[17]), .I2(GND_net), 
            .I3(n37719), .O(n8023[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_20 (.CI(n37719), .I0(n8053[17]), .I1(GND_net), .CO(n37720));
    SB_LUT4 add_3086_19_lut (.I0(GND_net), .I1(n8053[16]), .I2(GND_net), 
            .I3(n37718), .O(n8023[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_22_lut (.I0(GND_net), .I1(n9331[19]), .I2(GND_net), 
            .I3(n38410), .O(n8476[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_19 (.CI(n37718), .I0(n8053[16]), .I1(GND_net), .CO(n37719));
    SB_LUT4 add_3086_18_lut (.I0(GND_net), .I1(n8053[15]), .I2(GND_net), 
            .I3(n37717), .O(n8023[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_21_lut (.I0(GND_net), .I1(n9331[18]), .I2(GND_net), 
            .I3(n38409), .O(n8476[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_18 (.CI(n37717), .I0(n8053[15]), .I1(GND_net), .CO(n37718));
    SB_LUT4 add_3086_17_lut (.I0(GND_net), .I1(n8053[14]), .I2(GND_net), 
            .I3(n37716), .O(n8023[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_21 (.CI(n38409), .I0(n9331[18]), .I1(GND_net), .CO(n38410));
    SB_CARRY add_3086_17 (.CI(n37716), .I0(n8053[14]), .I1(GND_net), .CO(n37717));
    SB_LUT4 add_3086_16_lut (.I0(GND_net), .I1(n8053[13]), .I2(GND_net), 
            .I3(n37715), .O(n8023[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i146_2_lut (.I0(\Kd[2] ), .I1(n67[7]), .I2(GND_net), 
            .I3(GND_net), .O(n216));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3109_20_lut (.I0(GND_net), .I1(n9331[17]), .I2(GND_net), 
            .I3(n38408), .O(n8476[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_16 (.CI(n37715), .I0(n8053[13]), .I1(GND_net), .CO(n37716));
    SB_LUT4 add_3086_15_lut (.I0(GND_net), .I1(n8053[12]), .I2(GND_net), 
            .I3(n37714), .O(n8023[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_20 (.CI(n38408), .I0(n9331[17]), .I1(GND_net), .CO(n38409));
    SB_CARRY add_3086_15 (.CI(n37714), .I0(n8053[12]), .I1(GND_net), .CO(n37715));
    SB_LUT4 add_3086_14_lut (.I0(GND_net), .I1(n8053[11]), .I2(GND_net), 
            .I3(n37713), .O(n8023[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_19_lut (.I0(GND_net), .I1(n9331[16]), .I2(GND_net), 
            .I3(n38407), .O(n8476[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_3 (.CI(n38122), .I0(n16633[0]), .I1(n276), .CO(n38123));
    SB_CARRY add_3086_14 (.CI(n37713), .I0(n8053[11]), .I1(GND_net), .CO(n37714));
    SB_LUT4 add_3343_14_lut (.I0(GND_net), .I1(n14438[11]), .I2(GND_net), 
            .I3(n36815), .O(n14039[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_14 (.CI(n36815), .I0(n14438[11]), .I1(GND_net), 
            .CO(n36816));
    SB_LUT4 add_3516_2_lut (.I0(GND_net), .I1(n86_adj_3409), .I2(n182), 
            .I3(GND_net), .O(n16624[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_13_lut (.I0(GND_net), .I1(n8053[10]), .I2(GND_net), 
            .I3(n37712), .O(n8023[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_13_lut (.I0(GND_net), .I1(n14438[10]), .I2(GND_net), 
            .I3(n36814), .O(n14039[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_13 (.CI(n36814), .I0(n14438[10]), .I1(GND_net), 
            .CO(n36815));
    SB_CARRY add_3109_19 (.CI(n38407), .I0(n9331[16]), .I1(GND_net), .CO(n38408));
    SB_CARRY add_3516_2 (.CI(GND_net), .I0(n86_adj_3409), .I1(n182), .CO(n38122));
    SB_CARRY add_3086_13 (.CI(n37712), .I0(n8053[10]), .I1(GND_net), .CO(n37713));
    SB_LUT4 add_3343_12_lut (.I0(GND_net), .I1(n14438[9]), .I2(GND_net), 
            .I3(n36813), .O(n14039[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[8] ), 
            .I2(n66[8]), .I3(n36629), .O(n67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_12 (.CI(n36813), .I0(n14438[9]), .I1(GND_net), .CO(n36814));
    SB_CARRY sub_11_add_2_10 (.CI(n36629), .I0(\PID_CONTROLLER.err_prev[8] ), 
            .I1(n66[8]), .CO(n36630));
    SB_LUT4 add_3446_15_lut (.I0(GND_net), .I1(n16035[12]), .I2(GND_net), 
            .I3(n38121), .O(n15854[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_12_lut (.I0(GND_net), .I1(n8053[9]), .I2(GND_net), 
            .I3(n37711), .O(n8023[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_18_lut (.I0(GND_net), .I1(n9331[15]), .I2(GND_net), 
            .I3(n38406), .O(n8476[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_11_lut (.I0(GND_net), .I1(n14438[8]), .I2(GND_net), 
            .I3(n36812), .O(n14039[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[7] ), 
            .I2(n66[7]), .I3(n36628), .O(n67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_11 (.CI(n36812), .I0(n14438[8]), .I1(GND_net), .CO(n36813));
    SB_CARRY sub_11_add_2_9 (.CI(n36628), .I0(\PID_CONTROLLER.err_prev[7] ), 
            .I1(n66[7]), .CO(n36629));
    SB_LUT4 add_3446_14_lut (.I0(GND_net), .I1(n16035[11]), .I2(GND_net), 
            .I3(n38120), .O(n15854[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_18 (.CI(n38406), .I0(n9331[15]), .I1(GND_net), .CO(n38407));
    SB_CARRY add_3446_14 (.CI(n38120), .I0(n16035[11]), .I1(GND_net), 
            .CO(n38121));
    SB_CARRY add_3086_12 (.CI(n37711), .I0(n8053[9]), .I1(GND_net), .CO(n37712));
    SB_LUT4 add_3343_10_lut (.I0(GND_net), .I1(n14438[7]), .I2(GND_net), 
            .I3(n36811), .O(n14039[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_10 (.CI(n36811), .I0(n14438[7]), .I1(GND_net), .CO(n36812));
    SB_LUT4 add_3446_13_lut (.I0(GND_net), .I1(n16035[10]), .I2(GND_net), 
            .I3(n38119), .O(n15854[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_11_lut (.I0(GND_net), .I1(n8053[8]), .I2(GND_net), 
            .I3(n37710), .O(n8023[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_9_lut (.I0(GND_net), .I1(n14438[6]), .I2(GND_net), 
            .I3(n36810), .O(n14039[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_9 (.CI(n36810), .I0(n14438[6]), .I1(GND_net), .CO(n36811));
    SB_LUT4 add_3109_17_lut (.I0(GND_net), .I1(n9331[14]), .I2(GND_net), 
            .I3(n38405), .O(n8476[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i206_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3086_11 (.CI(n37710), .I0(n8053[8]), .I1(GND_net), .CO(n37711));
    SB_CARRY add_3446_13 (.CI(n38119), .I0(n16035[10]), .I1(GND_net), 
            .CO(n38120));
    SB_LUT4 add_3086_10_lut (.I0(GND_net), .I1(n8053[7]), .I2(GND_net), 
            .I3(n37709), .O(n8023[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_8_lut (.I0(GND_net), .I1(n14438[5]), .I2(n713_adj_3503), 
            .I3(n36809), .O(n14039[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[6] ), 
            .I2(n66[6]), .I3(n36627), .O(n67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_10 (.CI(n37709), .I0(n8053[7]), .I1(GND_net), .CO(n37710));
    SB_CARRY add_3343_8 (.CI(n36809), .I0(n14438[5]), .I1(n713_adj_3503), 
            .CO(n36810));
    SB_CARRY sub_11_add_2_8 (.CI(n36627), .I0(\PID_CONTROLLER.err_prev[6] ), 
            .I1(n66[6]), .CO(n36628));
    SB_LUT4 add_3446_12_lut (.I0(GND_net), .I1(n16035[9]), .I2(GND_net), 
            .I3(n38118), .O(n15854[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_9_lut (.I0(GND_net), .I1(n8053[6]), .I2(GND_net), 
            .I3(n37708), .O(n8023[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_7_lut (.I0(GND_net), .I1(n14438[4]), .I2(n616_adj_3505), 
            .I3(n36808), .O(n14039[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[5] ), 
            .I2(n66[5]), .I3(n36626), .O(n67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_7 (.CI(n36808), .I0(n14438[4]), .I1(n616_adj_3505), 
            .CO(n36809));
    SB_CARRY sub_11_add_2_7 (.CI(n36626), .I0(\PID_CONTROLLER.err_prev[5] ), 
            .I1(n66[5]), .CO(n36627));
    SB_CARRY add_3109_17 (.CI(n38405), .I0(n9331[14]), .I1(GND_net), .CO(n38406));
    SB_CARRY add_3446_12 (.CI(n38118), .I0(n16035[9]), .I1(GND_net), .CO(n38119));
    SB_LUT4 add_3109_16_lut (.I0(GND_net), .I1(n9331[13]), .I2(GND_net), 
            .I3(n38404), .O(n8476[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_9 (.CI(n37708), .I0(n8053[6]), .I1(GND_net), .CO(n37709));
    SB_LUT4 add_3446_11_lut (.I0(GND_net), .I1(n16035[8]), .I2(GND_net), 
            .I3(n38117), .O(n15854[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_6_lut (.I0(GND_net), .I1(n14438[3]), .I2(n519_adj_3507), 
            .I3(n36807), .O(n14039[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_8_lut (.I0(GND_net), .I1(n8053[5]), .I2(n689), .I3(n37707), 
            .O(n8023[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[4] ), 
            .I2(n66[4]), .I3(n36625), .O(n67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_6 (.CI(n36807), .I0(n14438[3]), .I1(n519_adj_3507), 
            .CO(n36808));
    SB_CARRY sub_11_add_2_6 (.CI(n36625), .I0(\PID_CONTROLLER.err_prev[4] ), 
            .I1(n66[4]), .CO(n36626));
    SB_CARRY add_3446_11 (.CI(n38117), .I0(n16035[8]), .I1(GND_net), .CO(n38118));
    SB_LUT4 add_3446_10_lut (.I0(GND_net), .I1(n16035[7]), .I2(GND_net), 
            .I3(n38116), .O(n15854[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_8 (.CI(n37707), .I0(n8053[5]), .I1(n689), .CO(n37708));
    SB_LUT4 add_3343_5_lut (.I0(GND_net), .I1(n14438[2]), .I2(n422_adj_3509), 
            .I3(n36806), .O(n14039[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[3] ), 
            .I2(n66[3]), .I3(n36624), .O(n67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_5 (.CI(n36806), .I0(n14438[2]), .I1(n422_adj_3509), 
            .CO(n36807));
    SB_CARRY add_3109_16 (.CI(n38404), .I0(n9331[13]), .I1(GND_net), .CO(n38405));
    SB_CARRY sub_11_add_2_5 (.CI(n36624), .I0(\PID_CONTROLLER.err_prev[3] ), 
            .I1(n66[3]), .CO(n36625));
    SB_LUT4 add_3109_15_lut (.I0(GND_net), .I1(n9331[12]), .I2(GND_net), 
            .I3(n38403), .O(n8476[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_10 (.CI(n38116), .I0(n16035[7]), .I1(GND_net), .CO(n38117));
    SB_LUT4 add_3086_7_lut (.I0(GND_net), .I1(n8053[4]), .I2(n592_adj_3511), 
            .I3(n37706), .O(n8023[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_4_lut (.I0(GND_net), .I1(n14438[1]), .I2(n325_adj_3512), 
            .I3(n36805), .O(n14039[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_9_lut (.I0(GND_net), .I1(n16035[6]), .I2(GND_net), 
            .I3(n38115), .O(n15854[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[2] ), 
            .I2(n66[2]), .I3(n36623), .O(n67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_7 (.CI(n37706), .I0(n8053[4]), .I1(n592_adj_3511), 
            .CO(n37707));
    SB_CARRY sub_11_add_2_4 (.CI(n36623), .I0(\PID_CONTROLLER.err_prev[2] ), 
            .I1(n66[2]), .CO(n36624));
    SB_LUT4 add_3086_6_lut (.I0(GND_net), .I1(n8053[3]), .I2(n495), .I3(n37705), 
            .O(n8023[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_4 (.CI(n36805), .I0(n14438[1]), .I1(n325_adj_3512), 
            .CO(n36806));
    SB_LUT4 add_3343_3_lut (.I0(GND_net), .I1(n14438[0]), .I2(n228_adj_3514), 
            .I3(n36804), .O(n14039[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_9 (.CI(n38115), .I0(n16035[6]), .I1(GND_net), .CO(n38116));
    SB_LUT4 sub_11_add_2_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[1] ), 
            .I2(n66[1]), .I3(n36622), .O(n67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_3 (.CI(n36622), .I0(\PID_CONTROLLER.err_prev[1] ), 
            .I1(n66[1]), .CO(n36623));
    SB_LUT4 add_3446_8_lut (.I0(GND_net), .I1(n16035[5]), .I2(n731), .I3(n38114), 
            .O(n15854[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_6 (.CI(n37705), .I0(n8053[3]), .I1(n495), .CO(n37706));
    SB_CARRY add_3343_3 (.CI(n36804), .I0(n14438[0]), .I1(n228_adj_3514), 
            .CO(n36805));
    SB_LUT4 sub_11_add_2_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[0] ), 
            .I2(n66[0]), .I3(VCC_net), .O(n67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_2 (.CI(VCC_net), .I0(\PID_CONTROLLER.err_prev[0] ), 
            .I1(n66[0]), .CO(n36622));
    SB_LUT4 add_3343_2_lut (.I0(GND_net), .I1(n38_adj_3517), .I2(n131_adj_3518), 
            .I3(GND_net), .O(n14039[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_25_lut (.I0(n852[14]), .I1(GND_net), .I2(PHASES_5__N_3046), 
            .I3(n36621), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3109_15 (.CI(n38403), .I0(n9331[12]), .I1(GND_net), .CO(n38404));
    SB_LUT4 unary_minus_70_add_3_24_lut (.I0(n852[18]), .I1(GND_net), .I2(n73[22]), 
            .I3(n36620), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_3086_5_lut (.I0(GND_net), .I1(n8053[2]), .I2(n398), .I3(n37704), 
            .O(n8023[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_8 (.CI(n38114), .I0(n16035[5]), .I1(n731), .CO(n38115));
    SB_LUT4 add_3109_14_lut (.I0(GND_net), .I1(n9331[11]), .I2(GND_net), 
            .I3(n38402), .O(n8476[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_5 (.CI(n37704), .I0(n8053[2]), .I1(n398), .CO(n37705));
    SB_LUT4 add_3446_7_lut (.I0(GND_net), .I1(n16035[4]), .I2(n634), .I3(n38113), 
            .O(n15854[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_4_lut (.I0(GND_net), .I1(n8053[1]), .I2(n301_adj_3522), 
            .I3(n37703), .O(n8023[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_4 (.CI(n37703), .I0(n8053[1]), .I1(n301_adj_3522), 
            .CO(n37704));
    SB_CARRY add_3446_7 (.CI(n38113), .I0(n16035[4]), .I1(n634), .CO(n38114));
    SB_LUT4 add_3086_3_lut (.I0(GND_net), .I1(n8053[0]), .I2(n204), .I3(n37702), 
            .O(n8023[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_2 (.CI(GND_net), .I0(n38_adj_3517), .I1(n131_adj_3518), 
            .CO(n36804));
    SB_CARRY unary_minus_70_add_3_24 (.CI(n36620), .I0(GND_net), .I1(n73[22]), 
            .CO(n36621));
    SB_LUT4 add_3363_20_lut (.I0(GND_net), .I1(n14797[17]), .I2(GND_net), 
            .I3(n36803), .O(n14438[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_23_lut (.I0(n852[10]), .I1(GND_net), .I2(n73[21]), 
            .I3(n36619), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mult_12_i89_2_lut (.I0(\Kd[1] ), .I1(n67[11]), .I2(GND_net), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3446_6_lut (.I0(GND_net), .I1(n16035[3]), .I2(n537), .I3(n38112), 
            .O(n15854[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_3 (.CI(n37702), .I0(n8053[0]), .I1(n204), .CO(n37703));
    SB_LUT4 add_3363_19_lut (.I0(GND_net), .I1(n14797[16]), .I2(GND_net), 
            .I3(n36802), .O(n14438[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_23 (.CI(n36619), .I0(GND_net), .I1(n73[21]), 
            .CO(n36620));
    SB_CARRY add_3109_14 (.CI(n38402), .I0(n9331[11]), .I1(GND_net), .CO(n38403));
    SB_LUT4 mult_12_i26_2_lut (.I0(\Kd[0] ), .I1(n67[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_3370));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i26_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3446_6 (.CI(n38112), .I0(n16035[3]), .I1(n537), .CO(n38113));
    SB_LUT4 add_3446_5_lut (.I0(GND_net), .I1(n16035[2]), .I2(n440), .I3(n38111), 
            .O(n15854[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_2_lut (.I0(GND_net), .I1(n14_adj_3525), .I2(n107), 
            .I3(GND_net), .O(n8023[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_2 (.CI(GND_net), .I0(n14_adj_3525), .I1(n107), .CO(n37702));
    SB_LUT4 add_3085_30_lut (.I0(GND_net), .I1(n8023[27]), .I2(GND_net), 
            .I3(n37701), .O(n7992[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_19 (.CI(n36802), .I0(n14797[16]), .I1(GND_net), 
            .CO(n36803));
    SB_LUT4 unary_minus_70_add_3_22_lut (.I0(n852[16]), .I1(GND_net), .I2(n73[20]), 
            .I3(n36618), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_3109_13_lut (.I0(GND_net), .I1(n9331[10]), .I2(GND_net), 
            .I3(n38401), .O(n8476[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_5 (.CI(n38111), .I0(n16035[2]), .I1(n440), .CO(n38112));
    SB_CARRY unary_minus_70_add_3_22 (.CI(n36618), .I0(GND_net), .I1(n73[20]), 
            .CO(n36619));
    SB_LUT4 add_3085_29_lut (.I0(GND_net), .I1(n8023[26]), .I2(GND_net), 
            .I3(n37700), .O(n7992[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_18_lut (.I0(GND_net), .I1(n14797[15]), .I2(GND_net), 
            .I3(n36801), .O(n14438[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_21_lut (.I0(n852[11]), .I1(GND_net), .I2(n73[19]), 
            .I3(n36617), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3085_29 (.CI(n37700), .I0(n8023[26]), .I1(GND_net), .CO(n37701));
    SB_CARRY unary_minus_70_add_3_21 (.CI(n36617), .I0(GND_net), .I1(n73[19]), 
            .CO(n36618));
    SB_LUT4 add_3446_4_lut (.I0(GND_net), .I1(n16035[1]), .I2(n343), .I3(n38110), 
            .O(n15854[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3085_28_lut (.I0(GND_net), .I1(n8023[25]), .I2(GND_net), 
            .I3(n37699), .O(n7992[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_18 (.CI(n36801), .I0(n14797[15]), .I1(GND_net), 
            .CO(n36802));
    SB_LUT4 unary_minus_70_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n73[18]), 
            .I3(n36616), .O(n852[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_28 (.CI(n37699), .I0(n8023[25]), .I1(GND_net), .CO(n37700));
    SB_CARRY add_3446_4 (.CI(n38110), .I0(n16035[1]), .I1(n343), .CO(n38111));
    SB_LUT4 add_3085_27_lut (.I0(GND_net), .I1(n8023[24]), .I2(GND_net), 
            .I3(n37698), .O(n7992[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_3_lut (.I0(GND_net), .I1(n16035[0]), .I2(n246), .I3(n38109), 
            .O(n15854[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_20 (.CI(n36616), .I0(GND_net), .I1(n73[18]), 
            .CO(n36617));
    SB_LUT4 unary_minus_70_add_3_19_lut (.I0(n852[15]), .I1(GND_net), .I2(n73[17]), 
            .I3(n36615), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3446_3 (.CI(n38109), .I0(n16035[0]), .I1(n246), .CO(n38110));
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[9]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3085_27 (.CI(n37698), .I0(n8023[24]), .I1(GND_net), .CO(n37699));
    SB_CARRY add_3109_13 (.CI(n38401), .I0(n9331[10]), .I1(GND_net), .CO(n38402));
    SB_LUT4 add_3109_12_lut (.I0(GND_net), .I1(n9331[9]), .I2(GND_net), 
            .I3(n38400), .O(n8476[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3085_26_lut (.I0(GND_net), .I1(n8023[23]), .I2(GND_net), 
            .I3(n37697), .O(n7992[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_2_lut (.I0(GND_net), .I1(n56), .I2(n149), .I3(GND_net), 
            .O(n15854[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_19 (.CI(n36615), .I0(GND_net), .I1(n73[17]), 
            .CO(n36616));
    SB_CARRY add_3085_26 (.CI(n37697), .I0(n8023[23]), .I1(GND_net), .CO(n37698));
    SB_LUT4 add_3085_25_lut (.I0(GND_net), .I1(n8023[22]), .I2(GND_net), 
            .I3(n37696), .O(n7992[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_25 (.CI(n37696), .I0(n8023[22]), .I1(GND_net), .CO(n37697));
    SB_LUT4 add_3363_17_lut (.I0(GND_net), .I1(n14797[14]), .I2(GND_net), 
            .I3(n36800), .O(n14438[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i87_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n128_adj_3446));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i87_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3363_17 (.CI(n36800), .I0(n14797[14]), .I1(GND_net), 
            .CO(n36801));
    SB_CARRY add_3109_12 (.CI(n38400), .I0(n9331[9]), .I1(GND_net), .CO(n38401));
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3445));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[0]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3085_24_lut (.I0(GND_net), .I1(n8023[21]), .I2(GND_net), 
            .I3(n37695), .O(n7992[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_2 (.CI(GND_net), .I0(n56), .I1(n149), .CO(n38109));
    SB_LUT4 add_3459_14_lut (.I0(GND_net), .I1(n16189[11]), .I2(GND_net), 
            .I3(n38108), .O(n16035[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_24 (.CI(n37695), .I0(n8023[21]), .I1(GND_net), .CO(n37696));
    SB_LUT4 add_3459_13_lut (.I0(GND_net), .I1(n16189[10]), .I2(GND_net), 
            .I3(n38107), .O(n16035[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3085_23_lut (.I0(GND_net), .I1(n8023[20]), .I2(GND_net), 
            .I3(n37694), .O(n7992[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_16_lut (.I0(GND_net), .I1(n14797[13]), .I2(GND_net), 
            .I3(n36799), .O(n14438[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_16 (.CI(n36799), .I0(n14797[13]), .I1(GND_net), 
            .CO(n36800));
    SB_LUT4 add_3109_11_lut (.I0(GND_net), .I1(n9331[8]), .I2(GND_net), 
            .I3(n38399), .O(n8476[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_13 (.CI(n38107), .I0(n16189[10]), .I1(GND_net), 
            .CO(n38108));
    SB_CARRY add_3085_23 (.CI(n37694), .I0(n8023[20]), .I1(GND_net), .CO(n37695));
    SB_LUT4 add_3459_12_lut (.I0(GND_net), .I1(n16189[9]), .I2(GND_net), 
            .I3(n38106), .O(n16035[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_11 (.CI(n38399), .I0(n9331[8]), .I1(GND_net), .CO(n38400));
    SB_LUT4 add_3085_22_lut (.I0(GND_net), .I1(n8023[19]), .I2(GND_net), 
            .I3(n37693), .O(n7992[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_22 (.CI(n37693), .I0(n8023[19]), .I1(GND_net), .CO(n37694));
    SB_LUT4 add_3085_21_lut (.I0(GND_net), .I1(n8023[18]), .I2(GND_net), 
            .I3(n37692), .O(n7992[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_15_lut (.I0(GND_net), .I1(n14797[12]), .I2(GND_net), 
            .I3(n36798), .O(n14438[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_21 (.CI(n37692), .I0(n8023[18]), .I1(GND_net), .CO(n37693));
    SB_LUT4 add_3085_20_lut (.I0(GND_net), .I1(n8023[17]), .I2(GND_net), 
            .I3(n37691), .O(n7992[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_10_lut (.I0(GND_net), .I1(n9331[7]), .I2(GND_net), 
            .I3(n38398), .O(n8476[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_12 (.CI(n38106), .I0(n16189[9]), .I1(GND_net), .CO(n38107));
    SB_CARRY add_3085_20 (.CI(n37691), .I0(n8023[17]), .I1(GND_net), .CO(n37692));
    SB_CARRY add_3109_10 (.CI(n38398), .I0(n9331[7]), .I1(GND_net), .CO(n38399));
    SB_LUT4 add_3085_19_lut (.I0(GND_net), .I1(n8023[16]), .I2(GND_net), 
            .I3(n37690), .O(n7992[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3459_11_lut (.I0(GND_net), .I1(n16189[8]), .I2(GND_net), 
            .I3(n38105), .O(n16035[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_19 (.CI(n37690), .I0(n8023[16]), .I1(GND_net), .CO(n37691));
    SB_CARRY add_3363_15 (.CI(n36798), .I0(n14797[12]), .I1(GND_net), 
            .CO(n36799));
    SB_LUT4 unary_minus_70_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n73[16]), 
            .I3(n36614), .O(n852[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_9_lut (.I0(GND_net), .I1(n9331[6]), .I2(GND_net), 
            .I3(n38397), .O(n8476[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_11 (.CI(n38105), .I0(n16189[8]), .I1(GND_net), .CO(n38106));
    SB_LUT4 add_3085_18_lut (.I0(GND_net), .I1(n8023[15]), .I2(GND_net), 
            .I3(n37689), .O(n7992[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3459_10_lut (.I0(GND_net), .I1(n16189[7]), .I2(GND_net), 
            .I3(n38104), .O(n16035[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_18 (.CI(n37689), .I0(n8023[15]), .I1(GND_net), .CO(n37690));
    SB_LUT4 add_3363_14_lut (.I0(GND_net), .I1(n14797[11]), .I2(GND_net), 
            .I3(n36797), .O(n14438[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_18 (.CI(n36614), .I0(GND_net), .I1(n73[16]), 
            .CO(n36615));
    SB_LUT4 add_3085_17_lut (.I0(GND_net), .I1(n8023[14]), .I2(GND_net), 
            .I3(n37688), .O(n7992[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_count_1048__i0 (.Q(pwm_count[0]), .C(clk32MHz), .D(n75[0]));   // verilog/motorControl.v(99[18:29])
    SB_CARRY add_3459_10 (.CI(n38104), .I0(n16189[7]), .I1(GND_net), .CO(n38105));
    SB_LUT4 add_3459_9_lut (.I0(GND_net), .I1(n16189[6]), .I2(GND_net), 
            .I3(n38103), .O(n16035[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n73[15]), 
            .I3(n36613), .O(n852[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_9 (.CI(n38397), .I0(n9331[6]), .I1(GND_net), .CO(n38398));
    SB_CARRY add_3459_9 (.CI(n38103), .I0(n16189[6]), .I1(GND_net), .CO(n38104));
    SB_LUT4 add_3459_8_lut (.I0(GND_net), .I1(n16189[5]), .I2(n734), .I3(n38102), 
            .O(n16035[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[10]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3085_17 (.CI(n37688), .I0(n8023[14]), .I1(GND_net), .CO(n37689));
    SB_LUT4 add_3085_16_lut (.I0(GND_net), .I1(n8023[13]), .I2(GND_net), 
            .I3(n37687), .O(n7992[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_8_lut (.I0(GND_net), .I1(n9331[5]), .I2(n545), .I3(n38396), 
            .O(n8476[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_8 (.CI(n38102), .I0(n16189[5]), .I1(n734), .CO(n38103));
    SB_CARRY add_3085_16 (.CI(n37687), .I0(n8023[13]), .I1(GND_net), .CO(n37688));
    SB_CARRY add_3363_14 (.CI(n36797), .I0(n14797[11]), .I1(GND_net), 
            .CO(n36798));
    SB_CARRY add_3109_8 (.CI(n38396), .I0(n9331[5]), .I1(n545), .CO(n38397));
    SB_LUT4 add_3459_7_lut (.I0(GND_net), .I1(n16189[4]), .I2(n637), .I3(n38101), 
            .O(n16035[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3085_15_lut (.I0(GND_net), .I1(n8023[12]), .I2(GND_net), 
            .I3(n37686), .O(n7992[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_7 (.CI(n38101), .I0(n16189[4]), .I1(n637), .CO(n38102));
    SB_CARRY add_3085_15 (.CI(n37686), .I0(n8023[12]), .I1(GND_net), .CO(n37687));
    SB_LUT4 add_3363_13_lut (.I0(GND_net), .I1(n14797[10]), .I2(GND_net), 
            .I3(n36796), .O(n14438[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_13 (.CI(n36796), .I0(n14797[10]), .I1(GND_net), 
            .CO(n36797));
    SB_LUT4 add_3459_6_lut (.I0(GND_net), .I1(n16189[3]), .I2(n540), .I3(n38100), 
            .O(n16035[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3085_14_lut (.I0(GND_net), .I1(n8023[11]), .I2(GND_net), 
            .I3(n37685), .O(n7992[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_7_lut (.I0(GND_net), .I1(n9331[4]), .I2(n472), .I3(n38395), 
            .O(n8476[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_14 (.CI(n37685), .I0(n8023[11]), .I1(GND_net), .CO(n37686));
    SB_CARRY add_3459_6 (.CI(n38100), .I0(n16189[3]), .I1(n540), .CO(n38101));
    SB_LUT4 add_3363_12_lut (.I0(GND_net), .I1(n14797[9]), .I2(GND_net), 
            .I3(n36795), .O(n14438[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3085_13_lut (.I0(GND_net), .I1(n8023[10]), .I2(GND_net), 
            .I3(n37684), .O(n7992[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_13 (.CI(n37684), .I0(n8023[10]), .I1(GND_net), .CO(n37685));
    SB_LUT4 add_3085_12_lut (.I0(GND_net), .I1(n8023[9]), .I2(GND_net), 
            .I3(n37683), .O(n7992[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_17 (.CI(n36613), .I0(GND_net), .I1(n73[15]), 
            .CO(n36614));
    SB_LUT4 add_3459_5_lut (.I0(GND_net), .I1(n16189[2]), .I2(n443_adj_3536), 
            .I3(n38099), .O(n16035[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n73[14]), 
            .I3(n36612), .O(n852[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_12 (.CI(n37683), .I0(n8023[9]), .I1(GND_net), .CO(n37684));
    SB_CARRY add_3363_12 (.CI(n36795), .I0(n14797[9]), .I1(GND_net), .CO(n36796));
    SB_CARRY unary_minus_70_add_3_16 (.CI(n36612), .I0(GND_net), .I1(n73[14]), 
            .CO(n36613));
    SB_CARRY add_3109_7 (.CI(n38395), .I0(n9331[4]), .I1(n472), .CO(n38396));
    SB_CARRY add_3459_5 (.CI(n38099), .I0(n16189[2]), .I1(n443_adj_3536), 
            .CO(n38100));
    SB_LUT4 add_3085_11_lut (.I0(GND_net), .I1(n8023[8]), .I2(GND_net), 
            .I3(n37682), .O(n7992[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3459_4_lut (.I0(GND_net), .I1(n16189[1]), .I2(n346), .I3(n38098), 
            .O(n16035[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_11 (.CI(n37682), .I0(n8023[8]), .I1(GND_net), .CO(n37683));
    SB_LUT4 add_3363_11_lut (.I0(GND_net), .I1(n14797[8]), .I2(GND_net), 
            .I3(n36794), .O(n14438[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_15_lut (.I0(n48196), .I1(GND_net), .I2(n73[13]), 
            .I3(n36611), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY unary_minus_70_add_3_15 (.CI(n36611), .I0(GND_net), .I1(n73[13]), 
            .CO(n36612));
    SB_LUT4 add_3109_6_lut (.I0(GND_net), .I1(n9331[3]), .I2(n399), .I3(n38394), 
            .O(n8476[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_4 (.CI(n38098), .I0(n16189[1]), .I1(n346), .CO(n38099));
    SB_LUT4 add_3085_10_lut (.I0(GND_net), .I1(n8023[7]), .I2(GND_net), 
            .I3(n37681), .O(n7992[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_32_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n6546[29]), 
            .I2(GND_net), .I3(n37192), .O(n5790[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_2137_31_lut (.I0(GND_net), .I1(n6546[28]), .I2(GND_net), 
            .I3(n37191), .O(n76[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_11 (.CI(n36794), .I0(n14797[8]), .I1(GND_net), .CO(n36795));
    SB_LUT4 add_3459_3_lut (.I0(GND_net), .I1(n16189[0]), .I2(n249), .I3(n38097), 
            .O(n16035[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_10 (.CI(n37681), .I0(n8023[7]), .I1(GND_net), .CO(n37682));
    SB_CARRY mult_10_add_2137_31 (.CI(n37191), .I0(n6546[28]), .I1(GND_net), 
            .CO(n37192));
    SB_LUT4 add_3363_10_lut (.I0(GND_net), .I1(n14797[7]), .I2(GND_net), 
            .I3(n36793), .O(n14438[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3085_9_lut (.I0(GND_net), .I1(n8023[6]), .I2(GND_net), 
            .I3(n37680), .O(n7992[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_9 (.CI(n37680), .I0(n8023[6]), .I1(GND_net), .CO(n37681));
    SB_LUT4 mult_10_add_2137_30_lut (.I0(GND_net), .I1(n6546[27]), .I2(GND_net), 
            .I3(n37190), .O(n76[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_30 (.CI(n37190), .I0(n6546[27]), .I1(GND_net), 
            .CO(n37191));
    SB_CARRY add_3459_3 (.CI(n38097), .I0(n16189[0]), .I1(n249), .CO(n38098));
    SB_LUT4 add_3085_8_lut (.I0(GND_net), .I1(n8023[5]), .I2(n686), .I3(n37679), 
            .O(n7992[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_29_lut (.I0(GND_net), .I1(n6546[26]), .I2(GND_net), 
            .I3(n37189), .O(n76[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_10 (.CI(n36793), .I0(n14797[7]), .I1(GND_net), .CO(n36794));
    SB_CARRY mult_10_add_2137_29 (.CI(n37189), .I0(n6546[26]), .I1(GND_net), 
            .CO(n37190));
    SB_LUT4 add_3363_9_lut (.I0(GND_net), .I1(n14797[6]), .I2(GND_net), 
            .I3(n36792), .O(n14438[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_6 (.CI(n38394), .I0(n9331[3]), .I1(n399), .CO(n38395));
    SB_LUT4 add_3459_2_lut (.I0(GND_net), .I1(n59), .I2(n152), .I3(GND_net), 
            .O(n16035[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_8 (.CI(n37679), .I0(n8023[5]), .I1(n686), .CO(n37680));
    SB_LUT4 mult_10_add_2137_28_lut (.I0(GND_net), .I1(n6546[25]), .I2(GND_net), 
            .I3(n37188), .O(n76[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_28 (.CI(n37188), .I0(n6546[25]), .I1(GND_net), 
            .CO(n37189));
    SB_CARRY add_3459_2 (.CI(GND_net), .I0(n59), .I1(n152), .CO(n38097));
    SB_LUT4 add_3085_7_lut (.I0(GND_net), .I1(n8023[4]), .I2(n589_adj_3541), 
            .I3(n37678), .O(n7992[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_27_lut (.I0(GND_net), .I1(n6546[24]), .I2(GND_net), 
            .I3(n37187), .O(n76[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_7 (.CI(n37678), .I0(n8023[4]), .I1(n589_adj_3541), 
            .CO(n37679));
    SB_CARRY add_3363_9 (.CI(n36792), .I0(n14797[6]), .I1(GND_net), .CO(n36793));
    SB_LUT4 add_3471_13_lut (.I0(GND_net), .I1(n16318[10]), .I2(GND_net), 
            .I3(n38096), .O(n16189[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_27 (.CI(n37187), .I0(n6546[24]), .I1(GND_net), 
            .CO(n37188));
    SB_LUT4 add_3085_6_lut (.I0(GND_net), .I1(n8023[3]), .I2(n492), .I3(n37677), 
            .O(n7992[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_8_lut (.I0(GND_net), .I1(n14797[5]), .I2(n716), .I3(n36791), 
            .O(n14438[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_5_lut (.I0(GND_net), .I1(n9331[2]), .I2(n326), .I3(n38393), 
            .O(n8476[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_26_lut (.I0(GND_net), .I1(n6546[23]), .I2(GND_net), 
            .I3(n37186), .O(n76[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_5 (.CI(n38393), .I0(n9331[2]), .I1(n326), .CO(n38394));
    SB_LUT4 add_3471_12_lut (.I0(GND_net), .I1(n16318[9]), .I2(GND_net), 
            .I3(n38095), .O(n16189[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_14_lut (.I0(n852[9]), .I1(GND_net), .I2(n73[12]), 
            .I3(n36610), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3471_12 (.CI(n38095), .I0(n16318[9]), .I1(GND_net), .CO(n38096));
    SB_CARRY add_3085_6 (.CI(n37677), .I0(n8023[3]), .I1(n492), .CO(n37678));
    SB_CARRY mult_10_add_2137_26 (.CI(n37186), .I0(n6546[23]), .I1(GND_net), 
            .CO(n37187));
    SB_LUT4 add_3085_5_lut (.I0(GND_net), .I1(n8023[2]), .I2(n395), .I3(n37676), 
            .O(n7992[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_8 (.CI(n36791), .I0(n14797[5]), .I1(n716), .CO(n36792));
    SB_CARRY add_3085_5 (.CI(n37676), .I0(n8023[2]), .I1(n395), .CO(n37677));
    SB_LUT4 mult_10_add_2137_25_lut (.I0(GND_net), .I1(n6546[22]), .I2(GND_net), 
            .I3(n37185), .O(n76[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_7_lut (.I0(GND_net), .I1(n14797[4]), .I2(n619), .I3(n36790), 
            .O(n14438[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_25 (.CI(n37185), .I0(n6546[22]), .I1(GND_net), 
            .CO(n37186));
    SB_LUT4 add_3471_11_lut (.I0(GND_net), .I1(n16318[8]), .I2(GND_net), 
            .I3(n38094), .O(n16189[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i211_2_lut (.I0(\Kd[3] ), .I1(n67[7]), .I2(GND_net), 
            .I3(GND_net), .O(n313));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3085_4_lut (.I0(GND_net), .I1(n8023[1]), .I2(n298_adj_3545), 
            .I3(n37675), .O(n7992[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_24_lut (.I0(GND_net), .I1(n6546[21]), .I2(GND_net), 
            .I3(n37184), .O(n76[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_7 (.CI(n36790), .I0(n14797[4]), .I1(n619), .CO(n36791));
    SB_CARRY mult_10_add_2137_24 (.CI(n37184), .I0(n6546[21]), .I1(GND_net), 
            .CO(n37185));
    SB_LUT4 add_3363_6_lut (.I0(GND_net), .I1(n14797[3]), .I2(n522_adj_3547), 
            .I3(n36789), .O(n14438[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_14 (.CI(n36610), .I0(GND_net), .I1(n73[12]), 
            .CO(n36611));
    SB_LUT4 add_3109_4_lut (.I0(GND_net), .I1(n9331[1]), .I2(n253), .I3(n38392), 
            .O(n8476[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_11 (.CI(n38094), .I0(n16318[8]), .I1(GND_net), .CO(n38095));
    SB_CARRY add_3085_4 (.CI(n37675), .I0(n8023[1]), .I1(n298_adj_3545), 
            .CO(n37676));
    SB_LUT4 add_3085_3_lut (.I0(GND_net), .I1(n8023[0]), .I2(n201), .I3(n37674), 
            .O(n7992[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_23_lut (.I0(GND_net), .I1(n6546[20]), .I2(GND_net), 
            .I3(n37183), .O(n76[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_23 (.CI(n37183), .I0(n6546[20]), .I1(GND_net), 
            .CO(n37184));
    SB_LUT4 mult_10_add_2137_22_lut (.I0(GND_net), .I1(n6546[19]), .I2(GND_net), 
            .I3(n37182), .O(n76[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_22 (.CI(n37182), .I0(n6546[19]), .I1(GND_net), 
            .CO(n37183));
    SB_CARRY add_3085_3 (.CI(n37674), .I0(n8023[0]), .I1(n201), .CO(n37675));
    SB_LUT4 add_3085_2_lut (.I0(GND_net), .I1(n11_adj_3548), .I2(n104), 
            .I3(GND_net), .O(n7992[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_10_lut (.I0(GND_net), .I1(n16318[7]), .I2(GND_net), 
            .I3(n38093), .O(n16189[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_21_lut (.I0(GND_net), .I1(n6546[18]), .I2(GND_net), 
            .I3(n37181), .O(n76[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_21 (.CI(n37181), .I0(n6546[18]), .I1(GND_net), 
            .CO(n37182));
    SB_CARRY add_3085_2 (.CI(GND_net), .I0(n11_adj_3548), .I1(n104), .CO(n37674));
    SB_LUT4 mult_10_add_2137_20_lut (.I0(GND_net), .I1(n6546[17]), .I2(GND_net), 
            .I3(n37180), .O(n76[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i152_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n225_adj_3442));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i152_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_2137_20 (.CI(n37180), .I0(n6546[17]), .I1(GND_net), 
            .CO(n37181));
    SB_LUT4 mult_10_add_2137_19_lut (.I0(GND_net), .I1(n6546[16]), .I2(GND_net), 
            .I3(n37179), .O(n76[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_6 (.CI(n36789), .I0(n14797[3]), .I1(n522_adj_3547), 
            .CO(n36790));
    SB_CARRY mult_10_add_2137_19 (.CI(n37179), .I0(n6546[16]), .I1(GND_net), 
            .CO(n37180));
    SB_LUT4 add_3363_5_lut (.I0(GND_net), .I1(n14797[2]), .I2(n425_adj_3549), 
            .I3(n36788), .O(n14438[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n73[11]), 
            .I3(n36609), .O(n852[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_4 (.CI(n38392), .I0(n9331[1]), .I1(n253), .CO(n38393));
    SB_CARRY add_3471_10 (.CI(n38093), .I0(n16318[7]), .I1(GND_net), .CO(n38094));
    SB_LUT4 mult_12_add_2137_32_lut (.I0(n67[25]), .I1(n7960[29]), .I2(GND_net), 
            .I3(n37673), .O(n7065[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_2137_18_lut (.I0(GND_net), .I1(n6546[15]), .I2(GND_net), 
            .I3(n37178), .O(n76[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_18 (.CI(n37178), .I0(n6546[15]), .I1(GND_net), 
            .CO(n37179));
    SB_LUT4 add_3471_9_lut (.I0(GND_net), .I1(n16318[6]), .I2(GND_net), 
            .I3(n38092), .O(n16189[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_31_lut (.I0(GND_net), .I1(n7960[28]), .I2(GND_net), 
            .I3(n37672), .O(n191[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_9 (.CI(n38092), .I0(n16318[6]), .I1(GND_net), .CO(n38093));
    SB_LUT4 mult_10_add_2137_17_lut (.I0(GND_net), .I1(n6546[14]), .I2(GND_net), 
            .I3(n37177), .O(n76[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_17 (.CI(n37177), .I0(n6546[14]), .I1(GND_net), 
            .CO(n37178));
    SB_CARRY add_3363_5 (.CI(n36788), .I0(n14797[2]), .I1(n425_adj_3549), 
            .CO(n36789));
    SB_LUT4 add_3471_8_lut (.I0(GND_net), .I1(n16318[5]), .I2(n737), .I3(n38091), 
            .O(n16189[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_3_lut (.I0(GND_net), .I1(n9331[0]), .I2(n180_adj_3552), 
            .I3(n38391), .O(n8476[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_16_lut (.I0(GND_net), .I1(n6546[13]), .I2(GND_net), 
            .I3(n37176), .O(n76[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[11]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_12_add_2137_31 (.CI(n37672), .I0(n7960[28]), .I1(GND_net), 
            .CO(n37673));
    SB_CARRY mult_10_add_2137_16 (.CI(n37176), .I0(n6546[13]), .I1(GND_net), 
            .CO(n37177));
    SB_LUT4 mult_12_add_2137_30_lut (.I0(GND_net), .I1(n7960[27]), .I2(GND_net), 
            .I3(n37671), .O(n191[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_4_lut (.I0(GND_net), .I1(n14797[1]), .I2(n328_adj_3553), 
            .I3(n36787), .O(n14438[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_15_lut (.I0(GND_net), .I1(n6546[12]), .I2(GND_net), 
            .I3(n37175), .O(n76[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_3 (.CI(n38391), .I0(n9331[0]), .I1(n180_adj_3552), 
            .CO(n38392));
    SB_CARRY add_3471_8 (.CI(n38091), .I0(n16318[5]), .I1(n737), .CO(n38092));
    SB_LUT4 add_3471_7_lut (.I0(GND_net), .I1(n16318[4]), .I2(n640), .I3(n38090), 
            .O(n16189[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_30 (.CI(n37671), .I0(n7960[27]), .I1(GND_net), 
            .CO(n37672));
    SB_CARRY mult_10_add_2137_15 (.CI(n37175), .I0(n6546[12]), .I1(GND_net), 
            .CO(n37176));
    SB_LUT4 mult_10_add_2137_14_lut (.I0(GND_net), .I1(n6546[11]), .I2(GND_net), 
            .I3(n37174), .O(n76[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_7 (.CI(n38090), .I0(n16318[4]), .I1(n640), .CO(n38091));
    SB_LUT4 mult_12_add_2137_29_lut (.I0(GND_net), .I1(n7960[26]), .I2(GND_net), 
            .I3(n37670), .O(n191[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_14 (.CI(n37174), .I0(n6546[11]), .I1(GND_net), 
            .CO(n37175));
    SB_CARRY add_3363_4 (.CI(n36787), .I0(n14797[1]), .I1(n328_adj_3553), 
            .CO(n36788));
    SB_LUT4 add_3109_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n8476[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_13_lut (.I0(GND_net), .I1(n6546[10]), .I2(GND_net), 
            .I3(n37173), .O(n76[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_3_lut (.I0(GND_net), .I1(n14797[0]), .I2(n231_adj_3558), 
            .I3(n36786), .O(n14438[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_6_lut (.I0(GND_net), .I1(n16318[3]), .I2(n543), .I3(n38089), 
            .O(n16189[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_6 (.CI(n38089), .I0(n16318[3]), .I1(n543), .CO(n38090));
    SB_CARRY add_3109_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n38391));
    SB_CARRY mult_10_add_2137_13 (.CI(n37173), .I0(n6546[10]), .I1(GND_net), 
            .CO(n37174));
    SB_CARRY unary_minus_70_add_3_13 (.CI(n36609), .I0(GND_net), .I1(n73[11]), 
            .CO(n36610));
    SB_LUT4 add_3471_5_lut (.I0(GND_net), .I1(n16318[2]), .I2(n446_adj_3559), 
            .I3(n38088), .O(n16189[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_5 (.CI(n38088), .I0(n16318[2]), .I1(n446_adj_3559), 
            .CO(n38089));
    SB_CARRY mult_12_add_2137_29 (.CI(n37670), .I0(n7960[26]), .I1(GND_net), 
            .CO(n37671));
    SB_LUT4 mult_10_add_2137_12_lut (.I0(GND_net), .I1(n6546[9]), .I2(GND_net), 
            .I3(n37172), .O(n76[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_28_lut (.I0(GND_net), .I1(n7960[25]), .I2(GND_net), 
            .I3(n37669), .O(n191[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_4_lut (.I0(GND_net), .I1(n16318[1]), .I2(n349), .I3(n38087), 
            .O(n16189[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_12 (.CI(n37172), .I0(n6546[9]), .I1(GND_net), 
            .CO(n37173));
    SB_CARRY add_3471_4 (.CI(n38087), .I0(n16318[1]), .I1(n349), .CO(n38088));
    SB_CARRY mult_12_add_2137_28 (.CI(n37669), .I0(n7960[25]), .I1(GND_net), 
            .CO(n37670));
    SB_LUT4 mult_10_add_2137_11_lut (.I0(GND_net), .I1(n6546[8]), .I2(GND_net), 
            .I3(n37171), .O(n76[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_3 (.CI(n36786), .I0(n14797[0]), .I1(n231_adj_3558), 
            .CO(n36787));
    SB_CARRY mult_10_add_2137_11 (.CI(n37171), .I0(n6546[8]), .I1(GND_net), 
            .CO(n37172));
    SB_LUT4 add_3363_2_lut (.I0(GND_net), .I1(n41_adj_3563), .I2(n134_adj_3564), 
            .I3(GND_net), .O(n14438[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n73[10]), 
            .I3(n36608), .O(n852[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_10_lut (.I0(GND_net), .I1(n6546[7]), .I2(GND_net), 
            .I3(n37170), .O(n76[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_24_lut (.I0(GND_net), .I1(n8452[21]), .I2(GND_net), 
            .I3(n38390), .O(n1804[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_23_lut (.I0(GND_net), .I1(n8452[20]), .I2(GND_net), 
            .I3(n38389), .O(n1804[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_3_lut (.I0(GND_net), .I1(n16318[0]), .I2(n252), .I3(n38086), 
            .O(n16189[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_10 (.CI(n37170), .I0(n6546[7]), .I1(GND_net), 
            .CO(n37171));
    SB_CARRY add_3471_3 (.CI(n38086), .I0(n16318[0]), .I1(n252), .CO(n38087));
    SB_LUT4 mult_12_add_2137_27_lut (.I0(GND_net), .I1(n7960[24]), .I2(GND_net), 
            .I3(n37668), .O(n191[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_23 (.CI(n38389), .I0(n8452[20]), .I1(GND_net), 
            .CO(n38390));
    SB_CARRY mult_12_add_2137_27 (.CI(n37668), .I0(n7960[24]), .I1(GND_net), 
            .CO(n37669));
    SB_LUT4 mult_10_add_2137_9_lut (.I0(GND_net), .I1(n6546[6]), .I2(GND_net), 
            .I3(n37169), .O(n76[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_2_lut (.I0(GND_net), .I1(n62), .I2(n155), .I3(GND_net), 
            .O(n16189[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i276_2_lut (.I0(\Kd[4] ), .I1(n67[7]), .I2(GND_net), 
            .I3(GND_net), .O(n410));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[1]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_2137_9 (.CI(n37169), .I0(n6546[6]), .I1(GND_net), 
            .CO(n37170));
    SB_LUT4 mult_12_add_2137_26_lut (.I0(GND_net), .I1(n7960[23]), .I2(GND_net), 
            .I3(n37667), .O(n191[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_2 (.CI(GND_net), .I0(n62), .I1(n155), .CO(n38086));
    SB_LUT4 add_3108_23_lut (.I0(GND_net), .I1(n8476[20]), .I2(GND_net), 
            .I3(n38085), .O(n8452[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_26 (.CI(n37667), .I0(n7960[23]), .I1(GND_net), 
            .CO(n37668));
    SB_LUT4 mult_10_add_2137_8_lut (.I0(GND_net), .I1(n6546[5]), .I2(n680), 
            .I3(n37168), .O(n76[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_2 (.CI(GND_net), .I0(n41_adj_3563), .I1(n134_adj_3564), 
            .CO(n36786));
    SB_CARRY mult_10_add_2137_8 (.CI(n37168), .I0(n6546[5]), .I1(n680), 
            .CO(n37169));
    SB_LUT4 add_3501_10_lut (.I0(GND_net), .I1(n16575[7]), .I2(GND_net), 
            .I3(n36785), .O(n16509[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_12 (.CI(n36608), .I0(GND_net), .I1(n73[10]), 
            .CO(n36609));
    SB_LUT4 mult_10_add_2137_7_lut (.I0(GND_net), .I1(n6546[4]), .I2(n583), 
            .I3(n37167), .O(n76[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_25_lut (.I0(GND_net), .I1(n7960[22]), .I2(GND_net), 
            .I3(n37666), .O(n191[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_7 (.CI(n37167), .I0(n6546[4]), .I1(n583), 
            .CO(n37168));
    SB_LUT4 mult_10_i217_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n322_adj_3436));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1219_22_lut (.I0(GND_net), .I1(n8452[19]), .I2(GND_net), 
            .I3(n38388), .O(n1804[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_22_lut (.I0(GND_net), .I1(n8476[19]), .I2(GND_net), 
            .I3(n38084), .O(n8452[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_6_lut (.I0(GND_net), .I1(n6546[3]), .I2(n486), 
            .I3(n37166), .O(n76[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_25 (.CI(n37666), .I0(n7960[22]), .I1(GND_net), 
            .CO(n37667));
    SB_CARRY mult_10_add_2137_6 (.CI(n37166), .I0(n6546[3]), .I1(n486), 
            .CO(n37167));
    SB_LUT4 mult_10_add_2137_5_lut (.I0(GND_net), .I1(n6546[2]), .I2(n389), 
            .I3(n37165), .O(n76[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_22 (.CI(n38084), .I0(n8476[19]), .I1(GND_net), .CO(n38085));
    SB_LUT4 mult_12_add_2137_24_lut (.I0(GND_net), .I1(n7960[21]), .I2(GND_net), 
            .I3(n37665), .O(n191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_5 (.CI(n37165), .I0(n6546[2]), .I1(n389), 
            .CO(n37166));
    SB_LUT4 add_3108_21_lut (.I0(GND_net), .I1(n8476[18]), .I2(GND_net), 
            .I3(n38083), .O(n8452[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_4_lut (.I0(GND_net), .I1(n6546[1]), .I2(n292), 
            .I3(n37164), .O(n76[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3501_9_lut (.I0(GND_net), .I1(n16575[6]), .I2(GND_net), 
            .I3(n36784), .O(n16509[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[2]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[12]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3108_21 (.CI(n38083), .I0(n8476[18]), .I1(GND_net), .CO(n38084));
    SB_CARRY mult_10_add_2137_4 (.CI(n37164), .I0(n6546[1]), .I1(n292), 
            .CO(n37165));
    SB_CARRY add_3501_9 (.CI(n36784), .I0(n16575[6]), .I1(GND_net), .CO(n36785));
    SB_CARRY mult_14_add_1219_22 (.CI(n38388), .I0(n8452[19]), .I1(GND_net), 
            .CO(n38389));
    SB_LUT4 add_3108_20_lut (.I0(GND_net), .I1(n8476[17]), .I2(GND_net), 
            .I3(n38082), .O(n8452[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_24 (.CI(n37665), .I0(n7960[21]), .I1(GND_net), 
            .CO(n37666));
    SB_LUT4 mult_10_add_2137_3_lut (.I0(GND_net), .I1(n6546[0]), .I2(n195), 
            .I3(n37163), .O(n76[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_3 (.CI(n37163), .I0(n6546[0]), .I1(n195), 
            .CO(n37164));
    SB_CARRY add_3108_20 (.CI(n38082), .I0(n8476[17]), .I1(GND_net), .CO(n38083));
    SB_LUT4 mult_12_add_2137_23_lut (.I0(GND_net), .I1(n7960[20]), .I2(GND_net), 
            .I3(n37664), .O(n191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_2_lut (.I0(GND_net), .I1(n5_adj_3578), .I2(n98), 
            .I3(GND_net), .O(n76[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_19_lut (.I0(GND_net), .I1(n8476[16]), .I2(GND_net), 
            .I3(n38081), .O(n8452[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_23 (.CI(n37664), .I0(n7960[20]), .I1(GND_net), 
            .CO(n37665));
    SB_CARRY mult_10_add_2137_2 (.CI(GND_net), .I0(n5_adj_3578), .I1(n98), 
            .CO(n37163));
    SB_LUT4 add_3501_8_lut (.I0(GND_net), .I1(n16575[5]), .I2(n746), .I3(n36783), 
            .O(n16509[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3501_8 (.CI(n36783), .I0(n16575[5]), .I1(n746), .CO(n36784));
    SB_LUT4 mult_14_add_1219_21_lut (.I0(GND_net), .I1(n8452[18]), .I2(GND_net), 
            .I3(n38387), .O(n1804[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_19 (.CI(n38081), .I0(n8476[16]), .I1(GND_net), .CO(n38082));
    SB_LUT4 mult_12_add_2137_22_lut (.I0(GND_net), .I1(n7960[19]), .I2(GND_net), 
            .I3(n37663), .O(n191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_18_lut (.I0(GND_net), .I1(n8476[15]), .I2(GND_net), 
            .I3(n38080), .O(n8452[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_22 (.CI(n37663), .I0(n7960[19]), .I1(GND_net), 
            .CO(n37664));
    SB_LUT4 add_3501_7_lut (.I0(GND_net), .I1(n16575[4]), .I2(n649), .I3(n36782), 
            .O(n16509[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_7 (.CI(n36782), .I0(n16575[4]), .I1(n649), .CO(n36783));
    SB_LUT4 unary_minus_70_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n73[9]), 
            .I3(n36607), .O(n852[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_21 (.CI(n38387), .I0(n8452[18]), .I1(GND_net), 
            .CO(n38388));
    SB_CARRY add_3108_18 (.CI(n38080), .I0(n8476[15]), .I1(GND_net), .CO(n38081));
    SB_LUT4 mult_12_add_2137_21_lut (.I0(GND_net), .I1(n7960[18]), .I2(GND_net), 
            .I3(n37662), .O(n191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_17_lut (.I0(GND_net), .I1(n8476[14]), .I2(GND_net), 
            .I3(n38079), .O(n8452[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_21 (.CI(n37662), .I0(n7960[18]), .I1(GND_net), 
            .CO(n37663));
    SB_LUT4 add_3501_6_lut (.I0(GND_net), .I1(n16575[3]), .I2(n552), .I3(n36781), 
            .O(n16509[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_17 (.CI(n38079), .I0(n8476[14]), .I1(GND_net), .CO(n38080));
    SB_CARRY unary_minus_70_add_3_11 (.CI(n36607), .I0(GND_net), .I1(n73[9]), 
            .CO(n36608));
    SB_CARRY add_3501_6 (.CI(n36781), .I0(n16575[3]), .I1(n552), .CO(n36782));
    SB_LUT4 mult_12_add_2137_20_lut (.I0(GND_net), .I1(n7960[17]), .I2(GND_net), 
            .I3(n37661), .O(n191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n73[8]), 
            .I3(n36606), .O(n868)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_20 (.CI(n37661), .I0(n7960[17]), .I1(GND_net), 
            .CO(n37662));
    SB_LUT4 mult_12_add_2137_19_lut (.I0(GND_net), .I1(n7960[16]), .I2(GND_net), 
            .I3(n37660), .O(n191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_10 (.CI(n36606), .I0(GND_net), .I1(n73[8]), 
            .CO(n36607));
    SB_CARRY mult_12_add_2137_19 (.CI(n37660), .I0(n7960[16]), .I1(GND_net), 
            .CO(n37661));
    SB_LUT4 add_3108_16_lut (.I0(GND_net), .I1(n8476[13]), .I2(GND_net), 
            .I3(n38078), .O(n8452[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_18_lut (.I0(GND_net), .I1(n7960[15]), .I2(GND_net), 
            .I3(n37659), .O(n191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_20_lut (.I0(GND_net), .I1(n8452[17]), .I2(GND_net), 
            .I3(n38386), .O(n1804[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_16 (.CI(n38078), .I0(n8476[13]), .I1(GND_net), .CO(n38079));
    SB_CARRY mult_14_add_1219_20 (.CI(n38386), .I0(n8452[17]), .I1(GND_net), 
            .CO(n38387));
    SB_LUT4 unary_minus_70_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n73[7]), 
            .I3(n36605), .O(n869)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_15_lut (.I0(GND_net), .I1(n8476[12]), .I2(GND_net), 
            .I3(n38077), .O(n8452[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_18 (.CI(n37659), .I0(n7960[15]), .I1(GND_net), 
            .CO(n37660));
    SB_LUT4 mult_12_add_2137_17_lut (.I0(GND_net), .I1(n7960[14]), .I2(GND_net), 
            .I3(n37658), .O(n191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_9 (.CI(n36605), .I0(GND_net), .I1(n73[7]), 
            .CO(n36606));
    SB_CARRY add_3108_15 (.CI(n38077), .I0(n8476[12]), .I1(GND_net), .CO(n38078));
    SB_LUT4 add_3501_5_lut (.I0(GND_net), .I1(n16575[2]), .I2(n455_adj_3588), 
            .I3(n36780), .O(n16509[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_31_lut (.I0(GND_net), .I1(n7764[28]), .I2(GND_net), 
            .I3(n37155), .O(n6546[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_17 (.CI(n37658), .I0(n7960[14]), .I1(GND_net), 
            .CO(n37659));
    SB_LUT4 add_3010_30_lut (.I0(GND_net), .I1(n7764[27]), .I2(GND_net), 
            .I3(n37154), .O(n6546[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_16_lut (.I0(GND_net), .I1(n7960[13]), .I2(GND_net), 
            .I3(n37657), .O(n191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_16 (.CI(n37657), .I0(n7960[13]), .I1(GND_net), 
            .CO(n37658));
    SB_LUT4 mult_14_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_add_2137_15_lut (.I0(GND_net), .I1(n7960[12]), .I2(GND_net), 
            .I3(n37656), .O(n191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_30 (.CI(n37154), .I0(n7764[27]), .I1(GND_net), .CO(n37155));
    SB_LUT4 add_3108_14_lut (.I0(GND_net), .I1(n8476[11]), .I2(GND_net), 
            .I3(n38076), .O(n8452[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_15 (.CI(n37656), .I0(n7960[12]), .I1(GND_net), 
            .CO(n37657));
    SB_LUT4 add_3010_29_lut (.I0(GND_net), .I1(n7764[26]), .I2(GND_net), 
            .I3(n37153), .O(n6546[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_29 (.CI(n37153), .I0(n7764[26]), .I1(GND_net), .CO(n37154));
    SB_LUT4 add_3010_28_lut (.I0(GND_net), .I1(n7764[25]), .I2(GND_net), 
            .I3(n37152), .O(n6546[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_5 (.CI(n36780), .I0(n16575[2]), .I1(n455_adj_3588), 
            .CO(n36781));
    SB_LUT4 mult_12_add_2137_14_lut (.I0(GND_net), .I1(n7960[11]), .I2(GND_net), 
            .I3(n37655), .O(n191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n73[6]), 
            .I3(n36604), .O(n870)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_28 (.CI(n37152), .I0(n7764[25]), .I1(GND_net), .CO(n37153));
    SB_CARRY add_3108_14 (.CI(n38076), .I0(n8476[11]), .I1(GND_net), .CO(n38077));
    SB_LUT4 add_3501_4_lut (.I0(GND_net), .I1(n16575[1]), .I2(n358), .I3(n36779), 
            .O(n16509[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i282_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n419_adj_3432));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3010_27_lut (.I0(GND_net), .I1(n7764[24]), .I2(GND_net), 
            .I3(n37151), .O(n6546[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_19_lut (.I0(GND_net), .I1(n8452[16]), .I2(GND_net), 
            .I3(n38385), .O(n1804[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_14 (.CI(n37655), .I0(n7960[11]), .I1(GND_net), 
            .CO(n37656));
    SB_LUT4 add_3108_13_lut (.I0(GND_net), .I1(n8476[10]), .I2(GND_net), 
            .I3(n38075), .O(n8452[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_19 (.CI(n38385), .I0(n8452[16]), .I1(GND_net), 
            .CO(n38386));
    SB_CARRY unary_minus_70_add_3_8 (.CI(n36604), .I0(GND_net), .I1(n73[6]), 
            .CO(n36605));
    SB_CARRY add_3501_4 (.CI(n36779), .I0(n16575[1]), .I1(n358), .CO(n36780));
    SB_CARRY add_3010_27 (.CI(n37151), .I0(n7764[24]), .I1(GND_net), .CO(n37152));
    SB_LUT4 mult_12_add_2137_13_lut (.I0(GND_net), .I1(n7960[10]), .I2(GND_net), 
            .I3(n37654), .O(n191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_26_lut (.I0(GND_net), .I1(n7764[23]), .I2(GND_net), 
            .I3(n37150), .O(n6546[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n73[5]), 
            .I3(n36603), .O(n871)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_7 (.CI(n36603), .I0(GND_net), .I1(n73[5]), 
            .CO(n36604));
    SB_CARRY add_3010_26 (.CI(n37150), .I0(n7764[23]), .I1(GND_net), .CO(n37151));
    SB_LUT4 mult_12_i341_2_lut (.I0(\Kd[5] ), .I1(n67[7]), .I2(GND_net), 
            .I3(GND_net), .O(n507));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[13]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3010_25_lut (.I0(GND_net), .I1(n7764[22]), .I2(GND_net), 
            .I3(n37149), .O(n6546[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_13 (.CI(n37654), .I0(n7960[10]), .I1(GND_net), 
            .CO(n37655));
    SB_CARRY add_3108_13 (.CI(n38075), .I0(n8476[10]), .I1(GND_net), .CO(n38076));
    SB_LUT4 add_3108_12_lut (.I0(GND_net), .I1(n8476[9]), .I2(GND_net), 
            .I3(n38074), .O(n8452[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_12_lut (.I0(GND_net), .I1(n7960[9]), .I2(GND_net), 
            .I3(n37653), .O(n191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[3]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[14]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3010_25 (.CI(n37149), .I0(n7764[22]), .I1(GND_net), .CO(n37150));
    SB_CARRY mult_12_add_2137_12 (.CI(n37653), .I0(n7960[9]), .I1(GND_net), 
            .CO(n37654));
    SB_LUT4 add_3010_24_lut (.I0(GND_net), .I1(n7764[21]), .I2(GND_net), 
            .I3(n37148), .O(n6546[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_24 (.CI(n37148), .I0(n7764[21]), .I1(GND_net), .CO(n37149));
    SB_CARRY add_3108_12 (.CI(n38074), .I0(n8476[9]), .I1(GND_net), .CO(n38075));
    SB_LUT4 mult_12_add_2137_11_lut (.I0(GND_net), .I1(n7960[8]), .I2(GND_net), 
            .I3(n37652), .O(n191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_23_lut (.I0(GND_net), .I1(n7764[20]), .I2(GND_net), 
            .I3(n37147), .O(n6546[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3501_3_lut (.I0(GND_net), .I1(n16575[0]), .I2(n261), .I3(n36778), 
            .O(n16509[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_18_lut (.I0(GND_net), .I1(n8452[15]), .I2(GND_net), 
            .I3(n38384), .O(n1804[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_11_lut (.I0(GND_net), .I1(n8476[8]), .I2(GND_net), 
            .I3(n38073), .O(n8452[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_23 (.CI(n37147), .I0(n7764[20]), .I1(GND_net), .CO(n37148));
    SB_LUT4 unary_minus_70_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n73[4]), 
            .I3(n36602), .O(n872)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_3 (.CI(n36778), .I0(n16575[0]), .I1(n261), .CO(n36779));
    SB_CARRY mult_12_add_2137_11 (.CI(n37652), .I0(n7960[8]), .I1(GND_net), 
            .CO(n37653));
    SB_CARRY mult_14_add_1219_18 (.CI(n38384), .I0(n8452[15]), .I1(GND_net), 
            .CO(n38385));
    SB_CARRY add_3108_11 (.CI(n38073), .I0(n8476[8]), .I1(GND_net), .CO(n38074));
    SB_LUT4 add_3010_22_lut (.I0(GND_net), .I1(n7764[19]), .I2(GND_net), 
            .I3(n37146), .O(n6546[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_10_lut (.I0(GND_net), .I1(n7960[7]), .I2(GND_net), 
            .I3(n37651), .O(n191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_22 (.CI(n37146), .I0(n7764[19]), .I1(GND_net), .CO(n37147));
    SB_CARRY unary_minus_70_add_3_6 (.CI(n36602), .I0(GND_net), .I1(n73[4]), 
            .CO(n36603));
    SB_LUT4 add_3010_21_lut (.I0(GND_net), .I1(n7764[18]), .I2(GND_net), 
            .I3(n37145), .O(n6546[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_17_lut (.I0(GND_net), .I1(n8452[14]), .I2(GND_net), 
            .I3(n38383), .O(n1804[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_10_lut (.I0(GND_net), .I1(n8476[7]), .I2(GND_net), 
            .I3(n38072), .O(n8452[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_10 (.CI(n37651), .I0(n7960[7]), .I1(GND_net), 
            .CO(n37652));
    SB_CARRY add_3010_21 (.CI(n37145), .I0(n7764[18]), .I1(GND_net), .CO(n37146));
    SB_LUT4 mult_12_add_2137_9_lut (.I0(GND_net), .I1(n7960[6]), .I2(GND_net), 
            .I3(n37650), .O(n191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_10 (.CI(n38072), .I0(n8476[7]), .I1(GND_net), .CO(n38073));
    SB_LUT4 add_3501_2_lut (.I0(GND_net), .I1(n71), .I2(n164), .I3(GND_net), 
            .O(n16509[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_9 (.CI(n37650), .I0(n7960[6]), .I1(GND_net), 
            .CO(n37651));
    SB_LUT4 add_3108_9_lut (.I0(GND_net), .I1(n8476[6]), .I2(GND_net), 
            .I3(n38071), .O(n8452[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_17 (.CI(n38383), .I0(n8452[14]), .I1(GND_net), 
            .CO(n38384));
    SB_CARRY add_3501_2 (.CI(GND_net), .I0(n71), .I1(n164), .CO(n36778));
    SB_LUT4 add_3010_20_lut (.I0(GND_net), .I1(n7764[17]), .I2(GND_net), 
            .I3(n37144), .O(n6546[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_8_lut (.I0(GND_net), .I1(n7960[5]), .I2(n680_adj_3597), 
            .I3(n37649), .O(n191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_8 (.CI(n37649), .I0(n7960[5]), .I1(n680_adj_3597), 
            .CO(n37650));
    SB_CARRY add_3010_20 (.CI(n37144), .I0(n7764[17]), .I1(GND_net), .CO(n37145));
    SB_CARRY add_3108_9 (.CI(n38071), .I0(n8476[6]), .I1(GND_net), .CO(n38072));
    SB_LUT4 add_3010_19_lut (.I0(GND_net), .I1(n7764[16]), .I2(GND_net), 
            .I3(n37143), .O(n6546[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_7_lut (.I0(GND_net), .I1(n7960[4]), .I2(n583_adj_3598), 
            .I3(n37648), .O(n191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_19 (.CI(n37143), .I0(n7764[16]), .I1(GND_net), .CO(n37144));
    SB_LUT4 add_3010_18_lut (.I0(GND_net), .I1(n7764[15]), .I2(GND_net), 
            .I3(n37142), .O(n6546[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n516_adj_3428));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3010_18 (.CI(n37142), .I0(n7764[15]), .I1(GND_net), .CO(n37143));
    SB_LUT4 unary_minus_70_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n73[3]), 
            .I3(n36601), .O(n873)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_17_lut (.I0(GND_net), .I1(n7764[14]), .I2(GND_net), 
            .I3(n37141), .O(n6546[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i406_2_lut (.I0(\Kd[6] ), .I1(n67[7]), .I2(GND_net), 
            .I3(GND_net), .O(n604));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[15]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_12_add_2137_7 (.CI(n37648), .I0(n7960[4]), .I1(n583_adj_3598), 
            .CO(n37649));
    SB_CARRY unary_minus_70_add_3_5 (.CI(n36601), .I0(GND_net), .I1(n73[3]), 
            .CO(n36602));
    SB_LUT4 unary_minus_70_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n73[2]), 
            .I3(n36600), .O(n874)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_16_lut (.I0(GND_net), .I1(n8452[13]), .I2(GND_net), 
            .I3(n38382), .O(n1804[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_8_lut (.I0(GND_net), .I1(n8476[5]), .I2(n545), .I3(n38070), 
            .O(n8452[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_6_lut (.I0(GND_net), .I1(n7960[3]), .I2(n486_adj_3601), 
            .I3(n37647), .O(n191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_4 (.CI(n36600), .I0(GND_net), .I1(n73[2]), 
            .CO(n36601));
    SB_CARRY mult_14_add_1219_16 (.CI(n38382), .I0(n8452[13]), .I1(GND_net), 
            .CO(n38383));
    SB_CARRY add_3108_8 (.CI(n38070), .I0(n8476[5]), .I1(n545), .CO(n38071));
    SB_CARRY mult_12_add_2137_6 (.CI(n37647), .I0(n7960[3]), .I1(n486_adj_3601), 
            .CO(n37648));
    SB_LUT4 mult_12_add_2137_5_lut (.I0(GND_net), .I1(n7960[2]), .I2(n389_adj_3603), 
            .I3(n37646), .O(n191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_7_lut (.I0(GND_net), .I1(n8476[4]), .I2(n472), .I3(n38069), 
            .O(n8452[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_17 (.CI(n37141), .I0(n7764[14]), .I1(GND_net), .CO(n37142));
    SB_CARRY mult_12_add_2137_5 (.CI(n37646), .I0(n7960[2]), .I1(n389_adj_3603), 
            .CO(n37647));
    SB_LUT4 mult_14_add_1219_15_lut (.I0(GND_net), .I1(n8452[12]), .I2(GND_net), 
            .I3(n38381), .O(n1804[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_16_lut (.I0(GND_net), .I1(n7764[13]), .I2(GND_net), 
            .I3(n37140), .O(n6546[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_15 (.CI(n38381), .I0(n8452[12]), .I1(GND_net), 
            .CO(n38382));
    SB_CARRY add_3108_7 (.CI(n38069), .I0(n8476[4]), .I1(n472), .CO(n38070));
    SB_LUT4 mult_12_add_2137_4_lut (.I0(GND_net), .I1(n7960[1]), .I2(n292_adj_3604), 
            .I3(n37645), .O(n191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_4 (.CI(n37645), .I0(n7960[1]), .I1(n292_adj_3604), 
            .CO(n37646));
    SB_CARRY add_3010_16 (.CI(n37140), .I0(n7764[13]), .I1(GND_net), .CO(n37141));
    SB_LUT4 mult_14_add_1219_14_lut (.I0(GND_net), .I1(n8452[11]), .I2(GND_net), 
            .I3(n38380), .O(n1804[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_6_lut (.I0(GND_net), .I1(n8476[3]), .I2(n399), .I3(n38068), 
            .O(n8452[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_3_lut (.I0(GND_net), .I1(n7960[0]), .I2(n195_adj_3605), 
            .I3(n37644), .O(n191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_15_lut (.I0(GND_net), .I1(n7764[12]), .I2(GND_net), 
            .I3(n37139), .O(n6546[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_3 (.CI(n37644), .I0(n7960[0]), .I1(n195_adj_3605), 
            .CO(n37645));
    SB_LUT4 mult_12_add_2137_2_lut (.I0(GND_net), .I1(n5_adj_3607), .I2(n98_adj_3608), 
            .I3(GND_net), .O(n191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_15 (.CI(n37139), .I0(n7764[12]), .I1(GND_net), .CO(n37140));
    SB_LUT4 add_3010_14_lut (.I0(GND_net), .I1(n7764[11]), .I2(GND_net), 
            .I3(n37138), .O(n6546[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n73[1]), 
            .I3(n36599), .O(n875)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_6 (.CI(n38068), .I0(n8476[3]), .I1(n399), .CO(n38069));
    SB_CARRY mult_12_add_2137_2 (.CI(GND_net), .I0(n5_adj_3607), .I1(n98_adj_3608), 
            .CO(n37644));
    SB_LUT4 add_3149_21_lut (.I0(GND_net), .I1(n10122[18]), .I2(GND_net), 
            .I3(n37643), .O(n9331[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_14 (.CI(n37138), .I0(n7764[11]), .I1(GND_net), .CO(n37139));
    SB_CARRY unary_minus_70_add_3_3 (.CI(n36599), .I0(GND_net), .I1(n73[1]), 
            .CO(n36600));
    SB_LUT4 add_3010_13_lut (.I0(GND_net), .I1(n7764[10]), .I2(GND_net), 
            .I3(n37137), .O(n6546[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_5_lut (.I0(GND_net), .I1(n8476[2]), .I2(n326), .I3(n38067), 
            .O(n8452[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_20_lut (.I0(GND_net), .I1(n10122[17]), .I2(GND_net), 
            .I3(n37642), .O(n9331[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_13 (.CI(n37137), .I0(n7764[10]), .I1(GND_net), .CO(n37138));
    SB_CARRY add_3149_20 (.CI(n37642), .I0(n10122[17]), .I1(GND_net), 
            .CO(n37643));
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n613_adj_3426));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3010_12_lut (.I0(GND_net), .I1(n7764[9]), .I2(GND_net), 
            .I3(n37136), .O(n6546[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_19_lut (.I0(GND_net), .I1(n10122[16]), .I2(GND_net), 
            .I3(n37641), .O(n9331[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_14 (.CI(n38380), .I0(n8452[11]), .I1(GND_net), 
            .CO(n38381));
    SB_CARRY add_3108_5 (.CI(n38067), .I0(n8476[2]), .I1(n326), .CO(n38068));
    SB_CARRY add_3149_19 (.CI(n37641), .I0(n10122[16]), .I1(GND_net), 
            .CO(n37642));
    SB_CARRY add_3010_12 (.CI(n37136), .I0(n7764[9]), .I1(GND_net), .CO(n37137));
    SB_LUT4 unary_minus_70_add_3_2_lut (.I0(n28668), .I1(GND_net), .I2(n73[0]), 
            .I3(VCC_net), .O(n46539)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3108_4_lut (.I0(GND_net), .I1(n8476[1]), .I2(n253), .I3(n38066), 
            .O(n8452[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_4 (.CI(n38066), .I0(n8476[1]), .I1(n253), .CO(n38067));
    SB_LUT4 mult_14_add_1219_13_lut (.I0(GND_net), .I1(n8452[10]), .I2(GND_net), 
            .I3(n38379), .O(n1804[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_3_lut (.I0(GND_net), .I1(n8476[0]), .I2(n180_adj_3552), 
            .I3(n38065), .O(n8452[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_18_lut (.I0(GND_net), .I1(n10122[15]), .I2(GND_net), 
            .I3(n37640), .O(n9331[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_11_lut (.I0(GND_net), .I1(n7764[8]), .I2(GND_net), 
            .I3(n37135), .O(n6546[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_18 (.CI(n37640), .I0(n10122[15]), .I1(GND_net), 
            .CO(n37641));
    SB_CARRY add_3010_11 (.CI(n37135), .I0(n7764[8]), .I1(GND_net), .CO(n37136));
    SB_LUT4 add_3010_10_lut (.I0(GND_net), .I1(n7764[7]), .I2(GND_net), 
            .I3(n37134), .O(n6546[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_3 (.CI(n38065), .I0(n8476[0]), .I1(n180_adj_3552), 
            .CO(n38066));
    SB_LUT4 add_3149_17_lut (.I0(GND_net), .I1(n10122[14]), .I2(GND_net), 
            .I3(n37639), .O(n9331[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_10 (.CI(n37134), .I0(n7764[7]), .I1(GND_net), .CO(n37135));
    SB_CARRY add_3149_17 (.CI(n37639), .I0(n10122[14]), .I1(GND_net), 
            .CO(n37640));
    SB_LUT4 add_3010_9_lut (.I0(GND_net), .I1(n7764[6]), .I2(GND_net), 
            .I3(n37133), .O(n6546[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[16]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3010_9 (.CI(n37133), .I0(n7764[6]), .I1(GND_net), .CO(n37134));
    SB_CARRY mult_14_add_1219_13 (.CI(n38379), .I0(n8452[10]), .I1(GND_net), 
            .CO(n38380));
    SB_LUT4 mult_14_add_1219_12_lut (.I0(GND_net), .I1(n8452[9]), .I2(GND_net), 
            .I3(n38378), .O(n1804[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_8_lut (.I0(GND_net), .I1(n7764[5]), .I2(n683), .I3(n37132), 
            .O(n6546[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_12 (.CI(n38378), .I0(n8452[9]), .I1(GND_net), 
            .CO(n38379));
    SB_LUT4 add_3108_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n8452[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_16_lut (.I0(GND_net), .I1(n10122[13]), .I2(GND_net), 
            .I3(n37638), .O(n9331[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_8 (.CI(n37132), .I0(n7764[5]), .I1(n683), .CO(n37133));
    SB_CARRY add_3108_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n38065));
    SB_CARRY add_3149_16 (.CI(n37638), .I0(n10122[13]), .I1(GND_net), 
            .CO(n37639));
    SB_LUT4 add_3010_7_lut (.I0(GND_net), .I1(n7764[4]), .I2(n586), .I3(n37131), 
            .O(n6546[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_15_lut (.I0(GND_net), .I1(n10122[12]), .I2(GND_net), 
            .I3(n37637), .O(n9331[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_15 (.CI(n37637), .I0(n10122[12]), .I1(GND_net), 
            .CO(n37638));
    SB_CARRY add_3010_7 (.CI(n37131), .I0(n7764[4]), .I1(n586), .CO(n37132));
    SB_LUT4 add_3010_6_lut (.I0(GND_net), .I1(n7764[3]), .I2(n489), .I3(n37130), 
            .O(n6546[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_6 (.CI(n37130), .I0(n7764[3]), .I1(n489), .CO(n37131));
    SB_LUT4 add_3107_8_lut (.I0(GND_net), .I1(n9323[5]), .I2(n752_adj_3611), 
            .I3(n38064), .O(n8443[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_14_lut (.I0(GND_net), .I1(n10122[11]), .I2(GND_net), 
            .I3(n37636), .O(n9331[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3107_7_lut (.I0(GND_net), .I1(n9323[4]), .I2(n655), .I3(n38063), 
            .O(n8443[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_5_lut (.I0(GND_net), .I1(n7764[2]), .I2(n392), .I3(n37129), 
            .O(n6546[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_14 (.CI(n37636), .I0(n10122[11]), .I1(GND_net), 
            .CO(n37637));
    SB_CARRY add_3010_5 (.CI(n37129), .I0(n7764[2]), .I1(n392), .CO(n37130));
    SB_LUT4 add_3010_4_lut (.I0(GND_net), .I1(n7764[1]), .I2(n295_adj_3612), 
            .I3(n37128), .O(n6546[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_4 (.CI(n37128), .I0(n7764[1]), .I1(n295_adj_3612), 
            .CO(n37129));
    SB_CARRY add_3107_7 (.CI(n38063), .I0(n9323[4]), .I1(n655), .CO(n38064));
    SB_LUT4 add_3149_13_lut (.I0(GND_net), .I1(n10122[10]), .I2(GND_net), 
            .I3(n37635), .O(n9331[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_13 (.CI(n37635), .I0(n10122[10]), .I1(GND_net), 
            .CO(n37636));
    SB_LUT4 add_3107_6_lut (.I0(GND_net), .I1(n9323[3]), .I2(n558_adj_3613), 
            .I3(n38062), .O(n8443[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_12_lut (.I0(GND_net), .I1(n10122[9]), .I2(GND_net), 
            .I3(n37634), .O(n9331[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_3_lut (.I0(GND_net), .I1(n7764[0]), .I2(n198), .I3(n37127), 
            .O(n6546[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_3 (.CI(n37127), .I0(n7764[0]), .I1(n198), .CO(n37128));
    SB_LUT4 add_3010_2_lut (.I0(GND_net), .I1(n8_adj_3614), .I2(n101), 
            .I3(GND_net), .O(n6546[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_12 (.CI(n37634), .I0(n10122[9]), .I1(GND_net), .CO(n37635));
    SB_CARRY add_3010_2 (.CI(GND_net), .I0(n8_adj_3614), .I1(n101), .CO(n37127));
    SB_LUT4 add_3077_30_lut (.I0(GND_net), .I1(n9129[27]), .I2(GND_net), 
            .I3(n37126), .O(n7764[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_11_lut (.I0(GND_net), .I1(n10122[8]), .I2(GND_net), 
            .I3(n37633), .O(n9331[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_11_lut (.I0(GND_net), .I1(n8452[8]), .I2(GND_net), 
            .I3(n38377), .O(n1804[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3107_6 (.CI(n38062), .I0(n9323[3]), .I1(n558_adj_3613), 
            .CO(n38063));
    SB_LUT4 add_3107_5_lut (.I0(GND_net), .I1(n9323[2]), .I2(n461_c), 
            .I3(n38061), .O(n8443[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_11 (.CI(n37633), .I0(n10122[8]), .I1(GND_net), .CO(n37634));
    SB_LUT4 add_3077_29_lut (.I0(GND_net), .I1(n9129[26]), .I2(GND_net), 
            .I3(n37125), .O(n7764[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_10_lut (.I0(GND_net), .I1(n10122[7]), .I2(GND_net), 
            .I3(n37632), .O(n9331[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_10 (.CI(n37632), .I0(n10122[7]), .I1(GND_net), .CO(n37633));
    SB_LUT4 add_3149_9_lut (.I0(GND_net), .I1(n10122[6]), .I2(GND_net), 
            .I3(n37631), .O(n9331[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_9 (.CI(n37631), .I0(n10122[6]), .I1(GND_net), .CO(n37632));
    SB_CARRY add_3077_29 (.CI(n37125), .I0(n9129[26]), .I1(GND_net), .CO(n37126));
    SB_LUT4 add_22497_33_lut (.I0(GND_net), .I1(n79[31]), .I2(n7065[0]), 
            .I3(n36772), .O(\PID_CONTROLLER.result_31__N_2994 [31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_28_lut (.I0(GND_net), .I1(n9129[25]), .I2(GND_net), 
            .I3(n37124), .O(n7764[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_32_lut (.I0(GND_net), .I1(n79[30]), .I2(n191[30]), 
            .I3(n36771), .O(\PID_CONTROLLER.result_31__N_2994 [30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n73[0]), 
            .CO(n36599));
    SB_CARRY mult_14_add_1219_11 (.CI(n38377), .I0(n8452[8]), .I1(GND_net), 
            .CO(n38378));
    SB_CARRY add_3107_5 (.CI(n38061), .I0(n9323[2]), .I1(n461_c), .CO(n38062));
    SB_LUT4 add_3149_8_lut (.I0(GND_net), .I1(n10122[5]), .I2(n545), .I3(n37630), 
            .O(n9331[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_28 (.CI(n37124), .I0(n9129[25]), .I1(GND_net), .CO(n37125));
    SB_LUT4 add_3077_27_lut (.I0(GND_net), .I1(n9129[24]), .I2(GND_net), 
            .I3(n37123), .O(n7764[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_27 (.CI(n37123), .I0(n9129[24]), .I1(GND_net), .CO(n37124));
    SB_LUT4 mult_10_i477_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n710_adj_3424));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i471_2_lut (.I0(\Kd[7] ), .I1(n67[7]), .I2(GND_net), 
            .I3(GND_net), .O(n701));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1219_10_lut (.I0(GND_net), .I1(n8452[7]), .I2(GND_net), 
            .I3(n38376), .O(n1804[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_26_lut (.I0(GND_net), .I1(n9129[23]), .I2(GND_net), 
            .I3(n37122), .O(n7764[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_26 (.CI(n37122), .I0(n9129[23]), .I1(GND_net), .CO(n37123));
    SB_LUT4 add_3107_4_lut (.I0(GND_net), .I1(n9323[1]), .I2(n364), .I3(n38060), 
            .O(n8443[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_8 (.CI(n37630), .I0(n10122[5]), .I1(n545), .CO(n37631));
    SB_LUT4 add_3077_25_lut (.I0(GND_net), .I1(n9129[22]), .I2(GND_net), 
            .I3(n37121), .O(n7764[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_32 (.CI(n36771), .I0(n79[30]), .I1(n191[30]), .CO(n36772));
    SB_CARRY add_3077_25 (.CI(n37121), .I0(n9129[22]), .I1(GND_net), .CO(n37122));
    SB_LUT4 add_22497_31_lut (.I0(GND_net), .I1(n79[29]), .I2(n191[29]), 
            .I3(n36770), .O(\PID_CONTROLLER.result_31__N_2994 [29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_10 (.CI(n38376), .I0(n8452[7]), .I1(GND_net), 
            .CO(n38377));
    SB_CARRY add_3107_4 (.CI(n38060), .I0(n9323[1]), .I1(n364), .CO(n38061));
    SB_LUT4 add_3149_7_lut (.I0(GND_net), .I1(n10122[4]), .I2(n472), .I3(n37629), 
            .O(n9331[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_24_lut (.I0(GND_net), .I1(n9129[21]), .I2(GND_net), 
            .I3(n37120), .O(n7764[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_24 (.CI(n37120), .I0(n9129[21]), .I1(GND_net), .CO(n37121));
    SB_LUT4 add_3107_3_lut (.I0(GND_net), .I1(n9323[0]), .I2(n267), .I3(n38059), 
            .O(n8443[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_7 (.CI(n37629), .I0(n10122[4]), .I1(n472), .CO(n37630));
    SB_LUT4 add_3077_23_lut (.I0(GND_net), .I1(n9129[20]), .I2(GND_net), 
            .I3(n37119), .O(n7764[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_31 (.CI(n36770), .I0(n79[29]), .I1(n191[29]), .CO(n36771));
    SB_CARRY add_3077_23 (.CI(n37119), .I0(n9129[20]), .I1(GND_net), .CO(n37120));
    SB_LUT4 add_22497_30_lut (.I0(GND_net), .I1(n79[28]), .I2(n191[28]), 
            .I3(n36769), .O(\PID_CONTROLLER.result_31__N_2994 [28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_9_lut (.I0(GND_net), .I1(n8452[6]), .I2(GND_net), 
            .I3(n38375), .O(n1804[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3107_3 (.CI(n38059), .I0(n9323[0]), .I1(n267), .CO(n38060));
    SB_LUT4 add_3149_6_lut (.I0(GND_net), .I1(n10122[3]), .I2(n399), .I3(n37628), 
            .O(n9331[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_6 (.CI(n37628), .I0(n10122[3]), .I1(n399), .CO(n37629));
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[17]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3077_22_lut (.I0(GND_net), .I1(n9129[19]), .I2(GND_net), 
            .I3(n37118), .O(n7764[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3107_2_lut (.I0(GND_net), .I1(n86_adj_3617), .I2(n170_adj_3618), 
            .I3(GND_net), .O(n8443[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_5_lut (.I0(GND_net), .I1(n10122[2]), .I2(n326), .I3(n37627), 
            .O(n9331[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3107_2 (.CI(GND_net), .I0(n86_adj_3617), .I1(n170_adj_3618), 
            .CO(n38059));
    SB_CARRY add_3149_5 (.CI(n37627), .I0(n10122[2]), .I1(n326), .CO(n37628));
    SB_CARRY add_3077_22 (.CI(n37118), .I0(n9129[19]), .I1(GND_net), .CO(n37119));
    SB_LUT4 add_3077_21_lut (.I0(GND_net), .I1(n9129[18]), .I2(GND_net), 
            .I3(n37117), .O(n7764[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3106_9_lut (.I0(GND_net), .I1(n8443[6]), .I2(GND_net), 
            .I3(n38058), .O(n8433[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_4_lut (.I0(GND_net), .I1(n10122[1]), .I2(n253), .I3(n37626), 
            .O(n9331[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_21 (.CI(n37117), .I0(n9129[18]), .I1(GND_net), .CO(n37118));
    SB_CARRY add_22497_30 (.CI(n36769), .I0(n79[28]), .I1(n191[28]), .CO(n36770));
    SB_LUT4 add_3077_20_lut (.I0(GND_net), .I1(n9129[17]), .I2(GND_net), 
            .I3(n37116), .O(n7764[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_29_lut (.I0(GND_net), .I1(n79[27]), .I2(n191[27]), 
            .I3(n36768), .O(\PID_CONTROLLER.result_31__N_2994 [27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_9 (.CI(n38375), .I0(n8452[6]), .I1(GND_net), 
            .CO(n38376));
    SB_LUT4 add_3106_8_lut (.I0(GND_net), .I1(n8443[5]), .I2(n749_adj_3619), 
            .I3(n38057), .O(n8433[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_4 (.CI(n37626), .I0(n10122[1]), .I1(n253), .CO(n37627));
    SB_CARRY add_3077_20 (.CI(n37116), .I0(n9129[17]), .I1(GND_net), .CO(n37117));
    SB_LUT4 add_3077_19_lut (.I0(GND_net), .I1(n9129[16]), .I2(GND_net), 
            .I3(n37115), .O(n7764[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3106_8 (.CI(n38057), .I0(n8443[5]), .I1(n749_adj_3619), 
            .CO(n38058));
    SB_LUT4 add_3149_3_lut (.I0(GND_net), .I1(n10122[0]), .I2(n180_adj_3552), 
            .I3(n37625), .O(n9331[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_19 (.CI(n37115), .I0(n9129[16]), .I1(GND_net), .CO(n37116));
    SB_CARRY add_22497_29 (.CI(n36768), .I0(n79[27]), .I1(n191[27]), .CO(n36769));
    SB_LUT4 add_3077_18_lut (.I0(GND_net), .I1(n9129[15]), .I2(GND_net), 
            .I3(n37114), .O(n7764[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_3 (.CI(n37625), .I0(n10122[0]), .I1(n180_adj_3552), 
            .CO(n37626));
    SB_CARRY add_3077_18 (.CI(n37114), .I0(n9129[15]), .I1(GND_net), .CO(n37115));
    SB_LUT4 add_22497_28_lut (.I0(GND_net), .I1(n79[26]), .I2(n191[26]), 
            .I3(n36767), .O(\PID_CONTROLLER.result_31__N_2994 [26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_17_lut (.I0(GND_net), .I1(n9129[14]), .I2(GND_net), 
            .I3(n37113), .O(n7764[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_8_lut (.I0(GND_net), .I1(n8452[5]), .I2(n536), 
            .I3(n38374), .O(n1804[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n9331[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3106_7_lut (.I0(GND_net), .I1(n8443[4]), .I2(n652_adj_3621), 
            .I3(n38056), .O(n8433[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_8 (.CI(n38374), .I0(n8452[5]), .I1(n536), 
            .CO(n38375));
    SB_CARRY add_3077_17 (.CI(n37113), .I0(n9129[14]), .I1(GND_net), .CO(n37114));
    SB_CARRY add_3106_7 (.CI(n38056), .I0(n8443[4]), .I1(n652_adj_3621), 
            .CO(n38057));
    SB_CARRY add_3149_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n37625));
    SB_LUT4 add_3148_7_lut (.I0(GND_net), .I1(n44226), .I2(n658_adj_3622), 
            .I3(n37624), .O(n9323[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_16_lut (.I0(GND_net), .I1(n9129[13]), .I2(GND_net), 
            .I3(n37112), .O(n7764[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_6_lut (.I0(GND_net), .I1(n10115[3]), .I2(n564), .I3(n37623), 
            .O(n9323[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_16 (.CI(n37112), .I0(n9129[13]), .I1(GND_net), .CO(n37113));
    SB_CARRY add_3148_6 (.CI(n37623), .I0(n10115[3]), .I1(n564), .CO(n37624));
    SB_LUT4 add_3106_6_lut (.I0(GND_net), .I1(n8443[3]), .I2(n555_adj_3623), 
            .I3(n38055), .O(n8433[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3106_6 (.CI(n38055), .I0(n8443[3]), .I1(n555_adj_3623), 
            .CO(n38056));
    SB_LUT4 add_3148_5_lut (.I0(GND_net), .I1(n10850[2]), .I2(n464_adj_3624), 
            .I3(n37622), .O(n9323[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_15_lut (.I0(GND_net), .I1(n9129[12]), .I2(GND_net), 
            .I3(n37111), .O(n7764[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_15 (.CI(n37111), .I0(n9129[12]), .I1(GND_net), .CO(n37112));
    SB_CARRY add_22497_28 (.CI(n36767), .I0(n79[26]), .I1(n191[26]), .CO(n36768));
    SB_CARRY add_3148_5 (.CI(n37622), .I0(n10850[2]), .I1(n464_adj_3624), 
            .CO(n37623));
    SB_LUT4 add_3077_14_lut (.I0(GND_net), .I1(n9129[11]), .I2(GND_net), 
            .I3(n37110), .O(n7764[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_27_lut (.I0(GND_net), .I1(n79[25]), .I2(n191[25]), 
            .I3(n36766), .O(\PID_CONTROLLER.result_31__N_2994 [25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_14 (.CI(n37110), .I0(n9129[11]), .I1(GND_net), .CO(n37111));
    SB_LUT4 mult_14_add_1219_7_lut (.I0(GND_net), .I1(n8452[4]), .I2(n463_c), 
            .I3(n38373), .O(n1804[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3106_5_lut (.I0(GND_net), .I1(n8443[2]), .I2(n458_adj_3626), 
            .I3(n38054), .O(n8433[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3106_5 (.CI(n38054), .I0(n8443[2]), .I1(n458_adj_3626), 
            .CO(n38055));
    SB_LUT4 add_3148_4_lut (.I0(GND_net), .I1(n10115[1]), .I2(n370_adj_3627), 
            .I3(n37621), .O(n9323[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_13_lut (.I0(GND_net), .I1(n9129[10]), .I2(GND_net), 
            .I3(n37109), .O(n7764[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_4 (.CI(n37621), .I0(n10115[1]), .I1(n370_adj_3627), 
            .CO(n37622));
    SB_CARRY add_3077_13 (.CI(n37109), .I0(n9129[10]), .I1(GND_net), .CO(n37110));
    SB_LUT4 add_3106_4_lut (.I0(GND_net), .I1(n8443[1]), .I2(n361_adj_3628), 
            .I3(n38053), .O(n8433[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_12_lut (.I0(GND_net), .I1(n9129[9]), .I2(GND_net), 
            .I3(n37108), .O(n7764[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3106_4 (.CI(n38053), .I0(n8443[1]), .I1(n361_adj_3628), 
            .CO(n38054));
    SB_LUT4 add_3148_3_lut (.I0(GND_net), .I1(n10115[0]), .I2(n276_adj_3629), 
            .I3(n37620), .O(n9323[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_3 (.CI(n37620), .I0(n10115[0]), .I1(n276_adj_3629), 
            .CO(n37621));
    SB_CARRY add_3077_12 (.CI(n37108), .I0(n9129[9]), .I1(GND_net), .CO(n37109));
    SB_LUT4 add_3077_11_lut (.I0(GND_net), .I1(n9129[8]), .I2(GND_net), 
            .I3(n37107), .O(n7764[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_27 (.CI(n36766), .I0(n79[25]), .I1(n191[25]), .CO(n36767));
    SB_CARRY add_3077_11 (.CI(n37107), .I0(n9129[8]), .I1(GND_net), .CO(n37108));
    SB_LUT4 add_22497_26_lut (.I0(GND_net), .I1(n79[24]), .I2(n191[24]), 
            .I3(n36765), .O(\PID_CONTROLLER.result_31__N_2994 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_10_lut (.I0(GND_net), .I1(n9129[7]), .I2(GND_net), 
            .I3(n37106), .O(n7764[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_7 (.CI(n38373), .I0(n8452[4]), .I1(n463_c), 
            .CO(n38374));
    SB_LUT4 add_3106_3_lut (.I0(GND_net), .I1(n8443[0]), .I2(n264_adj_3630), 
            .I3(n38052), .O(n8433[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_2_lut (.I0(GND_net), .I1(n86_adj_3617), .I2(n182_adj_3631), 
            .I3(GND_net), .O(n9323[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_6_lut (.I0(GND_net), .I1(n8452[3]), .I2(n390), 
            .I3(n38372), .O(n1804[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_10 (.CI(n37106), .I0(n9129[7]), .I1(GND_net), .CO(n37107));
    SB_LUT4 add_3077_9_lut (.I0(GND_net), .I1(n9129[6]), .I2(GND_net), 
            .I3(n37105), .O(n7764[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_9 (.CI(n37105), .I0(n9129[6]), .I1(GND_net), .CO(n37106));
    SB_CARRY add_3106_3 (.CI(n38052), .I0(n8443[0]), .I1(n264_adj_3630), 
            .CO(n38053));
    SB_CARRY add_3148_2 (.CI(GND_net), .I0(n86_adj_3617), .I1(n182_adj_3631), 
            .CO(n37620));
    SB_LUT4 add_3077_8_lut (.I0(GND_net), .I1(n9129[5]), .I2(n686_adj_3632), 
            .I3(n37104), .O(n7764[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_26 (.CI(n36765), .I0(n79[24]), .I1(n191[24]), .CO(n36766));
    SB_CARRY add_3077_8 (.CI(n37104), .I0(n9129[5]), .I1(n686_adj_3632), 
            .CO(n37105));
    SB_LUT4 add_3106_2_lut (.I0(GND_net), .I1(n74_adj_3633), .I2(n167_adj_3634), 
            .I3(GND_net), .O(n8433[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_25_lut (.I0(GND_net), .I1(n79[23]), .I2(n191[23]), 
            .I3(n36764), .O(\PID_CONTROLLER.result_31__N_2994 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_20_lut (.I0(GND_net), .I1(n10856[17]), .I2(GND_net), 
            .I3(n37619), .O(n10122[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_6 (.CI(n38372), .I0(n8452[3]), .I1(n390), 
            .CO(n38373));
    SB_CARRY add_3106_2 (.CI(GND_net), .I0(n74_adj_3633), .I1(n167_adj_3634), 
            .CO(n38052));
    SB_LUT4 add_3077_7_lut (.I0(GND_net), .I1(n9129[4]), .I2(n589_adj_3635), 
            .I3(n37103), .O(n7764[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_19_lut (.I0(GND_net), .I1(n10856[16]), .I2(GND_net), 
            .I3(n37618), .O(n10122[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_25 (.CI(n36764), .I0(n79[23]), .I1(n191[23]), .CO(n36765));
    SB_CARRY add_3077_7 (.CI(n37103), .I0(n9129[4]), .I1(n589_adj_3635), 
            .CO(n37104));
    SB_CARRY add_3178_19 (.CI(n37618), .I0(n10856[16]), .I1(GND_net), 
            .CO(n37619));
    SB_LUT4 add_3077_6_lut (.I0(GND_net), .I1(n9129[3]), .I2(n492_adj_3636), 
            .I3(n37102), .O(n7764[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_24_lut (.I0(GND_net), .I1(n79[22]), .I2(n191[22]), 
            .I3(n36763), .O(\PID_CONTROLLER.result_31__N_2994 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3105_10_lut (.I0(GND_net), .I1(n8433[7]), .I2(GND_net), 
            .I3(n38051), .O(n8422[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_18_lut (.I0(GND_net), .I1(n10856[15]), .I2(GND_net), 
            .I3(n37617), .O(n10122[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_6 (.CI(n37102), .I0(n9129[3]), .I1(n492_adj_3636), 
            .CO(n37103));
    SB_CARRY add_3178_18 (.CI(n37617), .I0(n10856[15]), .I1(GND_net), 
            .CO(n37618));
    SB_LUT4 add_3077_5_lut (.I0(GND_net), .I1(n9129[2]), .I2(n395_adj_3637), 
            .I3(n37101), .O(n7764[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_24 (.CI(n36763), .I0(n79[22]), .I1(n191[22]), .CO(n36764));
    SB_CARRY add_3077_5 (.CI(n37101), .I0(n9129[2]), .I1(n395_adj_3637), 
            .CO(n37102));
    SB_LUT4 add_3105_9_lut (.I0(GND_net), .I1(n8433[6]), .I2(GND_net), 
            .I3(n38050), .O(n8422[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_17_lut (.I0(GND_net), .I1(n10856[14]), .I2(GND_net), 
            .I3(n37616), .O(n10122[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_23_lut (.I0(GND_net), .I1(n79[21]), .I2(n191[21]), 
            .I3(n36762), .O(\PID_CONTROLLER.result_31__N_2994 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_4_lut (.I0(GND_net), .I1(n9129[1]), .I2(n298_adj_3638), 
            .I3(n37100), .O(n7764[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_4 (.CI(n37100), .I0(n9129[1]), .I1(n298_adj_3638), 
            .CO(n37101));
    SB_LUT4 add_3077_3_lut (.I0(GND_net), .I1(n9129[0]), .I2(n201_adj_3639), 
            .I3(n37099), .O(n7764[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_17 (.CI(n37616), .I0(n10856[14]), .I1(GND_net), 
            .CO(n37617));
    SB_CARRY add_3077_3 (.CI(n37099), .I0(n9129[0]), .I1(n201_adj_3639), 
            .CO(n37100));
    SB_CARRY add_22497_23 (.CI(n36762), .I0(n79[21]), .I1(n191[21]), .CO(n36763));
    SB_LUT4 add_3077_2_lut (.I0(GND_net), .I1(n11_adj_3640), .I2(n104_adj_3641), 
            .I3(GND_net), .O(n7764[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_5_lut (.I0(GND_net), .I1(n8452[2]), .I2(n317), 
            .I3(n38371), .O(n1804[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_9 (.CI(n38050), .I0(n8433[6]), .I1(GND_net), .CO(n38051));
    SB_LUT4 add_3178_16_lut (.I0(GND_net), .I1(n10856[13]), .I2(GND_net), 
            .I3(n37615), .O(n10122[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_16 (.CI(n37615), .I0(n10856[13]), .I1(GND_net), 
            .CO(n37616));
    SB_LUT4 add_3178_15_lut (.I0(GND_net), .I1(n10856[12]), .I2(GND_net), 
            .I3(n37614), .O(n10122[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_5 (.CI(n38371), .I0(n8452[2]), .I1(n317), 
            .CO(n38372));
    SB_LUT4 add_22497_22_lut (.I0(GND_net), .I1(n79[20]), .I2(n191[20]), 
            .I3(n36761), .O(\PID_CONTROLLER.result_31__N_2994 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_15 (.CI(n37614), .I0(n10856[12]), .I1(GND_net), 
            .CO(n37615));
    SB_LUT4 add_3105_8_lut (.I0(GND_net), .I1(n8433[5]), .I2(n746_adj_3642), 
            .I3(n38049), .O(n8422[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_4_lut (.I0(GND_net), .I1(n8452[1]), .I2(n244_adj_3644), 
            .I3(n38370), .O(n1804[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_14_lut (.I0(GND_net), .I1(n10856[11]), .I2(GND_net), 
            .I3(n37613), .O(n10122[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_2 (.CI(GND_net), .I0(n11_adj_3640), .I1(n104_adj_3641), 
            .CO(n37099));
    SB_LUT4 add_3307_15_lut (.I0(GND_net), .I1(n13738[12]), .I2(GND_net), 
            .I3(n37098), .O(n13260[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3307_14_lut (.I0(GND_net), .I1(n13738[11]), .I2(GND_net), 
            .I3(n37097), .O(n13260[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_14 (.CI(n37097), .I0(n13738[11]), .I1(GND_net), 
            .CO(n37098));
    SB_CARRY add_3178_14 (.CI(n37613), .I0(n10856[11]), .I1(GND_net), 
            .CO(n37614));
    SB_LUT4 add_3307_13_lut (.I0(GND_net), .I1(n13738[10]), .I2(GND_net), 
            .I3(n37096), .O(n13260[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_13 (.CI(n37096), .I0(n13738[10]), .I1(GND_net), 
            .CO(n37097));
    SB_CARRY add_3105_8 (.CI(n38049), .I0(n8433[5]), .I1(n746_adj_3642), 
            .CO(n38050));
    SB_LUT4 add_3178_13_lut (.I0(GND_net), .I1(n10856[10]), .I2(GND_net), 
            .I3(n37612), .O(n10122[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_13 (.CI(n37612), .I0(n10856[10]), .I1(GND_net), 
            .CO(n37613));
    SB_LUT4 add_3178_12_lut (.I0(GND_net), .I1(n10856[9]), .I2(GND_net), 
            .I3(n37611), .O(n10122[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3105_7_lut (.I0(GND_net), .I1(n8433[4]), .I2(n649_adj_3645), 
            .I3(n38048), .O(n8422[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_7 (.CI(n38048), .I0(n8433[4]), .I1(n649_adj_3645), 
            .CO(n38049));
    SB_CARRY add_3178_12 (.CI(n37611), .I0(n10856[9]), .I1(GND_net), .CO(n37612));
    SB_LUT4 add_3105_6_lut (.I0(GND_net), .I1(n8433[3]), .I2(n552_adj_3646), 
            .I3(n38047), .O(n8422[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3307_12_lut (.I0(GND_net), .I1(n13738[9]), .I2(GND_net), 
            .I3(n37095), .O(n13260[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_11_lut (.I0(GND_net), .I1(n10856[8]), .I2(GND_net), 
            .I3(n37610), .O(n10122[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_11 (.CI(n37610), .I0(n10856[8]), .I1(GND_net), .CO(n37611));
    SB_LUT4 add_3178_10_lut (.I0(GND_net), .I1(n10856[7]), .I2(GND_net), 
            .I3(n37609), .O(n10122[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_10 (.CI(n37609), .I0(n10856[7]), .I1(GND_net), .CO(n37610));
    SB_LUT4 add_3178_9_lut (.I0(GND_net), .I1(n10856[6]), .I2(GND_net), 
            .I3(n37608), .O(n10122[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_12 (.CI(n37095), .I0(n13738[9]), .I1(GND_net), .CO(n37096));
    SB_CARRY add_3178_9 (.CI(n37608), .I0(n10856[6]), .I1(GND_net), .CO(n37609));
    SB_LUT4 add_3307_11_lut (.I0(GND_net), .I1(n13738[8]), .I2(GND_net), 
            .I3(n37094), .O(n13260[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_11 (.CI(n37094), .I0(n13738[8]), .I1(GND_net), .CO(n37095));
    SB_LUT4 add_3307_10_lut (.I0(GND_net), .I1(n13738[7]), .I2(GND_net), 
            .I3(n37093), .O(n13260[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_8_lut (.I0(GND_net), .I1(n10856[5]), .I2(n545), .I3(n37607), 
            .O(n10122[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_10 (.CI(n37093), .I0(n13738[7]), .I1(GND_net), .CO(n37094));
    SB_LUT4 add_3307_9_lut (.I0(GND_net), .I1(n13738[6]), .I2(GND_net), 
            .I3(n37092), .O(n13260[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_6 (.CI(n38047), .I0(n8433[3]), .I1(n552_adj_3646), 
            .CO(n38048));
    SB_CARRY mult_14_add_1219_4 (.CI(n38370), .I0(n8452[1]), .I1(n244_adj_3644), 
            .CO(n38371));
    SB_CARRY add_3178_8 (.CI(n37607), .I0(n10856[5]), .I1(n545), .CO(n37608));
    SB_LUT4 add_3105_5_lut (.I0(GND_net), .I1(n8433[2]), .I2(n455_adj_3647), 
            .I3(n38046), .O(n8422[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_9 (.CI(n37092), .I0(n13738[6]), .I1(GND_net), .CO(n37093));
    SB_CARRY add_22497_22 (.CI(n36761), .I0(n79[20]), .I1(n191[20]), .CO(n36762));
    SB_LUT4 add_3307_8_lut (.I0(GND_net), .I1(n13738[5]), .I2(n545), .I3(n37091), 
            .O(n13260[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_21_lut (.I0(GND_net), .I1(n79[19]), .I2(n191[19]), 
            .I3(n36760), .O(\PID_CONTROLLER.result_31__N_2994 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_5 (.CI(n38046), .I0(n8433[2]), .I1(n455_adj_3647), 
            .CO(n38047));
    SB_CARRY add_3307_8 (.CI(n37091), .I0(n13738[5]), .I1(n545), .CO(n37092));
    SB_LUT4 mult_14_add_1219_3_lut (.I0(GND_net), .I1(n8452[0]), .I2(n171_adj_3649), 
            .I3(n38369), .O(n1804[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_3 (.CI(n38369), .I0(n8452[0]), .I1(n171_adj_3649), 
            .CO(n38370));
    SB_LUT4 add_3105_4_lut (.I0(GND_net), .I1(n8433[1]), .I2(n358_adj_3650), 
            .I3(n38045), .O(n8422[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_7_lut (.I0(GND_net), .I1(n10856[4]), .I2(n472), .I3(n37606), 
            .O(n10122[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_7 (.CI(n37606), .I0(n10856[4]), .I1(n472), .CO(n37607));
    SB_CARRY add_3105_4 (.CI(n38045), .I0(n8433[1]), .I1(n358_adj_3650), 
            .CO(n38046));
    SB_LUT4 add_3178_6_lut (.I0(GND_net), .I1(n10856[3]), .I2(n399), .I3(n37605), 
            .O(n10122[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_6 (.CI(n37605), .I0(n10856[3]), .I1(n399), .CO(n37606));
    SB_LUT4 add_3178_5_lut (.I0(GND_net), .I1(n10856[2]), .I2(n326), .I3(n37604), 
            .O(n10122[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3307_7_lut (.I0(GND_net), .I1(n13738[4]), .I2(n472), .I3(n37090), 
            .O(n13260[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3105_3_lut (.I0(GND_net), .I1(n8433[0]), .I2(n261_adj_3651), 
            .I3(n38044), .O(n8422[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_5 (.CI(n37604), .I0(n10856[2]), .I1(n326), .CO(n37605));
    SB_CARRY add_3307_7 (.CI(n37090), .I0(n13738[4]), .I1(n472), .CO(n37091));
    SB_LUT4 add_3178_4_lut (.I0(GND_net), .I1(n10856[1]), .I2(n253), .I3(n37603), 
            .O(n10122[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3307_6_lut (.I0(GND_net), .I1(n13738[3]), .I2(n399), .I3(n37089), 
            .O(n13260[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n98_adj_3652), 
            .I3(GND_net), .O(n1804[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_3 (.CI(n38044), .I0(n8433[0]), .I1(n261_adj_3651), 
            .CO(n38045));
    SB_CARRY add_3178_4 (.CI(n37603), .I0(n10856[1]), .I1(n253), .CO(n37604));
    SB_CARRY add_3307_6 (.CI(n37089), .I0(n13738[3]), .I1(n399), .CO(n37090));
    SB_LUT4 add_3307_5_lut (.I0(GND_net), .I1(n13738[2]), .I2(n326), .I3(n37088), 
            .O(n13260[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_3_lut (.I0(GND_net), .I1(n10856[0]), .I2(n180_adj_3552), 
            .I3(n37602), .O(n10122[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_3 (.CI(n37602), .I0(n10856[0]), .I1(n180_adj_3552), 
            .CO(n37603));
    SB_CARRY add_3307_5 (.CI(n37088), .I0(n13738[2]), .I1(n326), .CO(n37089));
    SB_LUT4 add_3178_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n10122[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n98_adj_3652), 
            .CO(n38369));
    SB_LUT4 add_3105_2_lut (.I0(GND_net), .I1(n71_adj_3653), .I2(n164_adj_3654), 
            .I3(GND_net), .O(n8422[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n37602));
    SB_LUT4 add_3307_4_lut (.I0(GND_net), .I1(n13738[1]), .I2(n253), .I3(n37087), 
            .O(n13260[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_19_lut (.I0(GND_net), .I1(n11535[16]), .I2(GND_net), 
            .I3(n37601), .O(n10856[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_4 (.CI(n37087), .I0(n13738[1]), .I1(n253), .CO(n37088));
    SB_LUT4 add_3307_3_lut (.I0(GND_net), .I1(n13738[0]), .I2(n180_adj_3552), 
            .I3(n37086), .O(n13260[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_2 (.CI(GND_net), .I0(n71_adj_3653), .I1(n164_adj_3654), 
            .CO(n38044));
    SB_LUT4 add_3206_18_lut (.I0(GND_net), .I1(n11535[15]), .I2(GND_net), 
            .I3(n37600), .O(n10856[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_24_lut (.I0(GND_net), .I1(n1804[21]), .I2(GND_net), 
            .I3(n38367), .O(n1803[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_11_lut (.I0(GND_net), .I1(n8422[8]), .I2(GND_net), 
            .I3(n38043), .O(n8410[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_18 (.CI(n37600), .I0(n11535[15]), .I1(GND_net), 
            .CO(n37601));
    SB_LUT4 add_3206_17_lut (.I0(GND_net), .I1(n11535[14]), .I2(GND_net), 
            .I3(n37599), .O(n10856[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_21 (.CI(n36760), .I0(n79[19]), .I1(n191[19]), .CO(n36761));
    SB_LUT4 add_22497_20_lut (.I0(GND_net), .I1(n79[18]), .I2(n191[18]), 
            .I3(n36759), .O(\PID_CONTROLLER.result_31__N_2994 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_17 (.CI(n37599), .I0(n11535[14]), .I1(GND_net), 
            .CO(n37600));
    SB_CARRY add_3307_3 (.CI(n37086), .I0(n13738[0]), .I1(n180_adj_3552), 
            .CO(n37087));
    SB_LUT4 add_3307_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n13260[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_10_lut (.I0(GND_net), .I1(n8422[7]), .I2(GND_net), 
            .I3(n38042), .O(n8410[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_16_lut (.I0(GND_net), .I1(n11535[13]), .I2(GND_net), 
            .I3(n37598), .O(n10856[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n37086));
    SB_CARRY add_3206_16 (.CI(n37598), .I0(n11535[13]), .I1(GND_net), 
            .CO(n37599));
    SB_LUT4 add_3131_29_lut (.I0(GND_net), .I1(n9933[26]), .I2(GND_net), 
            .I3(n37085), .O(n9129[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_28_lut (.I0(GND_net), .I1(n9933[25]), .I2(GND_net), 
            .I3(n37084), .O(n9129[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_24 (.CI(n38367), .I0(n1804[21]), .I1(GND_net), 
            .CO(n1711));
    SB_CARRY add_3104_10 (.CI(n38042), .I0(n8422[7]), .I1(GND_net), .CO(n38043));
    SB_LUT4 add_3206_15_lut (.I0(GND_net), .I1(n11535[12]), .I2(GND_net), 
            .I3(n37597), .O(n10856[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_28 (.CI(n37084), .I0(n9933[25]), .I1(GND_net), .CO(n37085));
    SB_CARRY add_3206_15 (.CI(n37597), .I0(n11535[12]), .I1(GND_net), 
            .CO(n37598));
    SB_LUT4 add_3131_27_lut (.I0(GND_net), .I1(n9933[24]), .I2(GND_net), 
            .I3(n37083), .O(n9129[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_27 (.CI(n37083), .I0(n9933[24]), .I1(GND_net), .CO(n37084));
    SB_LUT4 add_3104_9_lut (.I0(GND_net), .I1(n8422[6]), .I2(GND_net), 
            .I3(n38041), .O(n8410[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_14_lut (.I0(GND_net), .I1(n11535[11]), .I2(GND_net), 
            .I3(n37596), .O(n10856[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_26_lut (.I0(GND_net), .I1(n9933[23]), .I2(GND_net), 
            .I3(n37082), .O(n9129[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_23_lut (.I0(GND_net), .I1(n1804[20]), .I2(GND_net), 
            .I3(n38366), .O(n1803[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3104_9 (.CI(n38041), .I0(n8422[6]), .I1(GND_net), .CO(n38042));
    SB_CARRY add_3206_14 (.CI(n37596), .I0(n11535[11]), .I1(GND_net), 
            .CO(n37597));
    SB_CARRY add_3131_26 (.CI(n37082), .I0(n9933[23]), .I1(GND_net), .CO(n37083));
    SB_LUT4 add_3131_25_lut (.I0(GND_net), .I1(n9933[22]), .I2(GND_net), 
            .I3(n37081), .O(n9129[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_8_lut (.I0(GND_net), .I1(n8422[5]), .I2(n743_adj_3655), 
            .I3(n38040), .O(n8410[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_13_lut (.I0(GND_net), .I1(n11535[10]), .I2(GND_net), 
            .I3(n37595), .O(n10856[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_25 (.CI(n37081), .I0(n9933[22]), .I1(GND_net), .CO(n37082));
    SB_CARRY add_22497_20 (.CI(n36759), .I0(n79[18]), .I1(n191[18]), .CO(n36760));
    SB_LUT4 add_3131_24_lut (.I0(GND_net), .I1(n9933[21]), .I2(GND_net), 
            .I3(n37080), .O(n9129[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_19_lut (.I0(GND_net), .I1(n79[17]), .I2(n191[17]), 
            .I3(n36758), .O(\PID_CONTROLLER.result_31__N_2994 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_23 (.CI(n38366), .I0(n1804[20]), .I1(GND_net), 
            .CO(n38367));
    SB_CARRY add_3104_8 (.CI(n38040), .I0(n8422[5]), .I1(n743_adj_3655), 
            .CO(n38041));
    SB_CARRY add_3206_13 (.CI(n37595), .I0(n11535[10]), .I1(GND_net), 
            .CO(n37596));
    SB_CARRY add_3131_24 (.CI(n37080), .I0(n9933[21]), .I1(GND_net), .CO(n37081));
    SB_LUT4 add_3131_23_lut (.I0(GND_net), .I1(n9933[20]), .I2(GND_net), 
            .I3(n37079), .O(n9129[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_7_lut (.I0(GND_net), .I1(n8422[4]), .I2(n646_adj_3656), 
            .I3(n38039), .O(n8410[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_12_lut (.I0(GND_net), .I1(n11535[9]), .I2(GND_net), 
            .I3(n37594), .O(n10856[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_23 (.CI(n37079), .I0(n9933[20]), .I1(GND_net), .CO(n37080));
    SB_CARRY add_22497_19 (.CI(n36758), .I0(n79[17]), .I1(n191[17]), .CO(n36759));
    SB_LUT4 add_3131_22_lut (.I0(GND_net), .I1(n9933[19]), .I2(GND_net), 
            .I3(n37078), .O(n9129[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_18_lut (.I0(GND_net), .I1(n79[16]), .I2(n191[16]), 
            .I3(n36757), .O(\PID_CONTROLLER.result_31__N_2994 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_22_lut (.I0(GND_net), .I1(n1804[19]), .I2(GND_net), 
            .I3(n38365), .O(n1803[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3104_7 (.CI(n38039), .I0(n8422[4]), .I1(n646_adj_3656), 
            .CO(n38040));
    SB_CARRY add_3206_12 (.CI(n37594), .I0(n11535[9]), .I1(GND_net), .CO(n37595));
    SB_CARRY add_3131_22 (.CI(n37078), .I0(n9933[19]), .I1(GND_net), .CO(n37079));
    SB_LUT4 add_3131_21_lut (.I0(GND_net), .I1(n9933[18]), .I2(GND_net), 
            .I3(n37077), .O(n9129[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_6_lut (.I0(GND_net), .I1(n8422[3]), .I2(n549_adj_3657), 
            .I3(n38038), .O(n8410[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_11_lut (.I0(GND_net), .I1(n11535[8]), .I2(GND_net), 
            .I3(n37593), .O(n10856[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_21 (.CI(n37077), .I0(n9933[18]), .I1(GND_net), .CO(n37078));
    SB_CARRY add_22497_18 (.CI(n36757), .I0(n79[16]), .I1(n191[16]), .CO(n36758));
    SB_LUT4 add_3131_20_lut (.I0(GND_net), .I1(n9933[17]), .I2(GND_net), 
            .I3(n37076), .O(n9129[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_17_lut (.I0(GND_net), .I1(n79[15]), .I2(n191[15]), 
            .I3(n36756), .O(\PID_CONTROLLER.result_31__N_2994 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_22 (.CI(n38365), .I0(n1804[19]), .I1(GND_net), 
            .CO(n38366));
    SB_CARRY add_3104_6 (.CI(n38038), .I0(n8422[3]), .I1(n549_adj_3657), 
            .CO(n38039));
    SB_CARRY add_3206_11 (.CI(n37593), .I0(n11535[8]), .I1(GND_net), .CO(n37594));
    SB_CARRY add_3131_20 (.CI(n37076), .I0(n9933[17]), .I1(GND_net), .CO(n37077));
    SB_LUT4 add_3131_19_lut (.I0(GND_net), .I1(n9933[16]), .I2(GND_net), 
            .I3(n37075), .O(n9129[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_5_lut (.I0(GND_net), .I1(n8422[2]), .I2(n452_adj_3658), 
            .I3(n38037), .O(n8410[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_10_lut (.I0(GND_net), .I1(n11535[7]), .I2(GND_net), 
            .I3(n37592), .O(n10856[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_19 (.CI(n37075), .I0(n9933[16]), .I1(GND_net), .CO(n37076));
    SB_CARRY add_22497_17 (.CI(n36756), .I0(n79[15]), .I1(n191[15]), .CO(n36757));
    SB_LUT4 add_3131_18_lut (.I0(GND_net), .I1(n9933[15]), .I2(GND_net), 
            .I3(n37074), .O(n9129[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_16_lut (.I0(GND_net), .I1(n79[14]), .I2(n191[14]), 
            .I3(n36755), .O(\PID_CONTROLLER.result_31__N_2994 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1218_21_lut (.I0(GND_net), .I1(n1804[18]), .I2(GND_net), 
            .I3(n38364), .O(n1803[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3104_5 (.CI(n38037), .I0(n8422[2]), .I1(n452_adj_3658), 
            .CO(n38038));
    SB_LUT4 mult_14_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3422));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i6_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3206_10 (.CI(n37592), .I0(n11535[7]), .I1(GND_net), .CO(n37593));
    SB_LUT4 add_3206_9_lut (.I0(GND_net), .I1(n11535[6]), .I2(GND_net), 
            .I3(n37591), .O(n10856[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_18 (.CI(n37074), .I0(n9933[15]), .I1(GND_net), .CO(n37075));
    SB_LUT4 add_3131_17_lut (.I0(GND_net), .I1(n9933[14]), .I2(GND_net), 
            .I3(n37073), .O(n9129[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_21 (.CI(n38364), .I0(n1804[18]), .I1(GND_net), 
            .CO(n38365));
    SB_LUT4 add_3104_4_lut (.I0(GND_net), .I1(n8422[1]), .I2(n355_adj_3659), 
            .I3(n38036), .O(n8410[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_9 (.CI(n37591), .I0(n11535[6]), .I1(GND_net), .CO(n37592));
    SB_CARRY add_3131_17 (.CI(n37073), .I0(n9933[14]), .I1(GND_net), .CO(n37074));
    SB_LUT4 add_3206_8_lut (.I0(GND_net), .I1(n11535[5]), .I2(n545), .I3(n37590), 
            .O(n10856[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_16_lut (.I0(GND_net), .I1(n9933[13]), .I2(GND_net), 
            .I3(n37072), .O(n9129[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_16 (.CI(n37072), .I0(n9933[13]), .I1(GND_net), .CO(n37073));
    SB_CARRY add_3104_4 (.CI(n38036), .I0(n8422[1]), .I1(n355_adj_3659), 
            .CO(n38037));
    SB_CARRY add_3206_8 (.CI(n37590), .I0(n11535[5]), .I1(n545), .CO(n37591));
    SB_LUT4 add_3131_15_lut (.I0(GND_net), .I1(n9933[12]), .I2(GND_net), 
            .I3(n37071), .O(n9129[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_7_lut (.I0(GND_net), .I1(n11535[4]), .I2(n472), .I3(n37589), 
            .O(n10856[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_15 (.CI(n37071), .I0(n9933[12]), .I1(GND_net), .CO(n37072));
    SB_LUT4 add_3131_14_lut (.I0(GND_net), .I1(n9933[11]), .I2(GND_net), 
            .I3(n37070), .O(n9129[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_20_lut (.I0(GND_net), .I1(n1804[17]), .I2(GND_net), 
            .I3(n38363), .O(n1803[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_3_lut (.I0(GND_net), .I1(n8422[0]), .I2(n258_adj_3660), 
            .I3(n38035), .O(n8410[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_7 (.CI(n37589), .I0(n11535[4]), .I1(n472), .CO(n37590));
    SB_LUT4 add_3206_6_lut (.I0(GND_net), .I1(n11535[3]), .I2(n399), .I3(n37588), 
            .O(n10856[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_14 (.CI(n37070), .I0(n9933[11]), .I1(GND_net), .CO(n37071));
    SB_DFFE \PID_CONTROLLER.integral_1049__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[0]));   // verilog/motorControl.v(34[21:33])
    SB_LUT4 add_3131_13_lut (.I0(GND_net), .I1(n9933[10]), .I2(GND_net), 
            .I3(n37069), .O(n9129[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_6 (.CI(n37588), .I0(n11535[3]), .I1(n399), .CO(n37589));
    SB_CARRY add_3104_3 (.CI(n38035), .I0(n8422[0]), .I1(n258_adj_3660), 
            .CO(n38036));
    SB_LUT4 add_3206_5_lut (.I0(GND_net), .I1(n11535[2]), .I2(n326), .I3(n37587), 
            .O(n10856[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_13 (.CI(n37069), .I0(n9933[10]), .I1(GND_net), .CO(n37070));
    SB_CARRY mult_14_add_1218_20 (.CI(n38363), .I0(n1804[17]), .I1(GND_net), 
            .CO(n38364));
    SB_LUT4 add_3131_12_lut (.I0(GND_net), .I1(n9933[9]), .I2(GND_net), 
            .I3(n37068), .O(n9129[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_19_lut (.I0(GND_net), .I1(n1804[16]), .I2(GND_net), 
            .I3(n38362), .O(n1803[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_5 (.CI(n37587), .I0(n11535[2]), .I1(n326), .CO(n37588));
    SB_LUT4 add_3104_2_lut (.I0(GND_net), .I1(n68_adj_3662), .I2(n161_adj_3663), 
            .I3(GND_net), .O(n8410[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_4_lut (.I0(GND_net), .I1(n11535[1]), .I2(n253), .I3(n37586), 
            .O(n10856[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_12 (.CI(n37068), .I0(n9933[9]), .I1(GND_net), .CO(n37069));
    SB_CARRY mult_14_add_1218_19 (.CI(n38362), .I0(n1804[16]), .I1(GND_net), 
            .CO(n38363));
    SB_CARRY add_3104_2 (.CI(GND_net), .I0(n68_adj_3662), .I1(n161_adj_3663), 
            .CO(n38035));
    SB_LUT4 add_3103_12_lut (.I0(GND_net), .I1(n8410[9]), .I2(GND_net), 
            .I3(n38034), .O(n8397[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_4 (.CI(n37586), .I0(n11535[1]), .I1(n253), .CO(n37587));
    SB_LUT4 add_3131_11_lut (.I0(GND_net), .I1(n9933[8]), .I2(GND_net), 
            .I3(n37067), .O(n9129[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_3_lut (.I0(GND_net), .I1(n11535[0]), .I2(n180_adj_3552), 
            .I3(n37585), .O(n10856[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_3 (.CI(n37585), .I0(n11535[0]), .I1(n180_adj_3552), 
            .CO(n37586));
    SB_CARRY add_3131_11 (.CI(n37067), .I0(n9933[8]), .I1(GND_net), .CO(n37068));
    SB_LUT4 add_3131_10_lut (.I0(GND_net), .I1(n9933[7]), .I2(GND_net), 
            .I3(n37066), .O(n9129[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_11_lut (.I0(GND_net), .I1(n8410[8]), .I2(GND_net), 
            .I3(n38033), .O(n8397[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n10856[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_10 (.CI(n37066), .I0(n9933[7]), .I1(GND_net), .CO(n37067));
    SB_CARRY add_3206_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n37585));
    SB_LUT4 add_3131_9_lut (.I0(GND_net), .I1(n9933[6]), .I2(GND_net), 
            .I3(n37065), .O(n9129[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_9 (.CI(n37065), .I0(n9933[6]), .I1(GND_net), .CO(n37066));
    SB_LUT4 mult_14_add_1218_18_lut (.I0(GND_net), .I1(n1804[15]), .I2(GND_net), 
            .I3(n38361), .O(n1803[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_8_lut (.I0(GND_net), .I1(n9933[5]), .I2(n689_adj_3664), 
            .I3(n37064), .O(n9129[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_18_lut (.I0(GND_net), .I1(n12161[15]), .I2(GND_net), 
            .I3(n37584), .O(n11535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_11 (.CI(n38033), .I0(n8410[8]), .I1(GND_net), .CO(n38034));
    SB_CARRY add_22497_16 (.CI(n36755), .I0(n79[14]), .I1(n191[14]), .CO(n36756));
    SB_LUT4 add_22497_15_lut (.I0(GND_net), .I1(n79[13]), .I2(n191[13]), 
            .I3(n36754), .O(\PID_CONTROLLER.result_31__N_2994 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_17_lut (.I0(GND_net), .I1(n12161[14]), .I2(GND_net), 
            .I3(n37583), .O(n11535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_8 (.CI(n37064), .I0(n9933[5]), .I1(n689_adj_3664), 
            .CO(n37065));
    SB_CARRY add_3233_17 (.CI(n37583), .I0(n12161[14]), .I1(GND_net), 
            .CO(n37584));
    SB_LUT4 add_3131_7_lut (.I0(GND_net), .I1(n9933[4]), .I2(n592_adj_3665), 
            .I3(n37063), .O(n9129[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_7 (.CI(n37063), .I0(n9933[4]), .I1(n592_adj_3665), 
            .CO(n37064));
    SB_LUT4 add_3103_10_lut (.I0(GND_net), .I1(n8410[7]), .I2(GND_net), 
            .I3(n38032), .O(n8397[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_16_lut (.I0(GND_net), .I1(n12161[13]), .I2(GND_net), 
            .I3(n37582), .O(n11535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_6_lut (.I0(GND_net), .I1(n9933[3]), .I2(n495_adj_3666), 
            .I3(n37062), .O(n9129[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_10 (.CI(n38032), .I0(n8410[7]), .I1(GND_net), .CO(n38033));
    SB_LUT4 add_3103_9_lut (.I0(GND_net), .I1(n8410[6]), .I2(GND_net), 
            .I3(n38031), .O(n8397[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_16 (.CI(n37582), .I0(n12161[13]), .I1(GND_net), 
            .CO(n37583));
    SB_CARRY add_3131_6 (.CI(n37062), .I0(n9933[3]), .I1(n495_adj_3666), 
            .CO(n37063));
    SB_LUT4 add_3233_15_lut (.I0(GND_net), .I1(n12161[12]), .I2(GND_net), 
            .I3(n37581), .O(n11535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_5_lut (.I0(GND_net), .I1(n9933[2]), .I2(n398_adj_3667), 
            .I3(n37061), .O(n9129[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_5 (.CI(n37061), .I0(n9933[2]), .I1(n398_adj_3667), 
            .CO(n37062));
    SB_CARRY mult_14_add_1218_18 (.CI(n38361), .I0(n1804[15]), .I1(GND_net), 
            .CO(n38362));
    SB_CARRY add_3103_9 (.CI(n38031), .I0(n8410[6]), .I1(GND_net), .CO(n38032));
    SB_CARRY add_3233_15 (.CI(n37581), .I0(n12161[12]), .I1(GND_net), 
            .CO(n37582));
    SB_LUT4 add_3131_4_lut (.I0(GND_net), .I1(n9933[1]), .I2(n301_adj_3668), 
            .I3(n37060), .O(n9129[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_14_lut (.I0(GND_net), .I1(n12161[11]), .I2(GND_net), 
            .I3(n37580), .O(n11535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_4 (.CI(n37060), .I0(n9933[1]), .I1(n301_adj_3668), 
            .CO(n37061));
    SB_LUT4 add_3131_3_lut (.I0(GND_net), .I1(n9933[0]), .I2(n204_adj_3669), 
            .I3(n37059), .O(n9129[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_8_lut (.I0(GND_net), .I1(n8410[5]), .I2(n740_adj_3670), 
            .I3(n38030), .O(n8397[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_14 (.CI(n37580), .I0(n12161[11]), .I1(GND_net), 
            .CO(n37581));
    SB_LUT4 add_3233_13_lut (.I0(GND_net), .I1(n12161[10]), .I2(GND_net), 
            .I3(n37579), .O(n11535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_3 (.CI(n37059), .I0(n9933[0]), .I1(n204_adj_3669), 
            .CO(n37060));
    SB_LUT4 add_3131_2_lut (.I0(GND_net), .I1(n14_adj_3671), .I2(n107_adj_3672), 
            .I3(GND_net), .O(n9129[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_15 (.CI(n36754), .I0(n79[13]), .I1(n191[13]), .CO(n36755));
    SB_LUT4 add_22497_14_lut (.I0(GND_net), .I1(n79[12]), .I2(n191[12]), 
            .I3(n36753), .O(\PID_CONTROLLER.result_31__N_2994 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_13 (.CI(n37579), .I0(n12161[10]), .I1(GND_net), 
            .CO(n37580));
    SB_LUT4 add_3233_12_lut (.I0(GND_net), .I1(n12161[9]), .I2(GND_net), 
            .I3(n37578), .O(n11535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_2 (.CI(GND_net), .I0(n14_adj_3671), .I1(n107_adj_3672), 
            .CO(n37059));
    SB_LUT4 add_3329_14_lut (.I0(GND_net), .I1(n14172[11]), .I2(GND_net), 
            .I3(n37058), .O(n13738[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_17_lut (.I0(GND_net), .I1(n1804[14]), .I2(GND_net), 
            .I3(n38360), .O(n1803[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_12 (.CI(n37578), .I0(n12161[9]), .I1(GND_net), .CO(n37579));
    SB_LUT4 add_3329_13_lut (.I0(GND_net), .I1(n14172[10]), .I2(GND_net), 
            .I3(n37057), .O(n13738[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_13 (.CI(n37057), .I0(n14172[10]), .I1(GND_net), 
            .CO(n37058));
    SB_CARRY add_22497_14 (.CI(n36753), .I0(n79[12]), .I1(n191[12]), .CO(n36754));
    SB_CARRY mult_14_add_1218_17 (.CI(n38360), .I0(n1804[14]), .I1(GND_net), 
            .CO(n38361));
    SB_CARRY add_3103_8 (.CI(n38030), .I0(n8410[5]), .I1(n740_adj_3670), 
            .CO(n38031));
    SB_LUT4 add_3329_12_lut (.I0(GND_net), .I1(n14172[9]), .I2(GND_net), 
            .I3(n37056), .O(n13738[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_12 (.CI(n37056), .I0(n14172[9]), .I1(GND_net), .CO(n37057));
    SB_LUT4 add_3233_11_lut (.I0(GND_net), .I1(n12161[8]), .I2(GND_net), 
            .I3(n37577), .O(n11535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_13_lut (.I0(GND_net), .I1(n79[11]), .I2(n191[11]), 
            .I3(n36752), .O(\PID_CONTROLLER.result_31__N_2994 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_13 (.CI(n36752), .I0(n79[11]), .I1(n191[11]), .CO(n36753));
    SB_CARRY add_3233_11 (.CI(n37577), .I0(n12161[8]), .I1(GND_net), .CO(n37578));
    SB_LUT4 add_3329_11_lut (.I0(GND_net), .I1(n14172[8]), .I2(GND_net), 
            .I3(n37055), .O(n13738[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_7_lut (.I0(GND_net), .I1(n8410[4]), .I2(n643_adj_3673), 
            .I3(n38029), .O(n8397[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_16_lut (.I0(GND_net), .I1(n1804[13]), .I2(GND_net), 
            .I3(n38359), .O(n1803[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_7 (.CI(n38029), .I0(n8410[4]), .I1(n643_adj_3673), 
            .CO(n38030));
    SB_CARRY add_3329_11 (.CI(n37055), .I0(n14172[8]), .I1(GND_net), .CO(n37056));
    SB_LUT4 add_3233_10_lut (.I0(GND_net), .I1(n12161[7]), .I2(GND_net), 
            .I3(n37576), .O(n11535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3329_10_lut (.I0(GND_net), .I1(n14172[7]), .I2(GND_net), 
            .I3(n37054), .O(n13738[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_10 (.CI(n37054), .I0(n14172[7]), .I1(GND_net), .CO(n37055));
    SB_LUT4 add_22497_12_lut (.I0(GND_net), .I1(n79[10]), .I2(n191[10]), 
            .I3(n36751), .O(\PID_CONTROLLER.result_31__N_2994 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_12 (.CI(n36751), .I0(n79[10]), .I1(n191[10]), .CO(n36752));
    SB_CARRY add_3233_10 (.CI(n37576), .I0(n12161[7]), .I1(GND_net), .CO(n37577));
    SB_LUT4 add_3233_9_lut (.I0(GND_net), .I1(n12161[6]), .I2(GND_net), 
            .I3(n37575), .O(n11535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_9 (.CI(n37575), .I0(n12161[6]), .I1(GND_net), .CO(n37576));
    SB_LUT4 add_3329_9_lut (.I0(GND_net), .I1(n14172[6]), .I2(GND_net), 
            .I3(n37053), .O(n13738[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_6_lut (.I0(GND_net), .I1(n8410[3]), .I2(n546_adj_3674), 
            .I3(n38028), .O(n8397[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_9 (.CI(n37053), .I0(n14172[6]), .I1(GND_net), .CO(n37054));
    SB_LUT4 add_3233_8_lut (.I0(GND_net), .I1(n12161[5]), .I2(n545), .I3(n37574), 
            .O(n11535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_6 (.CI(n38028), .I0(n8410[3]), .I1(n546_adj_3674), 
            .CO(n38029));
    SB_CARRY add_3233_8 (.CI(n37574), .I0(n12161[5]), .I1(n545), .CO(n37575));
    SB_LUT4 add_3329_8_lut (.I0(GND_net), .I1(n14172[5]), .I2(n545), .I3(n37052), 
            .O(n13738[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_16 (.CI(n38359), .I0(n1804[13]), .I1(GND_net), 
            .CO(n38360));
    SB_LUT4 add_22497_11_lut (.I0(GND_net), .I1(n79[9]), .I2(n191[9]), 
            .I3(n36750), .O(\PID_CONTROLLER.result_31__N_2994 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_5_lut (.I0(GND_net), .I1(n8410[2]), .I2(n449_adj_3675), 
            .I3(n38027), .O(n8397[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_15_lut (.I0(GND_net), .I1(n1804[12]), .I2(GND_net), 
            .I3(n38358), .O(n1803[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_7_lut (.I0(GND_net), .I1(n12161[4]), .I2(n472), .I3(n37573), 
            .O(n11535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_7 (.CI(n37573), .I0(n12161[4]), .I1(n472), .CO(n37574));
    SB_LUT4 add_3233_6_lut (.I0(GND_net), .I1(n12161[3]), .I2(n399), .I3(n37572), 
            .O(n11535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_8 (.CI(n37052), .I0(n14172[5]), .I1(n545), .CO(n37053));
    SB_LUT4 add_3329_7_lut (.I0(GND_net), .I1(n14172[4]), .I2(n472), .I3(n37051), 
            .O(n13738[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_11 (.CI(n36750), .I0(n79[9]), .I1(n191[9]), .CO(n36751));
    SB_CARRY add_3103_5 (.CI(n38027), .I0(n8410[2]), .I1(n449_adj_3675), 
            .CO(n38028));
    SB_CARRY add_3233_6 (.CI(n37572), .I0(n12161[3]), .I1(n399), .CO(n37573));
    SB_LUT4 add_3103_4_lut (.I0(GND_net), .I1(n8410[1]), .I2(n352_adj_3676), 
            .I3(n38026), .O(n8397[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_5_lut (.I0(GND_net), .I1(n12161[2]), .I2(n326), .I3(n37571), 
            .O(n11535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_10_lut (.I0(GND_net), .I1(n79[8]), .I2(n191[8]), 
            .I3(n36749), .O(\PID_CONTROLLER.result_31__N_2994 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_4 (.CI(n38026), .I0(n8410[1]), .I1(n352_adj_3676), 
            .CO(n38027));
    SB_CARRY add_3233_5 (.CI(n37571), .I0(n12161[2]), .I1(n326), .CO(n37572));
    SB_LUT4 add_3233_4_lut (.I0(GND_net), .I1(n12161[1]), .I2(n253), .I3(n37570), 
            .O(n11535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_7 (.CI(n37051), .I0(n14172[4]), .I1(n472), .CO(n37052));
    SB_LUT4 add_3329_6_lut (.I0(GND_net), .I1(n14172[3]), .I2(n399), .I3(n37050), 
            .O(n13738[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_10 (.CI(n36749), .I0(n79[8]), .I1(n191[8]), .CO(n36750));
    SB_LUT4 add_3103_3_lut (.I0(GND_net), .I1(n8410[0]), .I2(n255_adj_3677), 
            .I3(n38025), .O(n8397[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_15 (.CI(n38358), .I0(n1804[12]), .I1(GND_net), 
            .CO(n38359));
    SB_CARRY add_3233_4 (.CI(n37570), .I0(n12161[1]), .I1(n253), .CO(n37571));
    SB_LUT4 add_22497_9_lut (.I0(GND_net), .I1(n79[7]), .I2(n191[7]), 
            .I3(n36748), .O(\PID_CONTROLLER.result_31__N_2994 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_3 (.CI(n38025), .I0(n8410[0]), .I1(n255_adj_3677), 
            .CO(n38026));
    SB_LUT4 add_3233_3_lut (.I0(GND_net), .I1(n12161[0]), .I2(n180_adj_3552), 
            .I3(n37569), .O(n11535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_14_lut (.I0(GND_net), .I1(n1804[11]), .I2(GND_net), 
            .I3(n38357), .O(n1803[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_6 (.CI(n37050), .I0(n14172[3]), .I1(n399), .CO(n37051));
    SB_LUT4 add_3103_2_lut (.I0(GND_net), .I1(n65_adj_3678), .I2(n158_adj_3679), 
            .I3(GND_net), .O(n8397[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3329_5_lut (.I0(GND_net), .I1(n14172[2]), .I2(n326), .I3(n37049), 
            .O(n13738[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_3 (.CI(n37569), .I0(n12161[0]), .I1(n180_adj_3552), 
            .CO(n37570));
    SB_LUT4 add_3233_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n11535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n37569));
    SB_CARRY add_3329_5 (.CI(n37049), .I0(n14172[2]), .I1(n326), .CO(n37050));
    SB_CARRY mult_14_add_1218_14 (.CI(n38357), .I0(n1804[11]), .I1(GND_net), 
            .CO(n38358));
    SB_LUT4 add_3329_4_lut (.I0(GND_net), .I1(n14172[1]), .I2(n253), .I3(n37048), 
            .O(n13738[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_4 (.CI(n37048), .I0(n14172[1]), .I1(n253), .CO(n37049));
    SB_LUT4 add_3329_3_lut (.I0(GND_net), .I1(n14172[0]), .I2(n180_adj_3552), 
            .I3(n37047), .O(n13738[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_9 (.CI(n36748), .I0(n79[7]), .I1(n191[7]), .CO(n36749));
    SB_CARRY add_3329_3 (.CI(n37047), .I0(n14172[0]), .I1(n180_adj_3552), 
            .CO(n37048));
    SB_LUT4 add_3329_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n13738[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_2 (.CI(GND_net), .I0(n65_adj_3678), .I1(n158_adj_3679), 
            .CO(n38025));
    SB_LUT4 add_3259_17_lut (.I0(GND_net), .I1(n12736[14]), .I2(GND_net), 
            .I3(n37568), .O(n12161[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n37047));
    SB_LUT4 add_3102_13_lut (.I0(GND_net), .I1(n8397[10]), .I2(GND_net), 
            .I3(n38024), .O(n8383[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_16_lut (.I0(GND_net), .I1(n12736[13]), .I2(GND_net), 
            .I3(n37567), .O(n12161[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_28_lut (.I0(GND_net), .I1(n10675[25]), .I2(GND_net), 
            .I3(n37046), .O(n9933[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_8_lut (.I0(GND_net), .I1(n79[6]), .I2(n191[6]), 
            .I3(n36747), .O(\PID_CONTROLLER.result_31__N_2994 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_27_lut (.I0(GND_net), .I1(n10675[24]), .I2(GND_net), 
            .I3(n37045), .O(n9933[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_8 (.CI(n36747), .I0(n79[6]), .I1(n191[6]), .CO(n36748));
    SB_CARRY add_3170_27 (.CI(n37045), .I0(n10675[24]), .I1(GND_net), 
            .CO(n37046));
    SB_CARRY add_3259_16 (.CI(n37567), .I0(n12736[13]), .I1(GND_net), 
            .CO(n37568));
    SB_LUT4 add_22497_7_lut (.I0(GND_net), .I1(n79[5]), .I2(n191[5]), 
            .I3(n36746), .O(\PID_CONTROLLER.result_31__N_2994 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_13_lut (.I0(GND_net), .I1(n1804[10]), .I2(GND_net), 
            .I3(n38356), .O(n1803[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_7 (.CI(n36746), .I0(n79[5]), .I1(n191[5]), .CO(n36747));
    SB_LUT4 add_3259_15_lut (.I0(GND_net), .I1(n12736[12]), .I2(GND_net), 
            .I3(n37566), .O(n12161[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_6_lut (.I0(GND_net), .I1(n79[4]), .I2(n191[4]), 
            .I3(n36745), .O(\PID_CONTROLLER.result_31__N_2994 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3102_12_lut (.I0(GND_net), .I1(n8397[9]), .I2(GND_net), 
            .I3(n38023), .O(n8383[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_15 (.CI(n37566), .I0(n12736[12]), .I1(GND_net), 
            .CO(n37567));
    SB_LUT4 add_3170_26_lut (.I0(GND_net), .I1(n10675[23]), .I2(GND_net), 
            .I3(n37044), .O(n9933[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_26 (.CI(n37044), .I0(n10675[23]), .I1(GND_net), 
            .CO(n37045));
    SB_LUT4 add_3259_14_lut (.I0(GND_net), .I1(n12736[11]), .I2(GND_net), 
            .I3(n37565), .O(n12161[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_25_lut (.I0(GND_net), .I1(n10675[22]), .I2(GND_net), 
            .I3(n37043), .O(n9933[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_25 (.CI(n37043), .I0(n10675[22]), .I1(GND_net), 
            .CO(n37044));
    SB_CARRY add_3102_12 (.CI(n38023), .I0(n8397[9]), .I1(GND_net), .CO(n38024));
    SB_LUT4 add_3170_24_lut (.I0(GND_net), .I1(n10675[21]), .I2(GND_net), 
            .I3(n37042), .O(n9933[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_14 (.CI(n37565), .I0(n12736[11]), .I1(GND_net), 
            .CO(n37566));
    SB_LUT4 add_3102_11_lut (.I0(GND_net), .I1(n8397[8]), .I2(GND_net), 
            .I3(n38022), .O(n8383[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_24 (.CI(n37042), .I0(n10675[21]), .I1(GND_net), 
            .CO(n37043));
    SB_CARRY add_22497_6 (.CI(n36745), .I0(n79[4]), .I1(n191[4]), .CO(n36746));
    SB_CARRY mult_14_add_1218_13 (.CI(n38356), .I0(n1804[10]), .I1(GND_net), 
            .CO(n38357));
    SB_LUT4 add_3259_13_lut (.I0(GND_net), .I1(n12736[10]), .I2(GND_net), 
            .I3(n37564), .O(n12161[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_23_lut (.I0(GND_net), .I1(n10675[20]), .I2(GND_net), 
            .I3(n37041), .O(n9933[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_5_lut (.I0(GND_net), .I1(n79[3]), .I2(n191[3]), 
            .I3(n36744), .O(\PID_CONTROLLER.result_31__N_2994 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_11 (.CI(n38022), .I0(n8397[8]), .I1(GND_net), .CO(n38023));
    SB_LUT4 mult_14_add_1218_12_lut (.I0(GND_net), .I1(n1804[9]), .I2(GND_net), 
            .I3(n38355), .O(n1803[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_13 (.CI(n37564), .I0(n12736[10]), .I1(GND_net), 
            .CO(n37565));
    SB_CARRY add_3170_23 (.CI(n37041), .I0(n10675[20]), .I1(GND_net), 
            .CO(n37042));
    SB_LUT4 add_3102_10_lut (.I0(GND_net), .I1(n8397[7]), .I2(GND_net), 
            .I3(n38021), .O(n8383[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_12_lut (.I0(GND_net), .I1(n12736[9]), .I2(GND_net), 
            .I3(n37563), .O(n12161[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_22_lut (.I0(GND_net), .I1(n10675[19]), .I2(GND_net), 
            .I3(n37040), .O(n9933[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_22 (.CI(n37040), .I0(n10675[19]), .I1(GND_net), 
            .CO(n37041));
    SB_CARRY add_3259_12 (.CI(n37563), .I0(n12736[9]), .I1(GND_net), .CO(n37564));
    SB_CARRY add_3102_10 (.CI(n38021), .I0(n8397[7]), .I1(GND_net), .CO(n38022));
    SB_LUT4 add_3170_21_lut (.I0(GND_net), .I1(n10675[18]), .I2(GND_net), 
            .I3(n37039), .O(n9933[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_11_lut (.I0(GND_net), .I1(n12736[8]), .I2(GND_net), 
            .I3(n37562), .O(n12161[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_21 (.CI(n37039), .I0(n10675[18]), .I1(GND_net), 
            .CO(n37040));
    SB_LUT4 add_3170_20_lut (.I0(GND_net), .I1(n10675[17]), .I2(GND_net), 
            .I3(n37038), .O(n9933[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_11 (.CI(n37562), .I0(n12736[8]), .I1(GND_net), .CO(n37563));
    SB_CARRY add_3170_20 (.CI(n37038), .I0(n10675[17]), .I1(GND_net), 
            .CO(n37039));
    SB_LUT4 add_3102_9_lut (.I0(GND_net), .I1(n8397[6]), .I2(GND_net), 
            .I3(n38020), .O(n8383[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_19_lut (.I0(GND_net), .I1(n10675[16]), .I2(GND_net), 
            .I3(n37037), .O(n9933[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_12 (.CI(n38355), .I0(n1804[9]), .I1(GND_net), 
            .CO(n38356));
    SB_LUT4 add_3259_10_lut (.I0(GND_net), .I1(n12736[7]), .I2(GND_net), 
            .I3(n37561), .O(n12161[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_9 (.CI(n38020), .I0(n8397[6]), .I1(GND_net), .CO(n38021));
    SB_CARRY add_3170_19 (.CI(n37037), .I0(n10675[16]), .I1(GND_net), 
            .CO(n37038));
    SB_CARRY add_3259_10 (.CI(n37561), .I0(n12736[7]), .I1(GND_net), .CO(n37562));
    SB_LUT4 add_3170_18_lut (.I0(GND_net), .I1(n10675[15]), .I2(GND_net), 
            .I3(n37036), .O(n9933[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_9_lut (.I0(GND_net), .I1(n12736[6]), .I2(GND_net), 
            .I3(n37560), .O(n12161[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_5 (.CI(n36744), .I0(n79[3]), .I1(n191[3]), .CO(n36745));
    SB_CARRY add_3170_18 (.CI(n37036), .I0(n10675[15]), .I1(GND_net), 
            .CO(n37037));
    SB_CARRY add_3259_9 (.CI(n37560), .I0(n12736[6]), .I1(GND_net), .CO(n37561));
    SB_LUT4 add_3102_8_lut (.I0(GND_net), .I1(n8397[5]), .I2(n737_adj_3680), 
            .I3(n38019), .O(n8383[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_8 (.CI(n38019), .I0(n8397[5]), .I1(n737_adj_3680), 
            .CO(n38020));
    SB_LUT4 add_3259_8_lut (.I0(GND_net), .I1(n12736[5]), .I2(n545), .I3(n37559), 
            .O(n12161[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_8 (.CI(n37559), .I0(n12736[5]), .I1(n545), .CO(n37560));
    SB_LUT4 add_3170_17_lut (.I0(GND_net), .I1(n10675[14]), .I2(GND_net), 
            .I3(n37035), .O(n9933[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_17 (.CI(n37035), .I0(n10675[14]), .I1(GND_net), 
            .CO(n37036));
    SB_LUT4 add_22497_4_lut (.I0(GND_net), .I1(n79[2]), .I2(n191[2]), 
            .I3(n36743), .O(\PID_CONTROLLER.result_31__N_2994 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_11_lut (.I0(GND_net), .I1(n1804[8]), .I2(GND_net), 
            .I3(n38354), .O(n1803[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3102_7_lut (.I0(GND_net), .I1(n8397[4]), .I2(n640_adj_3681), 
            .I3(n38018), .O(n8383[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_7_lut (.I0(GND_net), .I1(n12736[4]), .I2(n472), .I3(n37558), 
            .O(n12161[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_16_lut (.I0(GND_net), .I1(n10675[13]), .I2(GND_net), 
            .I3(n37034), .O(n9933[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_16 (.CI(n37034), .I0(n10675[13]), .I1(GND_net), 
            .CO(n37035));
    SB_LUT4 add_3170_15_lut (.I0(GND_net), .I1(n10675[12]), .I2(GND_net), 
            .I3(n37033), .O(n9933[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_7 (.CI(n38018), .I0(n8397[4]), .I1(n640_adj_3681), 
            .CO(n38019));
    SB_CARRY add_3259_7 (.CI(n37558), .I0(n12736[4]), .I1(n472), .CO(n37559));
    SB_CARRY add_3170_15 (.CI(n37033), .I0(n10675[12]), .I1(GND_net), 
            .CO(n37034));
    SB_LUT4 add_3170_14_lut (.I0(GND_net), .I1(n10675[11]), .I2(GND_net), 
            .I3(n37032), .O(n9933[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3102_6_lut (.I0(GND_net), .I1(n8397[3]), .I2(n543_adj_3682), 
            .I3(n38017), .O(n8383[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_6_lut (.I0(GND_net), .I1(n12736[3]), .I2(n399), .I3(n37557), 
            .O(n12161[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_14 (.CI(n37032), .I0(n10675[11]), .I1(GND_net), 
            .CO(n37033));
    SB_CARRY add_3259_6 (.CI(n37557), .I0(n12736[3]), .I1(n399), .CO(n37558));
    SB_LUT4 add_3170_13_lut (.I0(GND_net), .I1(n10675[10]), .I2(GND_net), 
            .I3(n37031), .O(n9933[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_13 (.CI(n37031), .I0(n10675[10]), .I1(GND_net), 
            .CO(n37032));
    SB_LUT4 add_3170_12_lut (.I0(GND_net), .I1(n10675[9]), .I2(GND_net), 
            .I3(n37030), .O(n9933[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i102_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3170_12 (.CI(n37030), .I0(n10675[9]), .I1(GND_net), .CO(n37031));
    SB_LUT4 add_3170_11_lut (.I0(GND_net), .I1(n10675[8]), .I2(GND_net), 
            .I3(n37029), .O(n9933[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_11 (.CI(n38354), .I0(n1804[8]), .I1(GND_net), 
            .CO(n38355));
    SB_CARRY add_3102_6 (.CI(n38017), .I0(n8397[3]), .I1(n543_adj_3682), 
            .CO(n38018));
    SB_CARRY add_3170_11 (.CI(n37029), .I0(n10675[8]), .I1(GND_net), .CO(n37030));
    SB_LUT4 add_3259_5_lut (.I0(GND_net), .I1(n12736[2]), .I2(n326), .I3(n37556), 
            .O(n12161[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_4 (.CI(n36743), .I0(n79[2]), .I1(n191[2]), .CO(n36744));
    SB_CARRY add_3259_5 (.CI(n37556), .I0(n12736[2]), .I1(n326), .CO(n37557));
    SB_LUT4 add_22497_3_lut (.I0(GND_net), .I1(n79[1]), .I2(n191[1]), 
            .I3(n36742), .O(\PID_CONTROLLER.result_31__N_2994 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_4_lut (.I0(GND_net), .I1(n12736[1]), .I2(n253), .I3(n37555), 
            .O(n12161[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[4]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3102_5_lut (.I0(GND_net), .I1(n8397[2]), .I2(n446_adj_3683), 
            .I3(n38016), .O(n8383[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_10_lut (.I0(GND_net), .I1(n1804[7]), .I2(GND_net), 
            .I3(n38353), .O(n1803[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_5 (.CI(n38016), .I0(n8397[2]), .I1(n446_adj_3683), 
            .CO(n38017));
    SB_CARRY add_3259_4 (.CI(n37555), .I0(n12736[1]), .I1(n253), .CO(n37556));
    SB_LUT4 add_3170_10_lut (.I0(GND_net), .I1(n10675[7]), .I2(GND_net), 
            .I3(n37028), .O(n9933[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_3_lut (.I0(GND_net), .I1(n12736[0]), .I2(n180_adj_3552), 
            .I3(n37554), .O(n12161[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_3 (.CI(n36742), .I0(n79[1]), .I1(n191[1]), .CO(n36743));
    SB_CARRY add_3259_3 (.CI(n37554), .I0(n12736[0]), .I1(n180_adj_3552), 
            .CO(n37555));
    SB_LUT4 add_3259_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n12161[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_10 (.CI(n37028), .I0(n10675[7]), .I1(GND_net), .CO(n37029));
    SB_LUT4 add_3102_4_lut (.I0(GND_net), .I1(n8397[1]), .I2(n349_adj_3685), 
            .I3(n38015), .O(n8383[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n37554));
    SB_LUT4 add_3170_9_lut (.I0(GND_net), .I1(n10675[6]), .I2(GND_net), 
            .I3(n37027), .O(n9933[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_10 (.CI(n38353), .I0(n1804[7]), .I1(GND_net), 
            .CO(n38354));
    SB_CARRY add_3102_4 (.CI(n38015), .I0(n8397[1]), .I1(n349_adj_3685), 
            .CO(n38016));
    SB_CARRY add_3170_9 (.CI(n37027), .I0(n10675[6]), .I1(GND_net), .CO(n37028));
    SB_LUT4 add_3102_3_lut (.I0(GND_net), .I1(n8397[0]), .I2(n252_adj_3686), 
            .I3(n38014), .O(n8383[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_8_lut (.I0(GND_net), .I1(n10675[5]), .I2(n692_adj_3687), 
            .I3(n37026), .O(n9933[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_8 (.CI(n37026), .I0(n10675[5]), .I1(n692_adj_3687), 
            .CO(n37027));
    SB_LUT4 add_3170_7_lut (.I0(GND_net), .I1(n10675[4]), .I2(n595_adj_3688), 
            .I3(n37025), .O(n9933[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_9_lut (.I0(GND_net), .I1(n1804[6]), .I2(GND_net), 
            .I3(n38352), .O(n1803[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_7 (.CI(n37025), .I0(n10675[4]), .I1(n595_adj_3688), 
            .CO(n37026));
    SB_LUT4 add_3170_6_lut (.I0(GND_net), .I1(n10675[3]), .I2(n498_adj_3690), 
            .I3(n37024), .O(n9933[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_6 (.CI(n37024), .I0(n10675[3]), .I1(n498_adj_3690), 
            .CO(n37025));
    SB_CARRY mult_14_add_1218_9 (.CI(n38352), .I0(n1804[6]), .I1(GND_net), 
            .CO(n38353));
    SB_CARRY add_3102_3 (.CI(n38014), .I0(n8397[0]), .I1(n252_adj_3686), 
            .CO(n38015));
    SB_LUT4 mult_14_add_1218_8_lut (.I0(GND_net), .I1(n1804[5]), .I2(n533), 
            .I3(n38351), .O(n1803[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3102_2_lut (.I0(GND_net), .I1(n62_adj_3692), .I2(n155_adj_3693), 
            .I3(GND_net), .O(n8383[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22497_2_lut (.I0(GND_net), .I1(n79[0]), .I2(n191[0]), 
            .I3(GND_net), .O(\PID_CONTROLLER.result_31__N_2994 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22497_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22497_2 (.CI(GND_net), .I0(n79[0]), .I1(n191[0]), .CO(n36742));
    SB_CARRY add_3102_2 (.CI(GND_net), .I0(n62_adj_3692), .I1(n155_adj_3693), 
            .CO(n38014));
    SB_LUT4 add_3170_5_lut (.I0(GND_net), .I1(n10675[2]), .I2(n401_adj_3694), 
            .I3(n37023), .O(n9933[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_14_lut (.I0(GND_net), .I1(n8383[11]), .I2(GND_net), 
            .I3(n38013), .O(n8368[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_5 (.CI(n37023), .I0(n10675[2]), .I1(n401_adj_3694), 
            .CO(n37024));
    SB_CARRY mult_14_add_1218_8 (.CI(n38351), .I0(n1804[5]), .I1(n533), 
            .CO(n38352));
    SB_LUT4 add_3101_13_lut (.I0(GND_net), .I1(n8383[10]), .I2(GND_net), 
            .I3(n38012), .O(n8368[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_4_lut (.I0(GND_net), .I1(n10675[1]), .I2(n304_adj_3695), 
            .I3(n37022), .O(n9933[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_4 (.CI(n37022), .I0(n10675[1]), .I1(n304_adj_3695), 
            .CO(n37023));
    SB_LUT4 add_3170_3_lut (.I0(GND_net), .I1(n10675[0]), .I2(n207_adj_3696), 
            .I3(n37021), .O(n9933[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_3 (.CI(n37021), .I0(n10675[0]), .I1(n207_adj_3696), 
            .CO(n37022));
    SB_CARRY add_3101_13 (.CI(n38012), .I0(n8383[10]), .I1(GND_net), .CO(n38013));
    SB_LUT4 add_3170_2_lut (.I0(GND_net), .I1(n17_adj_3697), .I2(n110_adj_3698), 
            .I3(GND_net), .O(n9933[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_19_lut (.I0(GND_net), .I1(n15118[16]), .I2(GND_net), 
            .I3(n36741), .O(n14797[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_2 (.CI(GND_net), .I0(n17_adj_3697), .I1(n110_adj_3698), 
            .CO(n37021));
    SB_LUT4 add_3382_18_lut (.I0(GND_net), .I1(n15118[15]), .I2(GND_net), 
            .I3(n36740), .O(n14797[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3350_13_lut (.I0(GND_net), .I1(n14564[10]), .I2(GND_net), 
            .I3(n37020), .O(n14172[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_18 (.CI(n36740), .I0(n15118[15]), .I1(GND_net), 
            .CO(n36741));
    SB_LUT4 add_3382_17_lut (.I0(GND_net), .I1(n15118[14]), .I2(GND_net), 
            .I3(n36739), .O(n14797[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3350_12_lut (.I0(GND_net), .I1(n14564[9]), .I2(GND_net), 
            .I3(n37019), .O(n14172[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_12 (.CI(n37019), .I0(n14564[9]), .I1(GND_net), .CO(n37020));
    SB_LUT4 add_3350_11_lut (.I0(GND_net), .I1(n14564[8]), .I2(GND_net), 
            .I3(n37018), .O(n14172[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_7_lut (.I0(GND_net), .I1(n1804[4]), .I2(n460_c), 
            .I3(n38350), .O(n1803[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_11 (.CI(n37018), .I0(n14564[8]), .I1(GND_net), .CO(n37019));
    SB_LUT4 add_3101_12_lut (.I0(GND_net), .I1(n8383[9]), .I2(GND_net), 
            .I3(n38011), .O(n8368[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_12 (.CI(n38011), .I0(n8383[9]), .I1(GND_net), .CO(n38012));
    SB_LUT4 add_3350_10_lut (.I0(GND_net), .I1(n14564[7]), .I2(GND_net), 
            .I3(n37017), .O(n14172[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_11_lut (.I0(GND_net), .I1(n8383[8]), .I2(GND_net), 
            .I3(n38010), .O(n8368[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_10 (.CI(n37017), .I0(n14564[7]), .I1(GND_net), .CO(n37018));
    SB_LUT4 add_3350_9_lut (.I0(GND_net), .I1(n14564[6]), .I2(GND_net), 
            .I3(n37016), .O(n14172[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_9 (.CI(n37016), .I0(n14564[6]), .I1(GND_net), .CO(n37017));
    SB_CARRY mult_14_add_1218_7 (.CI(n38350), .I0(n1804[4]), .I1(n460_c), 
            .CO(n38351));
    SB_CARRY add_3101_11 (.CI(n38010), .I0(n8383[8]), .I1(GND_net), .CO(n38011));
    SB_LUT4 add_3350_8_lut (.I0(GND_net), .I1(n14564[5]), .I2(n545), .I3(n37015), 
            .O(n14172[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_8 (.CI(n37015), .I0(n14564[5]), .I1(n545), .CO(n37016));
    SB_LUT4 add_3350_7_lut (.I0(GND_net), .I1(n14564[4]), .I2(n472), .I3(n37014), 
            .O(n14172[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_10_lut (.I0(GND_net), .I1(n8383[7]), .I2(GND_net), 
            .I3(n38009), .O(n8368[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_7 (.CI(n37014), .I0(n14564[4]), .I1(n472), .CO(n37015));
    SB_LUT4 add_3350_6_lut (.I0(GND_net), .I1(n14564[3]), .I2(n399), .I3(n37013), 
            .O(n14172[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_6 (.CI(n37013), .I0(n14564[3]), .I1(n399), .CO(n37014));
    SB_CARRY add_3382_17 (.CI(n36739), .I0(n15118[14]), .I1(GND_net), 
            .CO(n36740));
    SB_CARRY add_3101_10 (.CI(n38009), .I0(n8383[7]), .I1(GND_net), .CO(n38010));
    SB_LUT4 mult_14_add_1218_6_lut (.I0(GND_net), .I1(n1804[3]), .I2(n387_c), 
            .I3(n38349), .O(n1803[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_9_lut (.I0(GND_net), .I1(n8383[6]), .I2(GND_net), 
            .I3(n38008), .O(n8368[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3350_5_lut (.I0(GND_net), .I1(n14564[2]), .I2(n326), .I3(n37012), 
            .O(n14172[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_9 (.CI(n38008), .I0(n8383[6]), .I1(GND_net), .CO(n38009));
    SB_CARRY add_3350_5 (.CI(n37012), .I0(n14564[2]), .I1(n326), .CO(n37013));
    SB_LUT4 add_3350_4_lut (.I0(GND_net), .I1(n14564[1]), .I2(n253), .I3(n37011), 
            .O(n14172[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_4 (.CI(n37011), .I0(n14564[1]), .I1(n253), .CO(n37012));
    SB_LUT4 add_3101_8_lut (.I0(GND_net), .I1(n8383[5]), .I2(n734_adj_3700), 
            .I3(n38007), .O(n8368[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3350_3_lut (.I0(GND_net), .I1(n14564[0]), .I2(n180_adj_3552), 
            .I3(n37010), .O(n14172[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_3 (.CI(n37010), .I0(n14564[0]), .I1(n180_adj_3552), 
            .CO(n37011));
    SB_LUT4 add_3350_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n14172[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_6 (.CI(n38349), .I0(n1804[3]), .I1(n387_c), 
            .CO(n38350));
    SB_LUT4 mult_12_i91_2_lut (.I0(\Kd[1] ), .I1(n67[12]), .I2(GND_net), 
            .I3(GND_net), .O(n134));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i91_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3101_8 (.CI(n38007), .I0(n8383[5]), .I1(n734_adj_3700), 
            .CO(n38008));
    SB_CARRY add_3350_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n37010));
    SB_LUT4 add_3382_16_lut (.I0(GND_net), .I1(n15118[13]), .I2(GND_net), 
            .I3(n36738), .O(n14797[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_16 (.CI(n36738), .I0(n15118[13]), .I1(GND_net), 
            .CO(n36739));
    SB_LUT4 add_3198_27_lut (.I0(GND_net), .I1(n11362[24]), .I2(GND_net), 
            .I3(n37009), .O(n10675[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_7_lut (.I0(GND_net), .I1(n8383[4]), .I2(n637_adj_3701), 
            .I3(n38006), .O(n8368[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_5_lut (.I0(GND_net), .I1(n1804[2]), .I2(n314_adj_3703), 
            .I3(n38348), .O(n1803[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_5 (.CI(n38348), .I0(n1804[2]), .I1(n314_adj_3703), 
            .CO(n38349));
    SB_LUT4 mult_14_add_1218_4_lut (.I0(GND_net), .I1(n1804[1]), .I2(n241_adj_3705), 
            .I3(n38347), .O(n1803[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_4 (.CI(n38347), .I0(n1804[1]), .I1(n241_adj_3705), 
            .CO(n38348));
    SB_LUT4 add_3198_26_lut (.I0(GND_net), .I1(n11362[23]), .I2(GND_net), 
            .I3(n37008), .O(n10675[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_3_lut (.I0(GND_net), .I1(n1804[0]), .I2(n168_adj_3707), 
            .I3(n38346), .O(n1803[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_15_lut (.I0(GND_net), .I1(n15118[12]), .I2(GND_net), 
            .I3(n36737), .O(n14797[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_7 (.CI(n38006), .I0(n8383[4]), .I1(n637_adj_3701), 
            .CO(n38007));
    SB_LUT4 add_3101_6_lut (.I0(GND_net), .I1(n8383[3]), .I2(n540_adj_3708), 
            .I3(n38005), .O(n8368[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_3 (.CI(n38346), .I0(n1804[0]), .I1(n168_adj_3707), 
            .CO(n38347));
    SB_CARRY add_3101_6 (.CI(n38005), .I0(n8383[3]), .I1(n540_adj_3708), 
            .CO(n38006));
    SB_LUT4 add_3101_5_lut (.I0(GND_net), .I1(n8383[2]), .I2(n443_adj_3709), 
            .I3(n38004), .O(n8368[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_15 (.CI(n36737), .I0(n15118[12]), .I1(GND_net), 
            .CO(n36738));
    SB_LUT4 add_3382_14_lut (.I0(GND_net), .I1(n15118[11]), .I2(GND_net), 
            .I3(n36736), .O(n14797[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_2_lut (.I0(GND_net), .I1(n26_adj_3710), .I2(n95), 
            .I3(GND_net), .O(n1803[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_5 (.CI(n38004), .I0(n8383[2]), .I1(n443_adj_3709), 
            .CO(n38005));
    SB_CARRY mult_14_add_1218_2 (.CI(GND_net), .I0(n26_adj_3710), .I1(n95), 
            .CO(n38346));
    SB_LUT4 add_3101_4_lut (.I0(GND_net), .I1(n8383[1]), .I2(n346_adj_3711), 
            .I3(n38003), .O(n8368[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_26 (.CI(n37008), .I0(n11362[23]), .I1(GND_net), 
            .CO(n37009));
    SB_LUT4 add_3198_25_lut (.I0(GND_net), .I1(n11362[22]), .I2(GND_net), 
            .I3(n37007), .O(n10675[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_4 (.CI(n38003), .I0(n8383[1]), .I1(n346_adj_3711), 
            .CO(n38004));
    SB_CARRY add_3198_25 (.CI(n37007), .I0(n11362[22]), .I1(GND_net), 
            .CO(n37008));
    SB_LUT4 add_3198_24_lut (.I0(GND_net), .I1(n11362[21]), .I2(GND_net), 
            .I3(n37006), .O(n10675[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_14 (.CI(n36736), .I0(n15118[11]), .I1(GND_net), 
            .CO(n36737));
    SB_CARRY add_3198_24 (.CI(n37006), .I0(n11362[21]), .I1(GND_net), 
            .CO(n37007));
    SB_LUT4 mult_14_add_1217_24_lut (.I0(GND_net), .I1(n1803[21]), .I2(GND_net), 
            .I3(n38344), .O(n1802[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_3_lut (.I0(GND_net), .I1(n8383[0]), .I2(n249_adj_3712), 
            .I3(n38002), .O(n8368[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_23_lut (.I0(GND_net), .I1(n11362[20]), .I2(GND_net), 
            .I3(n37005), .O(n10675[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_13_lut (.I0(GND_net), .I1(n15118[10]), .I2(GND_net), 
            .I3(n36735), .O(n14797[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_13 (.CI(n36735), .I0(n15118[10]), .I1(GND_net), 
            .CO(n36736));
    SB_CARRY add_3198_23 (.CI(n37005), .I0(n11362[20]), .I1(GND_net), 
            .CO(n37006));
    SB_LUT4 add_3198_22_lut (.I0(GND_net), .I1(n11362[19]), .I2(GND_net), 
            .I3(n37004), .O(n10675[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_22 (.CI(n37004), .I0(n11362[19]), .I1(GND_net), 
            .CO(n37005));
    SB_LUT4 add_3198_21_lut (.I0(GND_net), .I1(n11362[18]), .I2(GND_net), 
            .I3(n37003), .O(n10675[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_3 (.CI(n38002), .I0(n8383[0]), .I1(n249_adj_3712), 
            .CO(n38003));
    SB_CARRY add_3198_21 (.CI(n37003), .I0(n11362[18]), .I1(GND_net), 
            .CO(n37004));
    SB_LUT4 add_3382_12_lut (.I0(GND_net), .I1(n15118[9]), .I2(GND_net), 
            .I3(n36734), .O(n14797[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_12 (.CI(n36734), .I0(n15118[9]), .I1(GND_net), .CO(n36735));
    SB_LUT4 add_3198_20_lut (.I0(GND_net), .I1(n11362[17]), .I2(GND_net), 
            .I3(n37002), .O(n10675[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_20 (.CI(n37002), .I0(n11362[17]), .I1(GND_net), 
            .CO(n37003));
    SB_LUT4 add_3101_2_lut (.I0(GND_net), .I1(n59_adj_3713), .I2(n152_adj_3714), 
            .I3(GND_net), .O(n8368[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_19_lut (.I0(GND_net), .I1(n11362[16]), .I2(GND_net), 
            .I3(n37001), .O(n10675[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_19 (.CI(n37001), .I0(n11362[16]), .I1(GND_net), 
            .CO(n37002));
    SB_LUT4 add_3382_11_lut (.I0(GND_net), .I1(n15118[8]), .I2(GND_net), 
            .I3(n36733), .O(n14797[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_11 (.CI(n36733), .I0(n15118[8]), .I1(GND_net), .CO(n36734));
    SB_LUT4 add_3198_18_lut (.I0(GND_net), .I1(n11362[15]), .I2(GND_net), 
            .I3(n37000), .O(n10675[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_18 (.CI(n37000), .I0(n11362[15]), .I1(GND_net), 
            .CO(n37001));
    SB_CARRY mult_14_add_1217_24 (.CI(n38344), .I0(n1803[21]), .I1(GND_net), 
            .CO(n1707));
    SB_CARRY add_3101_2 (.CI(GND_net), .I0(n59_adj_3713), .I1(n152_adj_3714), 
            .CO(n38002));
    SB_LUT4 add_3382_10_lut (.I0(GND_net), .I1(n15118[7]), .I2(GND_net), 
            .I3(n36732), .O(n14797[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_17_lut (.I0(GND_net), .I1(n11362[14]), .I2(GND_net), 
            .I3(n36999), .O(n10675[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_17 (.CI(n36999), .I0(n11362[14]), .I1(GND_net), 
            .CO(n37000));
    SB_LUT4 mult_14_add_1217_23_lut (.I0(GND_net), .I1(n1803[20]), .I2(GND_net), 
            .I3(n38343), .O(n1802[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_16_lut (.I0(GND_net), .I1(n11362[13]), .I2(GND_net), 
            .I3(n36998), .O(n10675[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_16 (.CI(n36998), .I0(n11362[13]), .I1(GND_net), 
            .CO(n36999));
    SB_CARRY add_3382_10 (.CI(n36732), .I0(n15118[7]), .I1(GND_net), .CO(n36733));
    SB_LUT4 add_3382_9_lut (.I0(GND_net), .I1(n15118[6]), .I2(GND_net), 
            .I3(n36731), .O(n14797[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_15_lut (.I0(GND_net), .I1(n11362[12]), .I2(GND_net), 
            .I3(n36997), .O(n10675[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_15 (.CI(n36997), .I0(n11362[12]), .I1(GND_net), 
            .CO(n36998));
    SB_LUT4 add_3100_15_lut (.I0(GND_net), .I1(n8368[12]), .I2(GND_net), 
            .I3(n38001), .O(n8352[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_14_lut (.I0(GND_net), .I1(n8368[11]), .I2(GND_net), 
            .I3(n38000), .O(n8352[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_14_lut (.I0(GND_net), .I1(n11362[11]), .I2(GND_net), 
            .I3(n36996), .O(n10675[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_9 (.CI(n36731), .I0(n15118[6]), .I1(GND_net), .CO(n36732));
    SB_CARRY add_3198_14 (.CI(n36996), .I0(n11362[11]), .I1(GND_net), 
            .CO(n36997));
    SB_LUT4 add_3198_13_lut (.I0(GND_net), .I1(n11362[10]), .I2(GND_net), 
            .I3(n36995), .O(n10675[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_8_lut (.I0(GND_net), .I1(n15118[5]), .I2(n719), .I3(n36730), 
            .O(n14797[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_8 (.CI(n36730), .I0(n15118[5]), .I1(n719), .CO(n36731));
    SB_CARRY add_3198_13 (.CI(n36995), .I0(n11362[10]), .I1(GND_net), 
            .CO(n36996));
    SB_LUT4 add_3198_12_lut (.I0(GND_net), .I1(n11362[9]), .I2(GND_net), 
            .I3(n36994), .O(n10675[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_12 (.CI(n36994), .I0(n11362[9]), .I1(GND_net), .CO(n36995));
    SB_LUT4 add_3382_7_lut (.I0(GND_net), .I1(n15118[4]), .I2(n622), .I3(n36729), 
            .O(n14797[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_11_lut (.I0(GND_net), .I1(n11362[8]), .I2(GND_net), 
            .I3(n36993), .O(n10675[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_7 (.CI(n36729), .I0(n15118[4]), .I1(n622), .CO(n36730));
    SB_CARRY mult_14_add_1217_23 (.CI(n38343), .I0(n1803[20]), .I1(GND_net), 
            .CO(n38344));
    SB_LUT4 mult_14_add_1217_22_lut (.I0(GND_net), .I1(n1803[19]), .I2(GND_net), 
            .I3(n38342), .O(n1802[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_22 (.CI(n38342), .I0(n1803[19]), .I1(GND_net), 
            .CO(n38343));
    SB_CARRY add_3100_14 (.CI(n38000), .I0(n8368[11]), .I1(GND_net), .CO(n38001));
    SB_CARRY add_3198_11 (.CI(n36993), .I0(n11362[8]), .I1(GND_net), .CO(n36994));
    SB_LUT4 add_3198_10_lut (.I0(GND_net), .I1(n11362[7]), .I2(GND_net), 
            .I3(n36992), .O(n10675[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_6_lut (.I0(GND_net), .I1(n15118[3]), .I2(n525_adj_3715), 
            .I3(n36728), .O(n14797[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_6 (.CI(n36728), .I0(n15118[3]), .I1(n525_adj_3715), 
            .CO(n36729));
    SB_CARRY add_3198_10 (.CI(n36992), .I0(n11362[7]), .I1(GND_net), .CO(n36993));
    SB_LUT4 add_3198_9_lut (.I0(GND_net), .I1(n11362[6]), .I2(GND_net), 
            .I3(n36991), .O(n10675[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_13_lut (.I0(GND_net), .I1(n8368[10]), .I2(GND_net), 
            .I3(n37999), .O(n8352[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_9 (.CI(n36991), .I0(n11362[6]), .I1(GND_net), .CO(n36992));
    SB_CARRY add_3100_13 (.CI(n37999), .I0(n8368[10]), .I1(GND_net), .CO(n38000));
    SB_LUT4 add_3198_8_lut (.I0(GND_net), .I1(n11362[5]), .I2(n695_adj_3716), 
            .I3(n36990), .O(n10675[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_8 (.CI(n36990), .I0(n11362[5]), .I1(n695_adj_3716), 
            .CO(n36991));
    SB_LUT4 add_3198_7_lut (.I0(GND_net), .I1(n11362[4]), .I2(n598_adj_3717), 
            .I3(n36989), .O(n10675[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_12_lut (.I0(GND_net), .I1(n8368[9]), .I2(GND_net), 
            .I3(n37998), .O(n8352[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_7 (.CI(n36989), .I0(n11362[4]), .I1(n598_adj_3717), 
            .CO(n36990));
    SB_LUT4 add_3382_5_lut (.I0(GND_net), .I1(n15118[2]), .I2(n428), .I3(n36727), 
            .O(n14797[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_6_lut (.I0(GND_net), .I1(n11362[3]), .I2(n501_adj_3718), 
            .I3(n36988), .O(n10675[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_5 (.CI(n36727), .I0(n15118[2]), .I1(n428), .CO(n36728));
    SB_LUT4 mult_14_add_1217_21_lut (.I0(GND_net), .I1(n1803[18]), .I2(GND_net), 
            .I3(n38341), .O(n1802[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_12 (.CI(n37998), .I0(n8368[9]), .I1(GND_net), .CO(n37999));
    SB_CARRY add_3198_6 (.CI(n36988), .I0(n11362[3]), .I1(n501_adj_3718), 
            .CO(n36989));
    SB_LUT4 add_3198_5_lut (.I0(GND_net), .I1(n11362[2]), .I2(n404_adj_3719), 
            .I3(n36987), .O(n10675[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_5 (.CI(n36987), .I0(n11362[2]), .I1(n404_adj_3719), 
            .CO(n36988));
    SB_LUT4 add_3100_11_lut (.I0(GND_net), .I1(n8368[8]), .I2(GND_net), 
            .I3(n37997), .O(n8352[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_4_lut (.I0(GND_net), .I1(n11362[1]), .I2(n307_adj_3720), 
            .I3(n36986), .O(n10675[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_4_lut (.I0(GND_net), .I1(n15118[1]), .I2(n331), .I3(n36726), 
            .O(n14797[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_4 (.CI(n36986), .I0(n11362[1]), .I1(n307_adj_3720), 
            .CO(n36987));
    SB_CARRY add_3382_4 (.CI(n36726), .I0(n15118[1]), .I1(n331), .CO(n36727));
    SB_CARRY mult_14_add_1217_21 (.CI(n38341), .I0(n1803[18]), .I1(GND_net), 
            .CO(n38342));
    SB_CARRY add_3100_11 (.CI(n37997), .I0(n8368[8]), .I1(GND_net), .CO(n37998));
    SB_LUT4 add_3198_3_lut (.I0(GND_net), .I1(n11362[0]), .I2(n210_adj_3721), 
            .I3(n36985), .O(n10675[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_3 (.CI(n36985), .I0(n11362[0]), .I1(n210_adj_3721), 
            .CO(n36986));
    SB_LUT4 add_3100_10_lut (.I0(GND_net), .I1(n8368[7]), .I2(GND_net), 
            .I3(n37996), .O(n8352[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_2_lut (.I0(GND_net), .I1(n20_adj_3722), .I2(n113_adj_3723), 
            .I3(GND_net), .O(n10675[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_3_lut (.I0(GND_net), .I1(n15118[0]), .I2(n234_adj_3724), 
            .I3(n36725), .O(n14797[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_2 (.CI(GND_net), .I0(n20_adj_3722), .I1(n113_adj_3723), 
            .CO(n36985));
    SB_CARRY add_3382_3 (.CI(n36725), .I0(n15118[0]), .I1(n234_adj_3724), 
            .CO(n36726));
    SB_LUT4 mult_14_add_1217_20_lut (.I0(GND_net), .I1(n1803[17]), .I2(GND_net), 
            .I3(n38340), .O(n1802[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_10 (.CI(n37996), .I0(n8368[7]), .I1(GND_net), .CO(n37997));
    SB_LUT4 add_3370_12_lut (.I0(GND_net), .I1(n14916[9]), .I2(GND_net), 
            .I3(n36984), .O(n14564[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_11_lut (.I0(GND_net), .I1(n14916[8]), .I2(GND_net), 
            .I3(n36983), .O(n14564[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_20 (.CI(n38340), .I0(n1803[17]), .I1(GND_net), 
            .CO(n38341));
    SB_LUT4 add_3100_9_lut (.I0(GND_net), .I1(n8368[6]), .I2(GND_net), 
            .I3(n37995), .O(n8352[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_11 (.CI(n36983), .I0(n14916[8]), .I1(GND_net), .CO(n36984));
    SB_CARRY add_3100_9 (.CI(n37995), .I0(n8368[6]), .I1(GND_net), .CO(n37996));
    SB_LUT4 add_3370_10_lut (.I0(GND_net), .I1(n14916[7]), .I2(GND_net), 
            .I3(n36982), .O(n14564[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_2_lut (.I0(GND_net), .I1(n44), .I2(n137_adj_3725), 
            .I3(GND_net), .O(n14797[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_8_lut (.I0(GND_net), .I1(n8368[5]), .I2(n731_adj_3726), 
            .I3(n37994), .O(n8352[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_10 (.CI(n36982), .I0(n14916[7]), .I1(GND_net), .CO(n36983));
    SB_CARRY add_3382_2 (.CI(GND_net), .I0(n44), .I1(n137_adj_3725), .CO(n36725));
    SB_LUT4 add_3370_9_lut (.I0(GND_net), .I1(n14916[6]), .I2(GND_net), 
            .I3(n36981), .O(n14564[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_9 (.CI(n36981), .I0(n14916[6]), .I1(GND_net), .CO(n36982));
    SB_LUT4 mult_14_add_1217_19_lut (.I0(GND_net), .I1(n1803[16]), .I2(GND_net), 
            .I3(n38339), .O(n1802[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_8_lut (.I0(GND_net), .I1(n14916[5]), .I2(n545), .I3(n36980), 
            .O(n14564[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_8 (.CI(n37994), .I0(n8368[5]), .I1(n731_adj_3726), 
            .CO(n37995));
    SB_CARRY add_3370_8 (.CI(n36980), .I0(n14916[5]), .I1(n545), .CO(n36981));
    SB_LUT4 add_3370_7_lut (.I0(GND_net), .I1(n14916[4]), .I2(n472), .I3(n36979), 
            .O(n14564[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_7 (.CI(n36979), .I0(n14916[4]), .I1(n472), .CO(n36980));
    SB_LUT4 add_3100_7_lut (.I0(GND_net), .I1(n8368[4]), .I2(n634_adj_3727), 
            .I3(n37993), .O(n8352[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_19 (.CI(n38339), .I0(n1803[16]), .I1(GND_net), 
            .CO(n38340));
    SB_LUT4 add_3370_6_lut (.I0(GND_net), .I1(n14916[3]), .I2(n399), .I3(n36978), 
            .O(n14564[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_6 (.CI(n36978), .I0(n14916[3]), .I1(n399), .CO(n36979));
    SB_LUT4 add_3370_5_lut (.I0(GND_net), .I1(n14916[2]), .I2(n326), .I3(n36977), 
            .O(n14564[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_33_lut (.I0(GND_net), .I1(n7069[8]), 
            .I2(n5790[0]), .I3(n36724), .O(n79[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_5 (.CI(n36977), .I0(n14916[2]), .I1(n326), .CO(n36978));
    SB_LUT4 add_3370_4_lut (.I0(GND_net), .I1(n14916[1]), .I2(n253), .I3(n36976), 
            .O(n14564[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_4 (.CI(n36976), .I0(n14916[1]), .I1(n253), .CO(n36977));
    SB_LUT4 add_13_add_1_22497_add_1_32_lut (.I0(GND_net), .I1(n7069[7]), 
            .I2(n76[30]), .I3(n36723), .O(n79[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_32 (.CI(n36723), .I0(n7069[7]), .I1(n76[30]), 
            .CO(n36724));
    SB_CARRY add_3100_7 (.CI(n37993), .I0(n8368[4]), .I1(n634_adj_3727), 
            .CO(n37994));
    SB_LUT4 add_3370_3_lut (.I0(GND_net), .I1(n14916[0]), .I2(n180_adj_3552), 
            .I3(n36975), .O(n14564[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_31_lut (.I0(GND_net), .I1(n7069[6]), 
            .I2(n76[29]), .I3(n36722), .O(n79[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_31 (.CI(n36722), .I0(n7069[6]), .I1(n76[29]), 
            .CO(n36723));
    SB_LUT4 add_13_add_1_22497_add_1_30_lut (.I0(GND_net), .I1(n7069[5]), 
            .I2(n76[28]), .I3(n36721), .O(n79[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_3 (.CI(n36975), .I0(n14916[0]), .I1(n180_adj_3552), 
            .CO(n36976));
    SB_LUT4 add_3370_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n14564[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n36975));
    SB_LUT4 add_3100_6_lut (.I0(GND_net), .I1(n8368[3]), .I2(n537_adj_3728), 
            .I3(n37992), .O(n8352[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_26_lut (.I0(GND_net), .I1(n11996[23]), .I2(GND_net), 
            .I3(n36974), .O(n11362[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_25_lut (.I0(GND_net), .I1(n11996[22]), .I2(GND_net), 
            .I3(n36973), .O(n11362[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_18_lut (.I0(GND_net), .I1(n1803[15]), .I2(GND_net), 
            .I3(n38338), .O(n1802[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_18 (.CI(n38338), .I0(n1803[15]), .I1(GND_net), 
            .CO(n38339));
    SB_CARRY add_3225_25 (.CI(n36973), .I0(n11996[22]), .I1(GND_net), 
            .CO(n36974));
    SB_CARRY add_13_add_1_22497_add_1_30 (.CI(n36721), .I0(n7069[5]), .I1(n76[28]), 
            .CO(n36722));
    SB_LUT4 mult_14_add_1217_17_lut (.I0(GND_net), .I1(n1803[14]), .I2(GND_net), 
            .I3(n38337), .O(n1802[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_6 (.CI(n37992), .I0(n8368[3]), .I1(n537_adj_3728), 
            .CO(n37993));
    SB_CARRY mult_14_add_1217_17 (.CI(n38337), .I0(n1803[14]), .I1(GND_net), 
            .CO(n38338));
    SB_LUT4 add_13_add_1_22497_add_1_29_lut (.I0(GND_net), .I1(n7069[4]), 
            .I2(n76[27]), .I3(n36720), .O(n79[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_16_lut (.I0(GND_net), .I1(n1803[13]), .I2(GND_net), 
            .I3(n38336), .O(n1802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_5_lut (.I0(GND_net), .I1(n8368[2]), .I2(n440_adj_3729), 
            .I3(n37991), .O(n8352[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_5 (.CI(n37991), .I0(n8368[2]), .I1(n440_adj_3729), 
            .CO(n37992));
    SB_LUT4 add_3225_24_lut (.I0(GND_net), .I1(n11996[21]), .I2(GND_net), 
            .I3(n36972), .O(n11362[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_4_lut (.I0(GND_net), .I1(n8368[1]), .I2(n343_adj_3730), 
            .I3(n37990), .O(n8352[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_16 (.CI(n38336), .I0(n1803[13]), .I1(GND_net), 
            .CO(n38337));
    SB_CARRY add_3225_24 (.CI(n36972), .I0(n11996[21]), .I1(GND_net), 
            .CO(n36973));
    SB_LUT4 add_3225_23_lut (.I0(GND_net), .I1(n11996[20]), .I2(GND_net), 
            .I3(n36971), .O(n11362[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_4 (.CI(n37990), .I0(n8368[1]), .I1(n343_adj_3730), 
            .CO(n37991));
    SB_LUT4 add_3100_3_lut (.I0(GND_net), .I1(n8368[0]), .I2(n246_adj_3731), 
            .I3(n37989), .O(n8352[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_23 (.CI(n36971), .I0(n11996[20]), .I1(GND_net), 
            .CO(n36972));
    SB_LUT4 add_3225_22_lut (.I0(GND_net), .I1(n11996[19]), .I2(GND_net), 
            .I3(n36970), .O(n11362[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_15_lut (.I0(GND_net), .I1(n1803[12]), .I2(GND_net), 
            .I3(n38335), .O(n1802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_22 (.CI(n36970), .I0(n11996[19]), .I1(GND_net), 
            .CO(n36971));
    SB_CARRY add_3100_3 (.CI(n37989), .I0(n8368[0]), .I1(n246_adj_3731), 
            .CO(n37990));
    SB_LUT4 add_3225_21_lut (.I0(GND_net), .I1(n11996[18]), .I2(GND_net), 
            .I3(n36969), .O(n11362[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_21 (.CI(n36969), .I0(n11996[18]), .I1(GND_net), 
            .CO(n36970));
    SB_CARRY add_13_add_1_22497_add_1_29 (.CI(n36720), .I0(n7069[4]), .I1(n76[27]), 
            .CO(n36721));
    SB_LUT4 add_3225_20_lut (.I0(GND_net), .I1(n11996[17]), .I2(GND_net), 
            .I3(n36968), .O(n11362[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_20 (.CI(n36968), .I0(n11996[17]), .I1(GND_net), 
            .CO(n36969));
    SB_LUT4 add_3225_19_lut (.I0(GND_net), .I1(n11996[16]), .I2(GND_net), 
            .I3(n36967), .O(n11362[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_19 (.CI(n36967), .I0(n11996[16]), .I1(GND_net), 
            .CO(n36968));
    SB_LUT4 add_3100_2_lut (.I0(GND_net), .I1(n56_adj_3732), .I2(n149_adj_3733), 
            .I3(GND_net), .O(n8352[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_18_lut (.I0(GND_net), .I1(n11996[15]), .I2(GND_net), 
            .I3(n36966), .O(n11362[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_28_lut (.I0(GND_net), .I1(n7069[3]), 
            .I2(n76[26]), .I3(n36719), .O(n79[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_18 (.CI(n36966), .I0(n11996[15]), .I1(GND_net), 
            .CO(n36967));
    SB_CARRY add_13_add_1_22497_add_1_28 (.CI(n36719), .I0(n7069[3]), .I1(n76[26]), 
            .CO(n36720));
    SB_CARRY mult_14_add_1217_15 (.CI(n38335), .I0(n1803[12]), .I1(GND_net), 
            .CO(n38336));
    SB_CARRY add_3100_2 (.CI(GND_net), .I0(n56_adj_3732), .I1(n149_adj_3733), 
            .CO(n37989));
    SB_LUT4 add_13_add_1_22497_add_1_27_lut (.I0(GND_net), .I1(n7069[2]), 
            .I2(n76[25]), .I3(n36718), .O(n79[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_17_lut (.I0(GND_net), .I1(n11996[14]), .I2(GND_net), 
            .I3(n36965), .O(n11362[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_17 (.CI(n36965), .I0(n11996[14]), .I1(GND_net), 
            .CO(n36966));
    SB_LUT4 add_3099_16_lut (.I0(GND_net), .I1(n8352[13]), .I2(GND_net), 
            .I3(n37988), .O(n8335[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_27 (.CI(n36718), .I0(n7069[2]), .I1(n76[25]), 
            .CO(n36719));
    SB_LUT4 add_3225_16_lut (.I0(GND_net), .I1(n11996[13]), .I2(GND_net), 
            .I3(n36964), .O(n11362[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_26_lut (.I0(GND_net), .I1(n7069[1]), 
            .I2(n76[24]), .I3(n36717), .O(n79[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_16 (.CI(n36964), .I0(n11996[13]), .I1(GND_net), 
            .CO(n36965));
    SB_CARRY add_13_add_1_22497_add_1_26 (.CI(n36717), .I0(n7069[1]), .I1(n76[24]), 
            .CO(n36718));
    SB_LUT4 mult_14_add_1217_14_lut (.I0(GND_net), .I1(n1803[11]), .I2(GND_net), 
            .I3(n38334), .O(n1802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_25_lut (.I0(GND_net), .I1(n7069[0]), 
            .I2(n76[23]), .I3(n36716), .O(n79[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_15_lut (.I0(GND_net), .I1(n8352[12]), .I2(GND_net), 
            .I3(n37987), .O(n8335[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_15 (.CI(n37987), .I0(n8352[12]), .I1(GND_net), .CO(n37988));
    SB_CARRY mult_14_add_1217_14 (.CI(n38334), .I0(n1803[11]), .I1(GND_net), 
            .CO(n38335));
    SB_LUT4 add_3099_14_lut (.I0(GND_net), .I1(n8352[11]), .I2(GND_net), 
            .I3(n37986), .O(n8335[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_15_lut (.I0(GND_net), .I1(n11996[12]), .I2(GND_net), 
            .I3(n36963), .O(n11362[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_15 (.CI(n36963), .I0(n11996[12]), .I1(GND_net), 
            .CO(n36964));
    SB_CARRY add_3099_14 (.CI(n37986), .I0(n8352[11]), .I1(GND_net), .CO(n37987));
    SB_LUT4 add_3099_13_lut (.I0(GND_net), .I1(n8352[10]), .I2(GND_net), 
            .I3(n37985), .O(n8335[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n37507), .O(n82[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_14_lut (.I0(GND_net), .I1(n11996[11]), .I2(GND_net), 
            .I3(n36962), .O(n11362[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_25 (.CI(n36716), .I0(n7069[0]), .I1(n76[23]), 
            .CO(n36717));
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n37506), .O(n82[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_14 (.CI(n36962), .I0(n11996[11]), .I1(GND_net), 
            .CO(n36963));
    SB_LUT4 add_13_add_1_22497_add_1_24_lut (.I0(GND_net), .I1(n282[22]), 
            .I2(n76[22]), .I3(n36715), .O(n79[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_13_lut (.I0(GND_net), .I1(n11996[10]), .I2(GND_net), 
            .I3(n36961), .O(n11362[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_13_lut (.I0(GND_net), .I1(n1803[10]), .I2(GND_net), 
            .I3(n38333), .O(n1802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_13 (.CI(n38333), .I0(n1803[10]), .I1(GND_net), 
            .CO(n38334));
    SB_CARRY add_3099_13 (.CI(n37985), .I0(n8352[10]), .I1(GND_net), .CO(n37986));
    SB_CARRY \PID_CONTROLLER.integral_1049_add_4_10  (.CI(n37506), .I0(\PID_CONTROLLER.err[8] ), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n37507));
    SB_LUT4 mult_14_add_1217_12_lut (.I0(GND_net), .I1(n1803[9]), .I2(GND_net), 
            .I3(n38332), .O(n1802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_12 (.CI(n38332), .I0(n1803[9]), .I1(GND_net), 
            .CO(n38333));
    SB_CARRY add_3225_13 (.CI(n36961), .I0(n11996[10]), .I1(GND_net), 
            .CO(n36962));
    SB_LUT4 add_3225_12_lut (.I0(GND_net), .I1(n11996[9]), .I2(GND_net), 
            .I3(n36960), .O(n11362[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n37505), .O(n82[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_12_lut (.I0(GND_net), .I1(n8352[9]), .I2(GND_net), 
            .I3(n37984), .O(n8335[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1049_add_4_9  (.CI(n37505), .I0(\PID_CONTROLLER.err[7] ), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n37506));
    SB_CARRY add_3225_12 (.CI(n36960), .I0(n11996[9]), .I1(GND_net), .CO(n36961));
    SB_LUT4 add_3225_11_lut (.I0(GND_net), .I1(n11996[8]), .I2(GND_net), 
            .I3(n36959), .O(n11362[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_24 (.CI(n36715), .I0(n282[22]), .I1(n76[22]), 
            .CO(n36716));
    SB_CARRY add_3099_12 (.CI(n37984), .I0(n8352[9]), .I1(GND_net), .CO(n37985));
    SB_LUT4 add_13_add_1_22497_add_1_23_lut (.I0(GND_net), .I1(n282[21]), 
            .I2(n76[21]), .I3(n36714), .O(n79[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n37504), .O(n82[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_11 (.CI(n36959), .I0(n11996[8]), .I1(GND_net), .CO(n36960));
    SB_LUT4 add_3099_11_lut (.I0(GND_net), .I1(n8352[8]), .I2(GND_net), 
            .I3(n37983), .O(n8335[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1049_add_4_8  (.CI(n37504), .I0(\PID_CONTROLLER.err[6] ), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n37505));
    SB_CARRY add_3099_11 (.CI(n37983), .I0(n8352[8]), .I1(GND_net), .CO(n37984));
    SB_LUT4 mult_14_add_1217_11_lut (.I0(GND_net), .I1(n1803[8]), .I2(GND_net), 
            .I3(n38331), .O(n1802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n37503), .O(n82[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_10_lut (.I0(GND_net), .I1(n11996[7]), .I2(GND_net), 
            .I3(n36958), .O(n11362[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_10 (.CI(n36958), .I0(n11996[7]), .I1(GND_net), .CO(n36959));
    SB_CARRY mult_14_add_1217_11 (.CI(n38331), .I0(n1803[8]), .I1(GND_net), 
            .CO(n38332));
    SB_LUT4 add_3099_10_lut (.I0(GND_net), .I1(n8352[7]), .I2(GND_net), 
            .I3(n37982), .O(n8335[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_10 (.CI(n37982), .I0(n8352[7]), .I1(GND_net), .CO(n37983));
    SB_CARRY \PID_CONTROLLER.integral_1049_add_4_7  (.CI(n37503), .I0(\PID_CONTROLLER.err[5] ), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n37504));
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n37502), .O(n82[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1049_add_4_6  (.CI(n37502), .I0(\PID_CONTROLLER.err[4] ), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n37503));
    SB_LUT4 add_3099_9_lut (.I0(GND_net), .I1(n8352[6]), .I2(GND_net), 
            .I3(n37981), .O(n8335[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n37501), .O(n82[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_9_lut (.I0(GND_net), .I1(n11996[6]), .I2(GND_net), 
            .I3(n36957), .O(n11362[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1049_add_4_5  (.CI(n37501), .I0(\PID_CONTROLLER.err[3] ), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n37502));
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n37500), .O(n82[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_23 (.CI(n36714), .I0(n282[21]), .I1(n76[21]), 
            .CO(n36715));
    SB_LUT4 add_13_add_1_22497_add_1_22_lut (.I0(GND_net), .I1(n282[20]), 
            .I2(n76[20]), .I3(n36713), .O(n79[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_9 (.CI(n37981), .I0(n8352[6]), .I1(GND_net), .CO(n37982));
    SB_CARRY add_3225_9 (.CI(n36957), .I0(n11996[6]), .I1(GND_net), .CO(n36958));
    SB_CARRY \PID_CONTROLLER.integral_1049_add_4_4  (.CI(n37500), .I0(\PID_CONTROLLER.err[2] ), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n37501));
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n37499), .O(n82[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_10_lut (.I0(GND_net), .I1(n1803[7]), .I2(GND_net), 
            .I3(n38330), .O(n1802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1049_add_4_3  (.CI(n37499), .I0(\PID_CONTROLLER.err[1] ), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n37500));
    SB_LUT4 add_3225_8_lut (.I0(GND_net), .I1(n11996[5]), .I2(n698_adj_3737), 
            .I3(n36956), .O(n11362[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_10 (.CI(n38330), .I0(n1803[7]), .I1(GND_net), 
            .CO(n38331));
    SB_LUT4 add_3099_8_lut (.I0(GND_net), .I1(n8352[5]), .I2(n728_adj_3738), 
            .I3(n37980), .O(n8335[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_9_lut (.I0(GND_net), .I1(n1803[6]), .I2(GND_net), 
            .I3(n38329), .O(n1802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_8 (.CI(n37980), .I0(n8352[5]), .I1(n728_adj_3738), 
            .CO(n37981));
    SB_LUT4 \PID_CONTROLLER.integral_1049_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n82[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1049_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1049_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err[0] ), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n37499));
    SB_CARRY add_3225_8 (.CI(n36956), .I0(n11996[5]), .I1(n698_adj_3737), 
            .CO(n36957));
    SB_LUT4 add_3099_7_lut (.I0(GND_net), .I1(n8352[4]), .I2(n631_adj_3740), 
            .I3(n37979), .O(n8335[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1048_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_count[8] ), 
            .I3(n37498), .O(n75[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1048_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_7_lut (.I0(GND_net), .I1(n11996[4]), .I2(n601_adj_3741), 
            .I3(n36955), .O(n11362[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1048_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_count[7] ), 
            .I3(n37497), .O(n75[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1048_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_7 (.CI(n36955), .I0(n11996[4]), .I1(n601_adj_3741), 
            .CO(n36956));
    SB_CARRY add_13_add_1_22497_add_1_22 (.CI(n36713), .I0(n282[20]), .I1(n76[20]), 
            .CO(n36714));
    SB_CARRY pwm_count_1048_add_4_9 (.CI(n37497), .I0(GND_net), .I1(\pwm_count[7] ), 
            .CO(n37498));
    SB_LUT4 add_13_add_1_22497_add_1_21_lut (.I0(GND_net), .I1(n282[19]), 
            .I2(n76[19]), .I3(n36712), .O(n79[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_6_lut (.I0(GND_net), .I1(n11996[3]), .I2(n504_adj_3743), 
            .I3(n36954), .O(n11362[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1048_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_count[6] ), 
            .I3(n37496), .O(n75[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1048_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_6 (.CI(n36954), .I0(n11996[3]), .I1(n504_adj_3743), 
            .CO(n36955));
    SB_LUT4 add_3225_5_lut (.I0(GND_net), .I1(n11996[2]), .I2(n407_adj_3745), 
            .I3(n36953), .O(n11362[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_9 (.CI(n38329), .I0(n1803[6]), .I1(GND_net), 
            .CO(n38330));
    SB_CARRY add_3099_7 (.CI(n37979), .I0(n8352[4]), .I1(n631_adj_3740), 
            .CO(n37980));
    SB_CARRY pwm_count_1048_add_4_8 (.CI(n37496), .I0(GND_net), .I1(\pwm_count[6] ), 
            .CO(n37497));
    SB_CARRY add_3225_5 (.CI(n36953), .I0(n11996[2]), .I1(n407_adj_3745), 
            .CO(n36954));
    SB_LUT4 mult_14_add_1217_8_lut (.I0(GND_net), .I1(n1803[5]), .I2(n530), 
            .I3(n38328), .O(n1802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_21 (.CI(n36712), .I0(n282[19]), .I1(n76[19]), 
            .CO(n36713));
    SB_LUT4 add_13_add_1_22497_add_1_20_lut (.I0(GND_net), .I1(n282[18]), 
            .I2(n76[18]), .I3(n36711), .O(n79[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_4_lut (.I0(GND_net), .I1(n11996[1]), .I2(n310_adj_3747), 
            .I3(n36952), .O(n11362[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1048_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_count[5] ), 
            .I3(n37495), .O(n75[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1048_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1048_add_4_7 (.CI(n37495), .I0(GND_net), .I1(\pwm_count[5] ), 
            .CO(n37496));
    SB_CARRY add_3225_4 (.CI(n36952), .I0(n11996[1]), .I1(n310_adj_3747), 
            .CO(n36953));
    SB_CARRY add_13_add_1_22497_add_1_20 (.CI(n36711), .I0(n282[18]), .I1(n76[18]), 
            .CO(n36712));
    SB_LUT4 add_13_add_1_22497_add_1_19_lut (.I0(GND_net), .I1(n282[17]), 
            .I2(n76[17]), .I3(n36710), .O(n79[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1048_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_count[4] ), 
            .I3(n37494), .O(n75[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1048_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_3_lut (.I0(GND_net), .I1(n11996[0]), .I2(n213_adj_3750), 
            .I3(n36951), .O(n11362[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_3 (.CI(n36951), .I0(n11996[0]), .I1(n213_adj_3750), 
            .CO(n36952));
    SB_CARRY add_13_add_1_22497_add_1_19 (.CI(n36710), .I0(n282[17]), .I1(n76[17]), 
            .CO(n36711));
    SB_CARRY pwm_count_1048_add_4_6 (.CI(n37494), .I0(GND_net), .I1(\pwm_count[4] ), 
            .CO(n37495));
    SB_LUT4 pwm_count_1048_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_count[3] ), 
            .I3(n37493), .O(n75[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1048_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_8 (.CI(n38328), .I0(n1803[5]), .I1(n530), 
            .CO(n38329));
    SB_LUT4 add_3099_6_lut (.I0(GND_net), .I1(n8352[3]), .I2(n534_adj_3752), 
            .I3(n37978), .O(n8335[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_6 (.CI(n37978), .I0(n8352[3]), .I1(n534_adj_3752), 
            .CO(n37979));
    SB_CARRY pwm_count_1048_add_4_5 (.CI(n37493), .I0(GND_net), .I1(\pwm_count[3] ), 
            .CO(n37494));
    SB_LUT4 add_3225_2_lut (.I0(GND_net), .I1(n23_adj_3753), .I2(n116_adj_3754), 
            .I3(GND_net), .O(n11362[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i28_2_lut (.I0(\Kd[0] ), .I1(n67[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_13_add_1_22497_add_1_18_lut (.I0(GND_net), .I1(n282[16]), 
            .I2(n76[16]), .I3(n36709), .O(n79[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_2 (.CI(GND_net), .I0(n23_adj_3753), .I1(n116_adj_3754), 
            .CO(n36951));
    SB_LUT4 pwm_count_1048_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_count[2] ), 
            .I3(n37492), .O(n75[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1048_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_11_lut (.I0(GND_net), .I1(n15230[8]), .I2(GND_net), 
            .I3(n36950), .O(n14916[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_5_lut (.I0(GND_net), .I1(n8352[2]), .I2(n437_adj_3756), 
            .I3(n37977), .O(n8335[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_10_lut (.I0(GND_net), .I1(n15230[7]), .I2(GND_net), 
            .I3(n36949), .O(n14916[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_5 (.CI(n37977), .I0(n8352[2]), .I1(n437_adj_3756), 
            .CO(n37978));
    SB_LUT4 mult_12_i154_2_lut (.I0(\Kd[2] ), .I1(n67[11]), .I2(GND_net), 
            .I3(GND_net), .O(n228));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i154_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY pwm_count_1048_add_4_4 (.CI(n37492), .I0(GND_net), .I1(\pwm_count[2] ), 
            .CO(n37493));
    SB_CARRY add_3389_10 (.CI(n36949), .I0(n15230[7]), .I1(GND_net), .CO(n36950));
    SB_LUT4 add_3389_9_lut (.I0(GND_net), .I1(n15230[6]), .I2(GND_net), 
            .I3(n36948), .O(n14916[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_9 (.CI(n36948), .I0(n15230[6]), .I1(GND_net), .CO(n36949));
    SB_LUT4 pwm_count_1048_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_count[1] ), 
            .I3(n37491), .O(n75[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1048_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_18 (.CI(n36709), .I0(n282[16]), .I1(n76[16]), 
            .CO(n36710));
    SB_CARRY pwm_count_1048_add_4_3 (.CI(n37491), .I0(GND_net), .I1(\pwm_count[1] ), 
            .CO(n37492));
    SB_LUT4 add_3389_8_lut (.I0(GND_net), .I1(n15230[5]), .I2(n545), .I3(n36947), 
            .O(n14916[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_4_lut (.I0(GND_net), .I1(n8352[1]), .I2(n340_adj_3758), 
            .I3(n37976), .O(n8335[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1048_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[0]), 
            .I3(VCC_net), .O(n75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1048_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_4 (.CI(n37976), .I0(n8352[1]), .I1(n340_adj_3758), 
            .CO(n37977));
    SB_CARRY add_3389_8 (.CI(n36947), .I0(n15230[5]), .I1(n545), .CO(n36948));
    SB_LUT4 add_3389_7_lut (.I0(GND_net), .I1(n15230[4]), .I2(n472), .I3(n36946), 
            .O(n14916[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_17_lut (.I0(GND_net), .I1(n282[15]), 
            .I2(n76[15]), .I3(n36708), .O(n79[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_17 (.CI(n36708), .I0(n282[15]), .I1(n76[15]), 
            .CO(n36709));
    SB_CARRY pwm_count_1048_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_count[0]), 
            .CO(n37491));
    SB_CARRY add_3389_7 (.CI(n36946), .I0(n15230[4]), .I1(n472), .CO(n36947));
    SB_LUT4 mult_14_add_1217_7_lut (.I0(GND_net), .I1(n1803[4]), .I2(n457_c), 
            .I3(n38327), .O(n1802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_3_lut (.I0(GND_net), .I1(n8352[0]), .I2(n243_adj_3760), 
            .I3(n37975), .O(n8335[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_31_lut (.I0(GND_net), .I1(n7992[28]), .I2(GND_net), 
            .I3(n37490), .O(n7960[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_6_lut (.I0(GND_net), .I1(n15230[3]), .I2(n399), .I3(n36945), 
            .O(n14916[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_6 (.CI(n36945), .I0(n15230[3]), .I1(n399), .CO(n36946));
    SB_LUT4 add_13_add_1_22497_add_1_16_lut (.I0(GND_net), .I1(n282[14]), 
            .I2(n76[14]), .I3(n36707), .O(n79[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_5_lut (.I0(GND_net), .I1(n15230[2]), .I2(n326), .I3(n36944), 
            .O(n14916[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i2  (.Q(\PID_CONTROLLER.err_prev[1] ), 
           .C(clk32MHz), .D(n23966));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_13_add_1_22497_add_1_16 (.CI(n36707), .I0(n282[14]), .I1(n76[14]), 
            .CO(n36708));
    SB_DFF \PID_CONTROLLER.err_prev__i3  (.Q(\PID_CONTROLLER.err_prev[2] ), 
           .C(clk32MHz), .D(n23965));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3084_30_lut (.I0(GND_net), .I1(n7992[27]), .I2(GND_net), 
            .I3(n37489), .O(n7960[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_30_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i4  (.Q(\PID_CONTROLLER.err_prev[3] ), 
           .C(clk32MHz), .D(n23964));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3099_3 (.CI(n37975), .I0(n8352[0]), .I1(n243_adj_3760), 
            .CO(n37976));
    SB_CARRY add_3084_30 (.CI(n37489), .I0(n7992[27]), .I1(GND_net), .CO(n37490));
    SB_DFF \PID_CONTROLLER.err_prev__i5  (.Q(\PID_CONTROLLER.err_prev[4] ), 
           .C(clk32MHz), .D(n23963));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3084_29_lut (.I0(GND_net), .I1(n7992[26]), .I2(GND_net), 
            .I3(n37488), .O(n7960[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_29_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i6  (.Q(\PID_CONTROLLER.err_prev[5] ), 
           .C(clk32MHz), .D(n23962));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i7  (.Q(\PID_CONTROLLER.err_prev[6] ), 
           .C(clk32MHz), .D(n23961));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3084_29 (.CI(n37488), .I0(n7992[26]), .I1(GND_net), .CO(n37489));
    SB_DFF \PID_CONTROLLER.err_prev__i8  (.Q(\PID_CONTROLLER.err_prev[7] ), 
           .C(clk32MHz), .D(n23960));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3389_5 (.CI(n36944), .I0(n15230[2]), .I1(n326), .CO(n36945));
    SB_DFF \PID_CONTROLLER.err_prev__i9  (.Q(\PID_CONTROLLER.err_prev[8] ), 
           .C(clk32MHz), .D(n23959));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3389_4_lut (.I0(GND_net), .I1(n15230[1]), .I2(n253), .I3(n36943), 
            .O(n14916[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i10  (.Q(\PID_CONTROLLER.err_prev[9] ), 
           .C(clk32MHz), .D(n23958));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3389_4 (.CI(n36943), .I0(n15230[1]), .I1(n253), .CO(n36944));
    SB_DFF \PID_CONTROLLER.err_prev__i11  (.Q(\PID_CONTROLLER.err_prev[10] ), 
           .C(clk32MHz), .D(n23957));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY mult_14_add_1217_7 (.CI(n38327), .I0(n1803[4]), .I1(n457_c), 
            .CO(n38328));
    SB_LUT4 add_3099_2_lut (.I0(GND_net), .I1(n53_adj_3761), .I2(n146_adj_3762), 
            .I3(GND_net), .O(n8335[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i12  (.Q(\PID_CONTROLLER.err_prev[11] ), 
           .C(clk32MHz), .D(n23956));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3084_28_lut (.I0(GND_net), .I1(n7992[25]), .I2(GND_net), 
            .I3(n37487), .O(n7960[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_28_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i13  (.Q(\PID_CONTROLLER.err_prev[12] ), 
           .C(clk32MHz), .D(n23955));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3389_3_lut (.I0(GND_net), .I1(n15230[0]), .I2(n180_adj_3552), 
            .I3(n36942), .O(n14916[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i14  (.Q(\PID_CONTROLLER.err_prev[13] ), 
           .C(clk32MHz), .D(n23954));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3389_3 (.CI(n36942), .I0(n15230[0]), .I1(n180_adj_3552), 
            .CO(n36943));
    SB_DFF \PID_CONTROLLER.err_prev__i15  (.Q(\PID_CONTROLLER.err_prev[14] ), 
           .C(clk32MHz), .D(n23953));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3084_28 (.CI(n37487), .I0(n7992[25]), .I1(GND_net), .CO(n37488));
    SB_DFF \PID_CONTROLLER.err_prev__i16  (.Q(\PID_CONTROLLER.err_prev[15] ), 
           .C(clk32MHz), .D(n23952));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3084_27_lut (.I0(GND_net), .I1(n7992[24]), .I2(GND_net), 
            .I3(n37486), .O(n7960[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_27_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i17  (.Q(\PID_CONTROLLER.err_prev[16] ), 
           .C(clk32MHz), .D(n23951));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i18  (.Q(\PID_CONTROLLER.err_prev[17] ), 
           .C(clk32MHz), .D(n23950));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i19  (.Q(\PID_CONTROLLER.err_prev[18] ), 
           .C(clk32MHz), .D(n23949));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3389_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n14916[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i20  (.Q(\PID_CONTROLLER.err_prev[19] ), 
           .C(clk32MHz), .D(n23948));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_13_add_1_22497_add_1_15_lut (.I0(GND_net), .I1(n282[13]), 
            .I2(n76[13]), .I3(n36706), .O(n79[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i21  (.Q(\PID_CONTROLLER.err_prev[20] ), 
           .C(clk32MHz), .D(n23947));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3389_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n36942));
    SB_DFF \PID_CONTROLLER.err_prev__i22  (.Q(\PID_CONTROLLER.err_prev[21] ), 
           .C(clk32MHz), .D(n23946));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 mult_14_add_1217_6_lut (.I0(GND_net), .I1(n1803[3]), .I2(n384), 
            .I3(n38326), .O(n1802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_2 (.CI(GND_net), .I0(n53_adj_3761), .I1(n146_adj_3762), 
            .CO(n37975));
    SB_CARRY add_13_add_1_22497_add_1_15 (.CI(n36706), .I0(n282[13]), .I1(n76[13]), 
            .CO(n36707));
    SB_DFF \PID_CONTROLLER.err_prev__i23  (.Q(\PID_CONTROLLER.err_prev[22] ), 
           .C(clk32MHz), .D(n23945));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i24  (.Q(\PID_CONTROLLER.err_prev[23] ), 
           .C(clk32MHz), .D(n23944));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3098_17_lut (.I0(GND_net), .I1(n8335[14]), .I2(GND_net), 
            .I3(n37974), .O(n8317[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i25  (.Q(\PID_CONTROLLER.err_prev[31] ), 
           .C(clk32MHz), .D(n23943));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3084_27 (.CI(n37486), .I0(n7992[24]), .I1(GND_net), .CO(n37487));
    SB_LUT4 add_3098_16_lut (.I0(GND_net), .I1(n8335[13]), .I2(GND_net), 
            .I3(n37973), .O(n8317[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_26_lut (.I0(GND_net), .I1(n7992[23]), .I2(GND_net), 
            .I3(n37485), .O(n7960[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_16 (.CI(n37973), .I0(n8335[13]), .I1(GND_net), .CO(n37974));
    SB_CARRY add_3084_26 (.CI(n37485), .I0(n7992[23]), .I1(GND_net), .CO(n37486));
    SB_LUT4 add_3084_25_lut (.I0(GND_net), .I1(n7992[22]), .I2(GND_net), 
            .I3(n37484), .O(n7960[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_25 (.CI(n37484), .I0(n7992[22]), .I1(GND_net), .CO(n37485));
    SB_LUT4 add_3084_24_lut (.I0(GND_net), .I1(n7992[21]), .I2(GND_net), 
            .I3(n37483), .O(n7960[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_24 (.CI(n37483), .I0(n7992[21]), .I1(GND_net), .CO(n37484));
    SB_LUT4 add_13_add_1_22497_add_1_14_lut (.I0(GND_net), .I1(n282[12]), 
            .I2(n76[12]), .I3(n36705), .O(n79[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_23_lut (.I0(GND_net), .I1(n7992[20]), .I2(GND_net), 
            .I3(n37482), .O(n7960[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_6 (.CI(n38326), .I0(n1803[3]), .I1(n384), 
            .CO(n38327));
    SB_CARRY add_3084_23 (.CI(n37482), .I0(n7992[20]), .I1(GND_net), .CO(n37483));
    SB_DFF \PID_CONTROLLER.result_i1  (.Q(\PID_CONTROLLER.result [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [1]));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_13_add_1_22497_add_1_14 (.CI(n36705), .I0(n282[12]), .I1(n76[12]), 
            .CO(n36706));
    SB_LUT4 add_3098_15_lut (.I0(GND_net), .I1(n8335[12]), .I2(GND_net), 
            .I3(n37972), .O(n8317[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_22_lut (.I0(GND_net), .I1(n7992[19]), .I2(GND_net), 
            .I3(n37481), .O(n7960[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_5_lut (.I0(GND_net), .I1(n1803[2]), .I2(n311_adj_3764), 
            .I3(n38325), .O(n1802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_5 (.CI(n38325), .I0(n1803[2]), .I1(n311_adj_3764), 
            .CO(n38326));
    SB_CARRY add_3098_15 (.CI(n37972), .I0(n8335[12]), .I1(GND_net), .CO(n37973));
    SB_CARRY add_3084_22 (.CI(n37481), .I0(n7992[19]), .I1(GND_net), .CO(n37482));
    SB_LUT4 add_3084_21_lut (.I0(GND_net), .I1(n7992[18]), .I2(GND_net), 
            .I3(n37480), .O(n7960[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.result_i2  (.Q(\PID_CONTROLLER.result [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [2]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i3  (.Q(\PID_CONTROLLER.result [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [3]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i4  (.Q(\PID_CONTROLLER.result[4] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [4]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i5  (.Q(\PID_CONTROLLER.result[5] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [5]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i6  (.Q(\PID_CONTROLLER.result [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [6]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i7  (.Q(\PID_CONTROLLER.result[7] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [7]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i8  (.Q(\PID_CONTROLLER.result [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [8]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i9  (.Q(\PID_CONTROLLER.result [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [9]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i10  (.Q(\PID_CONTROLLER.result [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [10]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i11  (.Q(\PID_CONTROLLER.result [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [11]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i12  (.Q(\PID_CONTROLLER.result [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [12]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i13  (.Q(\PID_CONTROLLER.result [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [13]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i14  (.Q(\PID_CONTROLLER.result [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [14]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i15  (.Q(\PID_CONTROLLER.result [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [15]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i16  (.Q(\PID_CONTROLLER.result [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [16]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i17  (.Q(\PID_CONTROLLER.result [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [17]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i18  (.Q(\PID_CONTROLLER.result [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [18]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i19  (.Q(\PID_CONTROLLER.result [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [19]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i20  (.Q(\PID_CONTROLLER.result [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [20]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i21  (.Q(\PID_CONTROLLER.result [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [21]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i22  (.Q(\PID_CONTROLLER.result [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [22]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i23  (.Q(\PID_CONTROLLER.result [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [23]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i24  (.Q(\PID_CONTROLLER.result [24]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [24]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i25  (.Q(\PID_CONTROLLER.result [25]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [25]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i26  (.Q(\PID_CONTROLLER.result [26]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [26]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i27  (.Q(\PID_CONTROLLER.result [27]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [27]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i28  (.Q(\PID_CONTROLLER.result [28]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [28]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i29  (.Q(\PID_CONTROLLER.result [29]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [29]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i30  (.Q(\PID_CONTROLLER.result [30]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [30]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i31  (.Q(\PID_CONTROLLER.result [31]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [31]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err[1] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [1]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFFE PHASES_i1 (.Q(PIN_6_c_0), .C(clk32MHz), .E(n23562), .D(PHASES_5__N_2779[0]));   // verilog/motorControl.v(57[10] 100[6])
    SB_DFFE PHASES_i2 (.Q(PIN_5_c_1), .C(clk32MHz), .E(n23622), .D(PHASES_5__N_2779[1]));   // verilog/motorControl.v(57[10] 100[6])
    SB_DFFE PHASES_i3 (.Q(PIN_4_c_2), .C(clk32MHz), .E(n15_adj_3765), 
            .D(PHASES_5__N_2779[2]));   // verilog/motorControl.v(57[10] 100[6])
    SB_DFFE PHASES_i4 (.Q(PIN_3_c_3), .C(clk32MHz), .E(n23630), .D(PHASES_5__N_2779[3]));   // verilog/motorControl.v(57[10] 100[6])
    SB_DFFE PHASES_i5 (.Q(PIN_2_c_4), .C(clk32MHz), .E(n42681), .D(PHASES_5__N_2779[4]));   // verilog/motorControl.v(57[10] 100[6])
    SB_LUT4 add_13_add_1_22497_add_1_13_lut (.I0(GND_net), .I1(n282[11]), 
            .I2(n76[11]), .I3(n36704), .O(n79[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_14_lut (.I0(GND_net), .I1(n8335[11]), .I2(GND_net), 
            .I3(n37971), .O(n8317[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_21 (.CI(n37480), .I0(n7992[18]), .I1(GND_net), .CO(n37481));
    SB_LUT4 add_3251_25_lut (.I0(GND_net), .I1(n12579[22]), .I2(GND_net), 
            .I3(n36935), .O(n11996[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_13 (.CI(n36704), .I0(n282[11]), .I1(n76[11]), 
            .CO(n36705));
    SB_LUT4 add_3251_24_lut (.I0(GND_net), .I1(n12579[21]), .I2(GND_net), 
            .I3(n36934), .O(n11996[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_12_lut (.I0(GND_net), .I1(n282[10]), 
            .I2(n76[10]), .I3(n36703), .O(n79[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_12 (.CI(n36703), .I0(n282[10]), .I1(n76[10]), 
            .CO(n36704));
    SB_LUT4 add_3084_20_lut (.I0(GND_net), .I1(n7992[17]), .I2(GND_net), 
            .I3(n37479), .O(n7960[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_4_lut (.I0(GND_net), .I1(n1803[1]), .I2(n238_adj_3767), 
            .I3(n38324), .O(n1802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_14 (.CI(n37971), .I0(n8335[11]), .I1(GND_net), .CO(n37972));
    SB_CARRY add_3084_20 (.CI(n37479), .I0(n7992[17]), .I1(GND_net), .CO(n37480));
    SB_CARRY add_3251_24 (.CI(n36934), .I0(n12579[21]), .I1(GND_net), 
            .CO(n36935));
    SB_LUT4 add_3251_23_lut (.I0(GND_net), .I1(n12579[20]), .I2(GND_net), 
            .I3(n36933), .O(n11996[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_23 (.CI(n36933), .I0(n12579[20]), .I1(GND_net), 
            .CO(n36934));
    SB_LUT4 add_3251_22_lut (.I0(GND_net), .I1(n12579[19]), .I2(GND_net), 
            .I3(n36932), .O(n11996[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_4 (.CI(n38324), .I0(n1803[1]), .I1(n238_adj_3767), 
            .CO(n38325));
    SB_LUT4 add_3098_13_lut (.I0(GND_net), .I1(n8335[10]), .I2(GND_net), 
            .I3(n37970), .O(n8317[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_19_lut (.I0(GND_net), .I1(n7992[16]), .I2(GND_net), 
            .I3(n37478), .O(n7960[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_22 (.CI(n36932), .I0(n12579[19]), .I1(GND_net), 
            .CO(n36933));
    SB_LUT4 add_13_add_1_22497_add_1_11_lut (.I0(GND_net), .I1(n282[9]), 
            .I2(n76[9]), .I3(n36702), .O(n79[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_21_lut (.I0(GND_net), .I1(n12579[18]), .I2(GND_net), 
            .I3(n36931), .O(n11996[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_13 (.CI(n37970), .I0(n8335[10]), .I1(GND_net), .CO(n37971));
    SB_CARRY add_3084_19 (.CI(n37478), .I0(n7992[16]), .I1(GND_net), .CO(n37479));
    SB_CARRY add_3251_21 (.CI(n36931), .I0(n12579[18]), .I1(GND_net), 
            .CO(n36932));
    SB_LUT4 add_3251_20_lut (.I0(GND_net), .I1(n12579[17]), .I2(GND_net), 
            .I3(n36930), .O(n11996[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_11 (.CI(n36702), .I0(n282[9]), .I1(n76[9]), 
            .CO(n36703));
    SB_LUT4 add_13_add_1_22497_add_1_10_lut (.I0(GND_net), .I1(n282[8]), 
            .I2(n76[8]), .I3(n36701), .O(n79[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_3_lut (.I0(GND_net), .I1(n1803[0]), .I2(n165_adj_3769), 
            .I3(n38323), .O(n1802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_12_lut (.I0(GND_net), .I1(n8335[9]), .I2(GND_net), 
            .I3(n37969), .O(n8317[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_10 (.CI(n36701), .I0(n282[8]), .I1(n76[8]), 
            .CO(n36702));
    SB_LUT4 add_3084_18_lut (.I0(GND_net), .I1(n7992[15]), .I2(GND_net), 
            .I3(n37477), .O(n7960[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_18 (.CI(n37477), .I0(n7992[15]), .I1(GND_net), .CO(n37478));
    SB_CARRY add_3251_20 (.CI(n36930), .I0(n12579[17]), .I1(GND_net), 
            .CO(n36931));
    SB_LUT4 add_3251_19_lut (.I0(GND_net), .I1(n12579[16]), .I2(GND_net), 
            .I3(n36929), .O(n11996[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_19 (.CI(n36929), .I0(n12579[16]), .I1(GND_net), 
            .CO(n36930));
    SB_CARRY add_3098_12 (.CI(n37969), .I0(n8335[9]), .I1(GND_net), .CO(n37970));
    SB_LUT4 add_3084_17_lut (.I0(GND_net), .I1(n7992[14]), .I2(GND_net), 
            .I3(n37476), .O(n7960[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_18_lut (.I0(GND_net), .I1(n12579[15]), .I2(GND_net), 
            .I3(n36928), .O(n11996[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_18 (.CI(n36928), .I0(n12579[15]), .I1(GND_net), 
            .CO(n36929));
    SB_LUT4 add_3098_11_lut (.I0(GND_net), .I1(n8335[8]), .I2(GND_net), 
            .I3(n37968), .O(n8317[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_9_lut (.I0(GND_net), .I1(n282[7]), 
            .I2(n76[7]), .I3(n36700), .O(n79[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n6_adj_3771), 
            .I3(n36574), .O(n58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_17_lut (.I0(GND_net), .I1(n12579[14]), .I2(GND_net), 
            .I3(n36927), .O(n11996[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_9 (.CI(n36700), .I0(n282[7]), .I1(n76[7]), 
            .CO(n36701));
    SB_CARRY add_3084_17 (.CI(n37476), .I0(n7992[14]), .I1(GND_net), .CO(n37477));
    SB_CARRY mult_14_add_1217_3 (.CI(n38323), .I0(n1803[0]), .I1(n165_adj_3769), 
            .CO(n38324));
    SB_CARRY add_3098_11 (.CI(n37968), .I0(n8335[8]), .I1(GND_net), .CO(n37969));
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err[2] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [2]));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3084_16_lut (.I0(GND_net), .I1(n7992[13]), .I2(GND_net), 
            .I3(n37475), .O(n7960[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_17 (.CI(n36927), .I0(n12579[14]), .I1(GND_net), 
            .CO(n36928));
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err[3] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [3]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err[4] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [4]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err[5] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [5]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err[6] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [6]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err[7] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [7]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err[8] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [8]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err[9] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [9]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err[10] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [10]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err[11] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [11]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err[12] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [12]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err[13] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [13]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err[14] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [14]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err[15] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [15]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err[16] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [16]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err[17] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [17]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err[18] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [18]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err[19] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [19]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err[20] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [20]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err[21] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [21]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err[22] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [22]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i24  (.Q(\PID_CONTROLLER.err[23] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [23]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i25  (.Q(\PID_CONTROLLER.err[31] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [24]));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3251_16_lut (.I0(GND_net), .I1(n12579[13]), .I2(GND_net), 
            .I3(n36926), .O(n11996[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_16 (.CI(n37475), .I0(n7992[13]), .I1(GND_net), .CO(n37476));
    SB_CARRY add_3251_16 (.CI(n36926), .I0(n12579[13]), .I1(GND_net), 
            .CO(n36927));
    SB_LUT4 add_3098_10_lut (.I0(GND_net), .I1(n8335[7]), .I2(GND_net), 
            .I3(n37967), .O(n8317[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_15_lut (.I0(GND_net), .I1(n7992[12]), .I2(GND_net), 
            .I3(n37474), .O(n7960[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_15_lut (.I0(GND_net), .I1(n12579[12]), .I2(GND_net), 
            .I3(n36925), .O(n11996[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_8_lut (.I0(GND_net), .I1(n282[6]), 
            .I2(n76[6]), .I3(n36699), .O(n79[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n6_adj_3771), 
            .I3(n36573), .O(n58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_15 (.CI(n36925), .I0(n12579[12]), .I1(GND_net), 
            .CO(n36926));
    SB_LUT4 add_3251_14_lut (.I0(GND_net), .I1(n12579[11]), .I2(GND_net), 
            .I3(n36924), .O(n11996[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_14 (.CI(n36924), .I0(n12579[11]), .I1(GND_net), 
            .CO(n36925));
    SB_CARRY add_3098_10 (.CI(n37967), .I0(n8335[7]), .I1(GND_net), .CO(n37968));
    SB_CARRY add_13_add_1_22497_add_1_8 (.CI(n36699), .I0(n282[6]), .I1(n76[6]), 
            .CO(n36700));
    SB_LUT4 add_13_add_1_22497_add_1_7_lut (.I0(GND_net), .I1(n282[5]), 
            .I2(n76[5]), .I3(n36698), .O(n79[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_7 (.CI(n36698), .I0(n282[5]), .I1(n76[5]), 
            .CO(n36699));
    SB_CARRY add_3084_15 (.CI(n37474), .I0(n7992[12]), .I1(GND_net), .CO(n37475));
    SB_LUT4 add_3251_13_lut (.I0(GND_net), .I1(n12579[10]), .I2(GND_net), 
            .I3(n36923), .O(n11996[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_6_lut (.I0(GND_net), .I1(n282[4]), 
            .I2(n76[4]), .I3(n36697), .O(n79[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_13 (.CI(n36923), .I0(n12579[10]), .I1(GND_net), 
            .CO(n36924));
    SB_LUT4 add_3098_9_lut (.I0(GND_net), .I1(n8335[6]), .I2(GND_net), 
            .I3(n37966), .O(n8317[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_9 (.CI(n37966), .I0(n8335[6]), .I1(GND_net), .CO(n37967));
    SB_LUT4 mult_14_add_1217_2_lut (.I0(GND_net), .I1(n23_adj_3772), .I2(n92), 
            .I3(GND_net), .O(n1802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_2 (.CI(GND_net), .I0(n23_adj_3772), .I1(n92), 
            .CO(n38323));
    SB_LUT4 add_3084_14_lut (.I0(GND_net), .I1(n7992[11]), .I2(GND_net), 
            .I3(n37473), .O(n7960[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_12_lut (.I0(GND_net), .I1(n12579[9]), .I2(GND_net), 
            .I3(n36922), .O(n11996[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_6 (.CI(n36697), .I0(n282[4]), .I1(n76[4]), 
            .CO(n36698));
    SB_LUT4 mult_14_add_1216_24_lut (.I0(GND_net), .I1(n1802[21]), .I2(GND_net), 
            .I3(n38321), .O(n1801[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_14 (.CI(n37473), .I0(n7992[11]), .I1(GND_net), .CO(n37474));
    SB_CARRY add_3251_12 (.CI(n36922), .I0(n12579[9]), .I1(GND_net), .CO(n36923));
    SB_CARRY unary_minus_21_add_3_11 (.CI(n36573), .I0(GND_net), .I1(n6_adj_3771), 
            .CO(n36574));
    SB_CARRY mult_14_add_1216_24 (.CI(n38321), .I0(n1802[21]), .I1(GND_net), 
            .CO(n1703));
    SB_LUT4 mult_14_add_1216_23_lut (.I0(GND_net), .I1(n1802[20]), .I2(GND_net), 
            .I3(n38320), .O(n1801[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_8_lut (.I0(GND_net), .I1(n8335[5]), .I2(n725_adj_3773), 
            .I3(n37965), .O(n8317[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_13_lut (.I0(GND_net), .I1(n7992[10]), .I2(GND_net), 
            .I3(n37472), .O(n7960[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_11_lut (.I0(GND_net), .I1(n12579[8]), .I2(GND_net), 
            .I3(n36921), .O(n11996[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_11 (.CI(n36921), .I0(n12579[8]), .I1(GND_net), .CO(n36922));
    SB_CARRY add_3098_8 (.CI(n37965), .I0(n8335[5]), .I1(n725_adj_3773), 
            .CO(n37966));
    SB_CARRY add_3084_13 (.CI(n37472), .I0(n7992[10]), .I1(GND_net), .CO(n37473));
    SB_LUT4 add_3251_10_lut (.I0(GND_net), .I1(n12579[7]), .I2(GND_net), 
            .I3(n36920), .O(n11996[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_10 (.CI(n36920), .I0(n12579[7]), .I1(GND_net), .CO(n36921));
    SB_LUT4 add_3098_7_lut (.I0(GND_net), .I1(n8335[4]), .I2(n628_adj_3774), 
            .I3(n37964), .O(n8317[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_9_lut (.I0(GND_net), .I1(n12579[6]), .I2(GND_net), 
            .I3(n36919), .O(n11996[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27934_2_lut_3_lut (.I0(PHASES_5__N_3039[4]), .I1(hall3), .I2(PHASES_5__N_3039[3]), 
            .I3(GND_net), .O(n43441));   // verilog/motorControl.v(90[10:34])
    defparam i27934_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i2_3_lut_4_lut_adj_1384 (.I0(PHASES_5__N_3039[4]), .I1(hall3), 
            .I2(n934), .I3(PHASES_5__N_3039[3]), .O(n22379));   // verilog/motorControl.v(90[10:34])
    defparam i2_3_lut_4_lut_adj_1384.LUT_INIT = 16'hfff8;
    SB_CARRY add_3098_7 (.CI(n37964), .I0(n8335[4]), .I1(n628_adj_3774), 
            .CO(n37965));
    SB_LUT4 add_3084_12_lut (.I0(GND_net), .I1(n7992[9]), .I2(GND_net), 
            .I3(n37471), .O(n7960[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n61[8]), 
            .I3(n36572), .O(n58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_12 (.CI(n37471), .I0(n7992[9]), .I1(GND_net), .CO(n37472));
    SB_CARRY mult_14_add_1216_23 (.CI(n38320), .I0(n1802[20]), .I1(GND_net), 
            .CO(n38321));
    SB_LUT4 add_3084_11_lut (.I0(GND_net), .I1(n7992[8]), .I2(GND_net), 
            .I3(n37470), .O(n7960[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_9 (.CI(n36919), .I0(n12579[6]), .I1(GND_net), .CO(n36920));
    SB_CARRY add_3084_11 (.CI(n37470), .I0(n7992[8]), .I1(GND_net), .CO(n37471));
    SB_LUT4 i6310_3_lut_3_lut (.I0(PHASES_5__N_3039[4]), .I1(hall3), .I2(n19954), 
            .I3(GND_net), .O(n19616));   // verilog/motorControl.v(90[10:34])
    defparam i6310_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 mult_14_add_1216_22_lut (.I0(GND_net), .I1(n1802[19]), .I2(GND_net), 
            .I3(n38319), .O(n1801[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_10_lut (.I0(GND_net), .I1(n7992[7]), .I2(GND_net), 
            .I3(n37469), .O(n7960[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_8_lut (.I0(GND_net), .I1(n12579[5]), .I2(n701_adj_3776), 
            .I3(n36918), .O(n11996[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_5_lut (.I0(GND_net), .I1(n282[3]), 
            .I2(n76[3]), .I3(n36696), .O(n79[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1047__i1 (.Q(Kd_delay_counter[1]), .C(clk32MHz), 
           .D(n57[1]));   // verilog/motorControl.v(48[27:47])
    SB_LUT4 add_3098_6_lut (.I0(GND_net), .I1(n8335[3]), .I2(n531_adj_3777), 
            .I3(n37963), .O(n8317[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_5 (.CI(n36696), .I0(n282[3]), .I1(n76[3]), 
            .CO(n36697));
    SB_CARRY add_3084_10 (.CI(n37469), .I0(n7992[7]), .I1(GND_net), .CO(n37470));
    SB_CARRY mult_14_add_1216_22 (.CI(n38319), .I0(n1802[19]), .I1(GND_net), 
            .CO(n38320));
    SB_CARRY add_3098_6 (.CI(n37963), .I0(n8335[3]), .I1(n531_adj_3777), 
            .CO(n37964));
    SB_LUT4 add_3084_9_lut (.I0(GND_net), .I1(n7992[6]), .I2(GND_net), 
            .I3(n37468), .O(n7960[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_8 (.CI(n36918), .I0(n12579[5]), .I1(n701_adj_3776), 
            .CO(n36919));
    SB_LUT4 mult_12_i156_2_lut (.I0(\Kd[2] ), .I1(n67[12]), .I2(GND_net), 
            .I3(GND_net), .O(n231));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i221_2_lut (.I0(\Kd[3] ), .I1(n67[12]), .I2(GND_net), 
            .I3(GND_net), .O(n328));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i221_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_21_add_3_10 (.CI(n36572), .I0(GND_net), .I1(n61[8]), 
            .CO(n36573));
    SB_CARRY add_3084_9 (.CI(n37468), .I0(n7992[6]), .I1(GND_net), .CO(n37469));
    SB_LUT4 add_3251_7_lut (.I0(GND_net), .I1(n12579[4]), .I2(n604_adj_3778), 
            .I3(n36917), .O(n11996[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFE PHASES_i6 (.Q(PIN_1_c_5), .C(clk32MHz), .E(n42680), .D(PHASES_5__N_2779[5]));   // verilog/motorControl.v(57[10] 100[6])
    SB_LUT4 add_3084_8_lut (.I0(GND_net), .I1(n7992[5]), .I2(n683_adj_3779), 
            .I3(n37467), .O(n7960[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_7 (.CI(n36917), .I0(n12579[4]), .I1(n604_adj_3778), 
            .CO(n36918));
    SB_LUT4 add_3251_6_lut (.I0(GND_net), .I1(n12579[3]), .I2(n507_adj_3780), 
            .I3(n36916), .O(n11996[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_5_lut (.I0(GND_net), .I1(n8335[2]), .I2(n434_adj_3781), 
            .I3(n37962), .O(n8317[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_6 (.CI(n36916), .I0(n12579[3]), .I1(n507_adj_3780), 
            .CO(n36917));
    SB_LUT4 mult_14_add_1216_21_lut (.I0(GND_net), .I1(n1802[18]), .I2(GND_net), 
            .I3(n38318), .O(n1801[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_5_lut (.I0(GND_net), .I1(n12579[2]), .I2(n410_adj_3782), 
            .I3(n36915), .O(n11996[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_5 (.CI(n37962), .I0(n8335[2]), .I1(n434_adj_3781), 
            .CO(n37963));
    SB_LUT4 add_13_add_1_22497_add_1_4_lut (.I0(GND_net), .I1(n282[2]), 
            .I2(n76[2]), .I3(n36695), .O(n79[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_8 (.CI(n37467), .I0(n7992[5]), .I1(n683_adj_3779), 
            .CO(n37468));
    SB_CARRY add_3251_5 (.CI(n36915), .I0(n12579[2]), .I1(n410_adj_3782), 
            .CO(n36916));
    SB_CARRY mult_14_add_1216_21 (.CI(n38318), .I0(n1802[18]), .I1(GND_net), 
            .CO(n38319));
    SB_LUT4 add_3098_4_lut (.I0(GND_net), .I1(n8335[1]), .I2(n337_adj_3783), 
            .I3(n37961), .O(n8317[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_7_lut (.I0(GND_net), .I1(n7992[4]), .I2(n586_adj_3784), 
            .I3(n37466), .O(n7960[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_4_lut (.I0(GND_net), .I1(n12579[1]), .I2(n313_adj_3785), 
            .I3(n36914), .O(n11996[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_4 (.CI(n37961), .I0(n8335[1]), .I1(n337_adj_3783), 
            .CO(n37962));
    SB_CARRY add_3084_7 (.CI(n37466), .I0(n7992[4]), .I1(n586_adj_3784), 
            .CO(n37467));
    SB_CARRY add_3251_4 (.CI(n36914), .I0(n12579[1]), .I1(n313_adj_3785), 
            .CO(n36915));
    SB_LUT4 add_3084_6_lut (.I0(GND_net), .I1(n7992[3]), .I2(n489_adj_3786), 
            .I3(n37465), .O(n7960[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_3_lut (.I0(GND_net), .I1(n8335[0]), .I2(n240_adj_3787), 
            .I3(n37960), .O(n8317[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i219_2_lut (.I0(\Kd[3] ), .I1(n67[11]), .I2(GND_net), 
            .I3(GND_net), .O(n325));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i219_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3084_6 (.CI(n37465), .I0(n7992[3]), .I1(n489_adj_3786), 
            .CO(n37466));
    SB_LUT4 add_3251_3_lut (.I0(GND_net), .I1(n12579[0]), .I2(n216_adj_3788), 
            .I3(n36913), .O(n11996[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_3 (.CI(n37960), .I0(n8335[0]), .I1(n240_adj_3787), 
            .CO(n37961));
    SB_LUT4 mult_12_i284_2_lut (.I0(\Kd[4] ), .I1(n67[11]), .I2(GND_net), 
            .I3(GND_net), .O(n422));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i284_2_lut.LUT_INIT = 16'h8888;
    SB_DFF Kd_delay_counter_1047__i2 (.Q(Kd_delay_counter[2]), .C(clk32MHz), 
           .D(n57[2]));   // verilog/motorControl.v(48[27:47])
    SB_DFF Kd_delay_counter_1047__i3 (.Q(Kd_delay_counter[3]), .C(clk32MHz), 
           .D(n57[3]));   // verilog/motorControl.v(48[27:47])
    SB_DFF Kd_delay_counter_1047__i4 (.Q(Kd_delay_counter[4]), .C(clk32MHz), 
           .D(n57[4]));   // verilog/motorControl.v(48[27:47])
    SB_DFF Kd_delay_counter_1047__i5 (.Q(Kd_delay_counter[5]), .C(clk32MHz), 
           .D(n57[5]));   // verilog/motorControl.v(48[27:47])
    SB_DFF Kd_delay_counter_1047__i6 (.Q(Kd_delay_counter[6]), .C(clk32MHz), 
           .D(n57[6]));   // verilog/motorControl.v(48[27:47])
    SB_DFF pwm_count_1048__i1 (.Q(\pwm_count[1] ), .C(clk32MHz), .D(n75[1]));   // verilog/motorControl.v(99[18:29])
    SB_CARRY add_13_add_1_22497_add_1_4 (.CI(n36695), .I0(n282[2]), .I1(n76[2]), 
            .CO(n36696));
    SB_LUT4 add_3098_2_lut (.I0(GND_net), .I1(n50_adj_3790), .I2(n143_adj_3791), 
            .I3(GND_net), .O(n8317[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_3_lut (.I0(GND_net), .I1(n282[1]), 
            .I2(n76[1]), .I3(n36694), .O(n79[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_5_lut (.I0(GND_net), .I1(n7992[2]), .I2(n392_adj_3792), 
            .I3(n37464), .O(n7960[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_5 (.CI(n37464), .I0(n7992[2]), .I1(n392_adj_3792), 
            .CO(n37465));
    SB_CARRY add_3251_3 (.CI(n36913), .I0(n12579[0]), .I1(n216_adj_3788), 
            .CO(n36914));
    SB_CARRY add_13_add_1_22497_add_1_3 (.CI(n36694), .I0(n282[1]), .I1(n76[1]), 
            .CO(n36695));
    SB_LUT4 add_3251_2_lut (.I0(GND_net), .I1(n26_adj_3793), .I2(n119_adj_3794), 
            .I3(GND_net), .O(n11996[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22497_add_1_2_lut (.I0(GND_net), .I1(n282[0]), 
            .I2(n76[0]), .I3(GND_net), .O(n79[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22497_add_1_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_20_lut (.I0(GND_net), .I1(n1802[17]), .I2(GND_net), 
            .I3(n38317), .O(n1801[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_20 (.CI(n38317), .I0(n1802[17]), .I1(GND_net), 
            .CO(n38318));
    SB_CARRY add_3098_2 (.CI(GND_net), .I0(n50_adj_3790), .I1(n143_adj_3791), 
            .CO(n37960));
    SB_LUT4 add_3097_18_lut (.I0(GND_net), .I1(n8317[15]), .I2(GND_net), 
            .I3(n37959), .O(n8298[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_4_lut (.I0(GND_net), .I1(n7992[1]), .I2(n295_adj_3797), 
            .I3(n37463), .O(n7960[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_2 (.CI(GND_net), .I0(n26_adj_3793), .I1(n119_adj_3794), 
            .CO(n36913));
    SB_CARRY add_3084_4 (.CI(n37463), .I0(n7992[1]), .I1(n295_adj_3797), 
            .CO(n37464));
    SB_LUT4 add_3407_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(n36912), .O(n15230[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22497_add_1_2 (.CI(GND_net), .I0(n282[0]), .I1(n76[0]), 
            .CO(n36694));
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n61[7]), 
            .I3(n36571), .O(n413)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_9_lut (.I0(GND_net), .I1(n583_adj_3800), .I2(GND_net), 
            .I3(n36911), .O(n15230[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_17_lut (.I0(GND_net), .I1(n8317[14]), .I2(GND_net), 
            .I3(n37958), .O(n8298[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_3_lut (.I0(GND_net), .I1(n7992[0]), .I2(n198_adj_3801), 
            .I3(n37462), .O(n7960[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_9 (.CI(n36911), .I0(n583_adj_3800), .I1(GND_net), 
            .CO(n36912));
    SB_CARRY add_3084_3 (.CI(n37462), .I0(n7992[0]), .I1(n198_adj_3801), 
            .CO(n37463));
    SB_CARRY unary_minus_21_add_3_9 (.CI(n36571), .I0(GND_net), .I1(n61[7]), 
            .CO(n36572));
    SB_LUT4 add_3407_8_lut (.I0(GND_net), .I1(n510_adj_3802), .I2(n545), 
            .I3(n36910), .O(n15230[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_17 (.CI(n37958), .I0(n8317[14]), .I1(GND_net), .CO(n37959));
    SB_LUT4 mult_14_add_1216_19_lut (.I0(GND_net), .I1(n1802[16]), .I2(GND_net), 
            .I3(n38316), .O(n1801[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_16_lut (.I0(GND_net), .I1(n8317[13]), .I2(GND_net), 
            .I3(n37957), .O(n8298[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_2_lut (.I0(GND_net), .I1(n8_adj_3803), .I2(n101_adj_3804), 
            .I3(GND_net), .O(n7960[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_8 (.CI(n36910), .I0(n510_adj_3802), .I1(n545), .CO(n36911));
    SB_CARRY add_3084_2 (.CI(GND_net), .I0(n8_adj_3803), .I1(n101_adj_3804), 
            .CO(n37462));
    SB_LUT4 add_3407_7_lut (.I0(GND_net), .I1(n437_adj_3805), .I2(n472), 
            .I3(n36909), .O(n15230[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_7 (.CI(n36909), .I0(n437_adj_3805), .I1(n472), .CO(n36910));
    SB_CARRY mult_14_add_1216_19 (.CI(n38316), .I0(n1802[16]), .I1(GND_net), 
            .CO(n38317));
    SB_LUT4 add_3284_16_lut (.I0(GND_net), .I1(n13260[13]), .I2(GND_net), 
            .I3(n37461), .O(n12736[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_6_lut (.I0(GND_net), .I1(n364_adj_3806), .I2(n399), 
            .I3(n36908), .O(n15230[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_15_lut (.I0(GND_net), .I1(n13260[12]), .I2(GND_net), 
            .I3(n37460), .O(n12736[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_16 (.CI(n37957), .I0(n8317[13]), .I1(GND_net), .CO(n37958));
    SB_DFF pwm_count_1048__i2 (.Q(\pwm_count[2] ), .C(clk32MHz), .D(n75[2]));   // verilog/motorControl.v(99[18:29])
    SB_CARRY add_3407_6 (.CI(n36908), .I0(n364_adj_3806), .I1(n399), .CO(n36909));
    SB_CARRY add_3284_15 (.CI(n37460), .I0(n13260[12]), .I1(GND_net), 
            .CO(n37461));
    SB_LUT4 add_3407_5_lut (.I0(GND_net), .I1(n291), .I2(n326), .I3(n36907), 
            .O(n15230[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_14_lut (.I0(GND_net), .I1(n13260[11]), .I2(GND_net), 
            .I3(n37459), .O(n12736[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_5 (.CI(n36907), .I0(n291), .I1(n326), .CO(n36908));
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n61[6]), 
            .I3(n36570), .O(n58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_14 (.CI(n37459), .I0(n13260[11]), .I1(GND_net), 
            .CO(n37460));
    SB_LUT4 add_3407_4_lut (.I0(GND_net), .I1(n218_adj_3808), .I2(n253), 
            .I3(n36906), .O(n15230[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_8 (.CI(n36570), .I0(GND_net), .I1(n61[6]), 
            .CO(n36571));
    SB_LUT4 mult_14_add_1216_18_lut (.I0(GND_net), .I1(n1802[15]), .I2(GND_net), 
            .I3(n38315), .O(n1801[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_18 (.CI(n38315), .I0(n1802[15]), .I1(GND_net), 
            .CO(n38316));
    SB_CARRY add_3407_4 (.CI(n36906), .I0(n218_adj_3808), .I1(n253), .CO(n36907));
    SB_LUT4 add_3407_3_lut (.I0(GND_net), .I1(n145_adj_3809), .I2(n180_adj_3552), 
            .I3(n36905), .O(n15230[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_17_lut (.I0(GND_net), .I1(n1802[14]), .I2(GND_net), 
            .I3(n38314), .O(n1801[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_15_lut (.I0(GND_net), .I1(n8317[12]), .I2(GND_net), 
            .I3(n37956), .O(n8298[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_13_lut (.I0(GND_net), .I1(n13260[10]), .I2(GND_net), 
            .I3(n37458), .O(n12736[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_count_1048__i3 (.Q(\pwm_count[3] ), .C(clk32MHz), .D(n75[3]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1048__i4 (.Q(\pwm_count[4] ), .C(clk32MHz), .D(n75[4]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1048__i5 (.Q(\pwm_count[5] ), .C(clk32MHz), .D(n75[5]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1048__i6 (.Q(\pwm_count[6] ), .C(clk32MHz), .D(n75[6]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1048__i7 (.Q(\pwm_count[7] ), .C(clk32MHz), .D(n75[7]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1048__i8 (.Q(\pwm_count[8] ), .C(clk32MHz), .D(n75[8]));   // verilog/motorControl.v(99[18:29])
    SB_DFFE \PID_CONTROLLER.integral_1049__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[1]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1049__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[2]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1049__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[3]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1049__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[4]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1049__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[5]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1049__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[6]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1049__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[7]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1049__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[8]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1049__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(n55_adj_3661), .D(n82[9]));   // verilog/motorControl.v(34[21:33])
    SB_CARRY add_3284_13 (.CI(n37458), .I0(n13260[10]), .I1(GND_net), 
            .CO(n37459));
    SB_CARRY mult_14_add_1216_17 (.CI(n38314), .I0(n1802[14]), .I1(GND_net), 
            .CO(n38315));
    SB_LUT4 mult_14_add_1216_16_lut (.I0(GND_net), .I1(n1802[13]), .I2(GND_net), 
            .I3(n38313), .O(n1801[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_3 (.CI(n36905), .I0(n145_adj_3809), .I1(n180_adj_3552), 
            .CO(n36906));
    SB_CARRY add_3097_15 (.CI(n37956), .I0(n8317[12]), .I1(GND_net), .CO(n37957));
    SB_LUT4 add_3097_14_lut (.I0(GND_net), .I1(n8317[11]), .I2(GND_net), 
            .I3(n37955), .O(n8298[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_14 (.CI(n37955), .I0(n8317[11]), .I1(GND_net), .CO(n37956));
    SB_LUT4 add_3284_12_lut (.I0(GND_net), .I1(n13260[9]), .I2(GND_net), 
            .I3(n37457), .O(n12736[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_13_lut (.I0(GND_net), .I1(n8317[10]), .I2(GND_net), 
            .I3(n37954), .O(n8298[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_2_lut (.I0(GND_net), .I1(n72), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n15230[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_13 (.CI(n37954), .I0(n8317[10]), .I1(GND_net), .CO(n37955));
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n61[5]), 
            .I3(n36569), .O(n415)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_12 (.CI(n37457), .I0(n13260[9]), .I1(GND_net), .CO(n37458));
    SB_LUT4 add_3284_11_lut (.I0(GND_net), .I1(n13260[8]), .I2(GND_net), 
            .I3(n37456), .O(n12736[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_11 (.CI(n37456), .I0(n13260[8]), .I1(GND_net), .CO(n37457));
    SB_CARRY add_3407_2 (.CI(GND_net), .I0(n72), .I1(n107_adj_3557), .CO(n36905));
    SB_LUT4 add_3284_10_lut (.I0(GND_net), .I1(n13260[7]), .I2(GND_net), 
            .I3(n37455), .O(n12736[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_24_lut (.I0(GND_net), .I1(n13113[21]), .I2(GND_net), 
            .I3(n36904), .O(n12579[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_23_lut (.I0(GND_net), .I1(n13113[20]), .I2(GND_net), 
            .I3(n36903), .O(n12579[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i1  (.Q(\PID_CONTROLLER.err_prev[0] ), 
           .C(clk32MHz), .D(n23812));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3284_10 (.CI(n37455), .I0(n13260[7]), .I1(GND_net), .CO(n37456));
    SB_CARRY unary_minus_21_add_3_7 (.CI(n36569), .I0(GND_net), .I1(n61[5]), 
            .CO(n36570));
    SB_LUT4 add_3284_9_lut (.I0(GND_net), .I1(n13260[6]), .I2(GND_net), 
            .I3(n37454), .O(n12736[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n61[4]), 
            .I3(n36568), .O(n416)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_23 (.CI(n36903), .I0(n13113[20]), .I1(GND_net), 
            .CO(n36904));
    SB_CARRY unary_minus_21_add_3_6 (.CI(n36568), .I0(GND_net), .I1(n61[4]), 
            .CO(n36569));
    SB_LUT4 add_3276_22_lut (.I0(GND_net), .I1(n13113[19]), .I2(GND_net), 
            .I3(n36902), .O(n12579[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_9 (.CI(n37454), .I0(n13260[6]), .I1(GND_net), .CO(n37455));
    SB_LUT4 add_3097_12_lut (.I0(GND_net), .I1(n8317[9]), .I2(GND_net), 
            .I3(n37953), .O(n8298[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_22 (.CI(n36902), .I0(n13113[19]), .I1(GND_net), 
            .CO(n36903));
    SB_CARRY mult_14_add_1216_16 (.CI(n38313), .I0(n1802[13]), .I1(GND_net), 
            .CO(n38314));
    SB_CARRY add_3097_12 (.CI(n37953), .I0(n8317[9]), .I1(GND_net), .CO(n37954));
    SB_LUT4 add_3284_8_lut (.I0(GND_net), .I1(n13260[5]), .I2(n545), .I3(n37453), 
            .O(n12736[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_21_lut (.I0(GND_net), .I1(n13113[18]), .I2(GND_net), 
            .I3(n36901), .O(n12579[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_8 (.CI(n37453), .I0(n13260[5]), .I1(n545), .CO(n37454));
    SB_LUT4 mult_14_add_1216_15_lut (.I0(GND_net), .I1(n1802[12]), .I2(GND_net), 
            .I3(n38312), .O(n1801[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_7_lut (.I0(GND_net), .I1(n13260[4]), .I2(n472), .I3(n37452), 
            .O(n12736[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_21 (.CI(n36901), .I0(n13113[18]), .I1(GND_net), 
            .CO(n36902));
    SB_LUT4 add_3276_20_lut (.I0(GND_net), .I1(n13113[17]), .I2(GND_net), 
            .I3(n36900), .O(n12579[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_11_lut (.I0(GND_net), .I1(n8317[8]), .I2(GND_net), 
            .I3(n37952), .O(n8298[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_15 (.CI(n38312), .I0(n1802[12]), .I1(GND_net), 
            .CO(n38313));
    SB_CARRY add_3097_11 (.CI(n37952), .I0(n8317[8]), .I1(GND_net), .CO(n37953));
    SB_LUT4 add_3097_10_lut (.I0(GND_net), .I1(n8317[7]), .I2(GND_net), 
            .I3(n37951), .O(n8298[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_14_lut (.I0(GND_net), .I1(n1802[11]), .I2(GND_net), 
            .I3(n38311), .O(n1801[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_10 (.CI(n37951), .I0(n8317[7]), .I1(GND_net), .CO(n37952));
    SB_LUT4 add_3097_9_lut (.I0(GND_net), .I1(n8317[6]), .I2(GND_net), 
            .I3(n37950), .O(n8298[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_14 (.CI(n38311), .I0(n1802[11]), .I1(GND_net), 
            .CO(n38312));
    SB_LUT4 mult_14_add_1216_13_lut (.I0(GND_net), .I1(n1802[10]), .I2(GND_net), 
            .I3(n38310), .O(n1801[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_13 (.CI(n38310), .I0(n1802[10]), .I1(GND_net), 
            .CO(n38311));
    SB_LUT4 mult_14_add_1216_12_lut (.I0(GND_net), .I1(n1802[9]), .I2(GND_net), 
            .I3(n38309), .O(n1801[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_12 (.CI(n38309), .I0(n1802[9]), .I1(GND_net), 
            .CO(n38310));
    SB_CARRY add_3284_7 (.CI(n37452), .I0(n13260[4]), .I1(n472), .CO(n37453));
    SB_CARRY add_3097_9 (.CI(n37950), .I0(n8317[6]), .I1(GND_net), .CO(n37951));
    SB_LUT4 add_3284_6_lut (.I0(GND_net), .I1(n13260[3]), .I2(n399), .I3(n37451), 
            .O(n12736[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_8_lut (.I0(GND_net), .I1(n8317[5]), .I2(n722_adj_3813), 
            .I3(n37949), .O(n8298[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_11_lut (.I0(GND_net), .I1(n1802[8]), .I2(GND_net), 
            .I3(n38308), .O(n1801[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_6 (.CI(n37451), .I0(n13260[3]), .I1(n399), .CO(n37452));
    SB_CARRY add_3097_8 (.CI(n37949), .I0(n8317[5]), .I1(n722_adj_3813), 
            .CO(n37950));
    SB_LUT4 add_3284_5_lut (.I0(GND_net), .I1(n13260[2]), .I2(n326), .I3(n37450), 
            .O(n12736[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_7_lut (.I0(GND_net), .I1(n8317[4]), .I2(n625_adj_3814), 
            .I3(n37948), .O(n8298[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_11 (.CI(n38308), .I0(n1802[8]), .I1(GND_net), 
            .CO(n38309));
    SB_CARRY add_3284_5 (.CI(n37450), .I0(n13260[2]), .I1(n326), .CO(n37451));
    SB_CARRY add_3097_7 (.CI(n37948), .I0(n8317[4]), .I1(n625_adj_3814), 
            .CO(n37949));
    SB_LUT4 add_3284_4_lut (.I0(GND_net), .I1(n13260[1]), .I2(n253), .I3(n37449), 
            .O(n12736[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_6_lut (.I0(GND_net), .I1(n8317[3]), .I2(n528_adj_3815), 
            .I3(n37947), .O(n8298[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_10_lut (.I0(GND_net), .I1(n1802[7]), .I2(GND_net), 
            .I3(n38307), .O(n1801[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_4 (.CI(n37449), .I0(n13260[1]), .I1(n253), .CO(n37450));
    SB_CARRY add_3097_6 (.CI(n37947), .I0(n8317[3]), .I1(n528_adj_3815), 
            .CO(n37948));
    SB_LUT4 add_3284_3_lut (.I0(GND_net), .I1(n13260[0]), .I2(n180_adj_3552), 
            .I3(n37448), .O(n12736[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_5_lut (.I0(GND_net), .I1(n8317[2]), .I2(n431_adj_3816), 
            .I3(n37946), .O(n8298[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_10 (.CI(n38307), .I0(n1802[7]), .I1(GND_net), 
            .CO(n38308));
    SB_CARRY add_3097_5 (.CI(n37946), .I0(n8317[2]), .I1(n431_adj_3816), 
            .CO(n37947));
    SB_LUT4 add_3097_4_lut (.I0(GND_net), .I1(n8317[1]), .I2(n334_adj_3817), 
            .I3(n37945), .O(n8298[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_9_lut (.I0(GND_net), .I1(n1802[6]), .I2(GND_net), 
            .I3(n38306), .O(n1801[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_4 (.CI(n37945), .I0(n8317[1]), .I1(n334_adj_3817), 
            .CO(n37946));
    SB_LUT4 add_3097_3_lut (.I0(GND_net), .I1(n8317[0]), .I2(n237_adj_3818), 
            .I3(n37944), .O(n8298[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_9 (.CI(n38306), .I0(n1802[6]), .I1(GND_net), 
            .CO(n38307));
    SB_CARRY add_3097_3 (.CI(n37944), .I0(n8317[0]), .I1(n237_adj_3818), 
            .CO(n37945));
    SB_LUT4 add_3097_2_lut (.I0(GND_net), .I1(n47_adj_3819), .I2(n140_adj_3820), 
            .I3(GND_net), .O(n8298[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_8_lut (.I0(GND_net), .I1(n1802[5]), .I2(n527), 
            .I3(n38305), .O(n1801[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_2 (.CI(GND_net), .I0(n47_adj_3819), .I1(n140_adj_3820), 
            .CO(n37944));
    SB_LUT4 add_3096_19_lut (.I0(GND_net), .I1(n8298[16]), .I2(GND_net), 
            .I3(n37943), .O(n8278[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_8 (.CI(n38305), .I0(n1802[5]), .I1(n527), 
            .CO(n38306));
    SB_CARRY add_3284_3 (.CI(n37448), .I0(n13260[0]), .I1(n180_adj_3552), 
            .CO(n37449));
    SB_LUT4 add_3096_18_lut (.I0(GND_net), .I1(n8298[15]), .I2(GND_net), 
            .I3(n37942), .O(n8278[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_2_lut (.I0(GND_net), .I1(n35_adj_3556), .I2(n107_adj_3557), 
            .I3(GND_net), .O(n12736[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_18 (.CI(n37942), .I0(n8298[15]), .I1(GND_net), .CO(n37943));
    SB_LUT4 mult_14_add_1216_7_lut (.I0(GND_net), .I1(n1802[4]), .I2(n454), 
            .I3(n38304), .O(n1801[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_2 (.CI(GND_net), .I0(n35_adj_3556), .I1(n107_adj_3557), 
            .CO(n37448));
    SB_LUT4 add_3096_17_lut (.I0(GND_net), .I1(n8298[14]), .I2(GND_net), 
            .I3(n37941), .O(n8278[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1047_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[6]), .I3(n37447), .O(n57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1047_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_17 (.CI(n37941), .I0(n8298[14]), .I1(GND_net), .CO(n37942));
    SB_CARRY mult_14_add_1216_7 (.CI(n38304), .I0(n1802[4]), .I1(n454), 
            .CO(n38305));
    SB_LUT4 Kd_delay_counter_1047_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[5]), .I3(n37446), .O(n57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1047_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_16_lut (.I0(GND_net), .I1(n8298[13]), .I2(GND_net), 
            .I3(n37940), .O(n8278[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1047_add_4_7 (.CI(n37446), .I0(GND_net), .I1(Kd_delay_counter[5]), 
            .CO(n37447));
    SB_CARRY add_3096_16 (.CI(n37940), .I0(n8298[13]), .I1(GND_net), .CO(n37941));
    SB_LUT4 mult_14_add_1216_6_lut (.I0(GND_net), .I1(n1802[3]), .I2(n381), 
            .I3(n38303), .O(n1801[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1047_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[4]), .I3(n37445), .O(n57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1047_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_15_lut (.I0(GND_net), .I1(n8298[12]), .I2(GND_net), 
            .I3(n37939), .O(n8278[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_15 (.CI(n37939), .I0(n8298[12]), .I1(GND_net), .CO(n37940));
    SB_CARRY mult_14_add_1216_6 (.CI(n38303), .I0(n1802[3]), .I1(n381), 
            .CO(n38304));
    SB_LUT4 add_3096_14_lut (.I0(GND_net), .I1(n8298[11]), .I2(GND_net), 
            .I3(n37938), .O(n8278[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_14 (.CI(n37938), .I0(n8298[11]), .I1(GND_net), .CO(n37939));
    SB_LUT4 mult_14_add_1216_5_lut (.I0(GND_net), .I1(n1802[2]), .I2(n308_adj_3821), 
            .I3(n38302), .O(n1801[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_13_lut (.I0(GND_net), .I1(n8298[10]), .I2(GND_net), 
            .I3(n37937), .O(n8278[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_13 (.CI(n37937), .I0(n8298[10]), .I1(GND_net), .CO(n37938));
    SB_CARRY mult_14_add_1216_5 (.CI(n38302), .I0(n1802[2]), .I1(n308_adj_3821), 
            .CO(n38303));
    SB_LUT4 add_3096_12_lut (.I0(GND_net), .I1(n8298[9]), .I2(GND_net), 
            .I3(n37936), .O(n8278[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_12 (.CI(n37936), .I0(n8298[9]), .I1(GND_net), .CO(n37937));
    SB_LUT4 mult_14_add_1216_4_lut (.I0(GND_net), .I1(n1802[1]), .I2(n235_adj_3822), 
            .I3(n38301), .O(n1801[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_11_lut (.I0(GND_net), .I1(n8298[8]), .I2(GND_net), 
            .I3(n37935), .O(n8278[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_4 (.CI(n38301), .I0(n1802[1]), .I1(n235_adj_3822), 
            .CO(n38302));
    SB_LUT4 mult_14_add_1216_3_lut (.I0(GND_net), .I1(n1802[0]), .I2(n162), 
            .I3(n38300), .O(n1801[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_3 (.CI(n38300), .I0(n1802[0]), .I1(n162), 
            .CO(n38301));
    SB_LUT4 mult_14_add_1216_2_lut (.I0(GND_net), .I1(n20_adj_3823), .I2(n89), 
            .I3(GND_net), .O(n1801[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_2 (.CI(GND_net), .I0(n20_adj_3823), .I1(n89), 
            .CO(n38300));
    SB_LUT4 mult_14_add_1215_24_lut (.I0(GND_net), .I1(n1801[21]), .I2(GND_net), 
            .I3(n38298), .O(n1800[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_24 (.CI(n38298), .I0(n1801[21]), .I1(GND_net), 
            .CO(n1699));
    SB_LUT4 mult_14_add_1215_23_lut (.I0(GND_net), .I1(n1801[20]), .I2(GND_net), 
            .I3(n38297), .O(n1800[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_23 (.CI(n38297), .I0(n1801[20]), .I1(GND_net), 
            .CO(n38298));
    SB_CARRY add_3096_11 (.CI(n37935), .I0(n8298[8]), .I1(GND_net), .CO(n37936));
    SB_LUT4 add_3096_10_lut (.I0(GND_net), .I1(n8298[7]), .I2(GND_net), 
            .I3(n37934), .O(n8278[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_22_lut (.I0(GND_net), .I1(n1801[19]), .I2(GND_net), 
            .I3(n38296), .O(n1800[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_10 (.CI(n37934), .I0(n8298[7]), .I1(GND_net), .CO(n37935));
    SB_LUT4 add_3096_9_lut (.I0(GND_net), .I1(n8298[6]), .I2(GND_net), 
            .I3(n37933), .O(n8278[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_22 (.CI(n38296), .I0(n1801[19]), .I1(GND_net), 
            .CO(n38297));
    SB_CARRY add_3096_9 (.CI(n37933), .I0(n8298[6]), .I1(GND_net), .CO(n37934));
    SB_LUT4 add_3096_8_lut (.I0(GND_net), .I1(n8298[5]), .I2(n719_adj_3824), 
            .I3(n37932), .O(n8278[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_21_lut (.I0(GND_net), .I1(n1801[18]), .I2(GND_net), 
            .I3(n38295), .O(n1800[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_8 (.CI(n37932), .I0(n8298[5]), .I1(n719_adj_3824), 
            .CO(n37933));
    SB_LUT4 add_3096_7_lut (.I0(GND_net), .I1(n8298[4]), .I2(n622_adj_3825), 
            .I3(n37931), .O(n8278[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_21 (.CI(n38295), .I0(n1801[18]), .I1(GND_net), 
            .CO(n38296));
    SB_CARRY add_3096_7 (.CI(n37931), .I0(n8298[4]), .I1(n622_adj_3825), 
            .CO(n37932));
    SB_LUT4 add_3096_6_lut (.I0(GND_net), .I1(n8298[3]), .I2(n525_adj_3826), 
            .I3(n37930), .O(n8278[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_20_lut (.I0(GND_net), .I1(n1801[17]), .I2(GND_net), 
            .I3(n38294), .O(n1800[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_6 (.CI(n37930), .I0(n8298[3]), .I1(n525_adj_3826), 
            .CO(n37931));
    SB_LUT4 add_3096_5_lut (.I0(GND_net), .I1(n8298[2]), .I2(n428_adj_3827), 
            .I3(n37929), .O(n8278[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_20 (.CI(n38294), .I0(n1801[17]), .I1(GND_net), 
            .CO(n38295));
    SB_CARRY add_3096_5 (.CI(n37929), .I0(n8298[2]), .I1(n428_adj_3827), 
            .CO(n37930));
    SB_LUT4 add_3096_4_lut (.I0(GND_net), .I1(n8298[1]), .I2(n331_adj_3828), 
            .I3(n37928), .O(n8278[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_19_lut (.I0(GND_net), .I1(n1801[16]), .I2(GND_net), 
            .I3(n38293), .O(n1800[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_4 (.CI(n37928), .I0(n8298[1]), .I1(n331_adj_3828), 
            .CO(n37929));
    SB_LUT4 add_3096_3_lut (.I0(GND_net), .I1(n8298[0]), .I2(n234_adj_3829), 
            .I3(n37927), .O(n8278[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_19 (.CI(n38293), .I0(n1801[16]), .I1(GND_net), 
            .CO(n38294));
    SB_CARRY add_3096_3 (.CI(n37927), .I0(n8298[0]), .I1(n234_adj_3829), 
            .CO(n37928));
    SB_LUT4 add_3096_2_lut (.I0(GND_net), .I1(n44_adj_3830), .I2(n137_adj_3831), 
            .I3(GND_net), .O(n8278[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_18_lut (.I0(GND_net), .I1(n1801[15]), .I2(GND_net), 
            .I3(n38292), .O(n1800[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_2 (.CI(GND_net), .I0(n44_adj_3830), .I1(n137_adj_3831), 
            .CO(n37927));
    SB_LUT4 add_3095_20_lut (.I0(GND_net), .I1(n8278[17]), .I2(GND_net), 
            .I3(n37926), .O(n8257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_18 (.CI(n38292), .I0(n1801[15]), .I1(GND_net), 
            .CO(n38293));
    SB_LUT4 add_3095_19_lut (.I0(GND_net), .I1(n8278[16]), .I2(GND_net), 
            .I3(n37925), .O(n8257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_19 (.CI(n37925), .I0(n8278[16]), .I1(GND_net), .CO(n37926));
    SB_LUT4 mult_14_add_1215_17_lut (.I0(GND_net), .I1(n1801[14]), .I2(GND_net), 
            .I3(n38291), .O(n1800[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_18_lut (.I0(GND_net), .I1(n8278[15]), .I2(GND_net), 
            .I3(n37924), .O(n8257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_18 (.CI(n37924), .I0(n8278[15]), .I1(GND_net), .CO(n37925));
    SB_CARRY mult_14_add_1215_17 (.CI(n38291), .I0(n1801[14]), .I1(GND_net), 
            .CO(n38292));
    SB_LUT4 add_3095_17_lut (.I0(GND_net), .I1(n8278[14]), .I2(GND_net), 
            .I3(n37923), .O(n8257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_17 (.CI(n37923), .I0(n8278[14]), .I1(GND_net), .CO(n37924));
    SB_LUT4 mult_14_add_1215_16_lut (.I0(GND_net), .I1(n1801[13]), .I2(GND_net), 
            .I3(n38290), .O(n1800[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_16_lut (.I0(GND_net), .I1(n8278[13]), .I2(GND_net), 
            .I3(n37922), .O(n8257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_16 (.CI(n37922), .I0(n8278[13]), .I1(GND_net), .CO(n37923));
    SB_CARRY mult_14_add_1215_16 (.CI(n38290), .I0(n1801[13]), .I1(GND_net), 
            .CO(n38291));
    SB_LUT4 add_3095_15_lut (.I0(GND_net), .I1(n8278[12]), .I2(GND_net), 
            .I3(n37921), .O(n8257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_15 (.CI(n37921), .I0(n8278[12]), .I1(GND_net), .CO(n37922));
    SB_LUT4 mult_14_add_1215_15_lut (.I0(GND_net), .I1(n1801[12]), .I2(GND_net), 
            .I3(n38289), .O(n1800[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_14_lut (.I0(GND_net), .I1(n8278[11]), .I2(GND_net), 
            .I3(n37920), .O(n8257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_14 (.CI(n37920), .I0(n8278[11]), .I1(GND_net), .CO(n37921));
    SB_CARRY mult_14_add_1215_15 (.CI(n38289), .I0(n1801[12]), .I1(GND_net), 
            .CO(n38290));
    SB_LUT4 add_3095_13_lut (.I0(GND_net), .I1(n8278[10]), .I2(GND_net), 
            .I3(n37919), .O(n8257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_13 (.CI(n37919), .I0(n8278[10]), .I1(GND_net), .CO(n37920));
    SB_LUT4 mult_14_add_1215_14_lut (.I0(GND_net), .I1(n1801[11]), .I2(GND_net), 
            .I3(n38288), .O(n1800[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_12_lut (.I0(GND_net), .I1(n8278[9]), .I2(GND_net), 
            .I3(n37918), .O(n8257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_12 (.CI(n37918), .I0(n8278[9]), .I1(GND_net), .CO(n37919));
    SB_CARRY mult_14_add_1215_14 (.CI(n38288), .I0(n1801[11]), .I1(GND_net), 
            .CO(n38289));
    SB_LUT4 add_3095_11_lut (.I0(GND_net), .I1(n8278[8]), .I2(GND_net), 
            .I3(n37917), .O(n8257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_11 (.CI(n37917), .I0(n8278[8]), .I1(GND_net), .CO(n37918));
    SB_LUT4 mult_14_add_1215_13_lut (.I0(GND_net), .I1(n1801[10]), .I2(GND_net), 
            .I3(n38287), .O(n1800[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_10_lut (.I0(GND_net), .I1(n8278[7]), .I2(GND_net), 
            .I3(n37916), .O(n8257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_10 (.CI(n37916), .I0(n8278[7]), .I1(GND_net), .CO(n37917));
    SB_CARRY mult_14_add_1215_13 (.CI(n38287), .I0(n1801[10]), .I1(GND_net), 
            .CO(n38288));
    SB_LUT4 add_3095_9_lut (.I0(GND_net), .I1(n8278[6]), .I2(GND_net), 
            .I3(n37915), .O(n8257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_9 (.CI(n37915), .I0(n8278[6]), .I1(GND_net), .CO(n37916));
    SB_LUT4 mult_14_add_1215_12_lut (.I0(GND_net), .I1(n1801[9]), .I2(GND_net), 
            .I3(n38286), .O(n1800[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_8_lut (.I0(GND_net), .I1(n8278[5]), .I2(n716_adj_3832), 
            .I3(n37914), .O(n8257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_8 (.CI(n37914), .I0(n8278[5]), .I1(n716_adj_3832), 
            .CO(n37915));
    SB_CARRY mult_14_add_1215_12 (.CI(n38286), .I0(n1801[9]), .I1(GND_net), 
            .CO(n38287));
    SB_LUT4 add_3095_7_lut (.I0(GND_net), .I1(n8278[4]), .I2(n619_adj_3833), 
            .I3(n37913), .O(n8257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_7 (.CI(n37913), .I0(n8278[4]), .I1(n619_adj_3833), 
            .CO(n37914));
    SB_LUT4 mult_14_add_1215_11_lut (.I0(GND_net), .I1(n1801[8]), .I2(GND_net), 
            .I3(n38285), .O(n1800[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_6_lut (.I0(GND_net), .I1(n8278[3]), .I2(n522_adj_3834), 
            .I3(n37912), .O(n8257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_6 (.CI(n37912), .I0(n8278[3]), .I1(n522_adj_3834), 
            .CO(n37913));
    SB_CARRY mult_14_add_1215_11 (.CI(n38285), .I0(n1801[8]), .I1(GND_net), 
            .CO(n38286));
    SB_LUT4 mux_24_i2_3_lut (.I0(\PID_CONTROLLER.result [1]), .I1(n58[1]), 
            .I2(n421), .I3(GND_net), .O(n470));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i3_3_lut (.I0(\PID_CONTROLLER.result [2]), .I1(n58[2]), 
            .I2(n421), .I3(GND_net), .O(n469));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i4_3_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n58[3]), 
            .I2(n421), .I3(GND_net), .O(n468));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(pwm_23__N_2948), .I1(n28170), .I2(\PWMLimit[4] ), 
            .I3(n387), .O(n24432));   // verilog/motorControl.v(37[10:51])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1385 (.I0(pwm_23__N_2948), .I1(n28227), .I2(\PWMLimit[5] ), 
            .I3(n387), .O(n24433));   // verilog/motorControl.v(37[10:51])
    defparam i1_4_lut_adj_1385.LUT_INIT = 16'ha088;
    SB_LUT4 mux_24_i7_3_lut (.I0(\PID_CONTROLLER.result [6]), .I1(n58[6]), 
            .I2(n421), .I3(GND_net), .O(n465));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1386 (.I0(pwm_23__N_2948), .I1(n1), .I2(\PWMLimit[7] ), 
            .I3(n387), .O(n24435));   // verilog/motorControl.v(37[10:51])
    defparam i1_4_lut_adj_1386.LUT_INIT = 16'ha088;
    SB_LUT4 mux_24_i9_3_lut (.I0(\PID_CONTROLLER.result [8]), .I1(n58[8]), 
            .I2(n421), .I3(GND_net), .O(n463));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i10_3_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n58[9]), 
            .I2(n421), .I3(GND_net), .O(n462));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i11_3_lut (.I0(\PID_CONTROLLER.result [10]), .I1(n58[10]), 
            .I2(n421), .I3(GND_net), .O(n461));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i12_3_lut (.I0(\PID_CONTROLLER.result [11]), .I1(n58[10]), 
            .I2(n421), .I3(GND_net), .O(n460));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i13_3_lut (.I0(\PID_CONTROLLER.result [12]), .I1(n58[10]), 
            .I2(n421), .I3(GND_net), .O(n459));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i14_3_lut (.I0(\PID_CONTROLLER.result [13]), .I1(n58[10]), 
            .I2(n421), .I3(GND_net), .O(n458));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i15_3_lut (.I0(\PID_CONTROLLER.result [14]), .I1(n58[10]), 
            .I2(n421), .I3(GND_net), .O(n457));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i16_3_lut (.I0(\PID_CONTROLLER.result [15]), .I1(n58[10]), 
            .I2(n421), .I3(GND_net), .O(n456));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i17_3_lut (.I0(\PID_CONTROLLER.result [16]), .I1(n58[10]), 
            .I2(n421), .I3(GND_net), .O(n455));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1387 (.I0(pwm_23__N_2948), .I1(n46606), .I2(\PWMLimit[9] ), 
            .I3(n387), .O(n41482));
    defparam i1_4_lut_adj_1387.LUT_INIT = 16'ha088;
    SB_LUT4 pwm_23__I_816_i13_2_lut (.I0(\PID_CONTROLLER.result [6]), .I1(pwm_23__N_2951[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_3842));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i7_2_lut  (.I0(\deadband[3] ), 
            .I1(\PID_CONTROLLER.result [3]), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_3843));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i7_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i11_2_lut  (.I0(\deadband[5] ), 
            .I1(\PID_CONTROLLER.result[5] ), .I2(GND_net), .I3(GND_net), 
            .O(n11_adj_3844));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i11_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i13_2_lut  (.I0(\deadband[6] ), 
            .I1(\PID_CONTROLLER.result [6]), .I2(GND_net), .I3(GND_net), 
            .O(n13_adj_3845));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i13_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i17_2_lut  (.I0(\deadband[8] ), 
            .I1(\PID_CONTROLLER.result [8]), .I2(GND_net), .I3(GND_net), 
            .O(n17_adj_3846));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i17_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 i32211_4_lut (.I0(\deadband[9] ), .I1(n17_adj_3846), .I2(\PID_CONTROLLER.result [9]), 
            .I3(n9), .O(n47725));
    defparam i32211_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32205_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [11]), .I3(n47725), .O(n47719));
    defparam i32205_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i32219_3_lut (.I0(n15), .I1(n13_adj_3845), .I2(n11_adj_3844), 
            .I3(GND_net), .O(n47733));
    defparam i32219_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i32191_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [13]), 
            .I2(\PID_CONTROLLER.result [14]), .I3(n47733), .O(n47705));
    defparam i32191_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i32171_4_lut (.I0(\PID_CONTROLLER.result [17]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(\deadband[9] ), .I3(n15), .O(n47685));
    defparam i32171_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i30_4_lut  (.I0(\PID_CONTROLLER.result[7] ), 
            .I1(\PID_CONTROLLER.result [17]), .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [16]), 
            .O(n30_adj_3849));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i30_4_lut .LUT_INIT = 16'h8f0e;
    SB_LUT4 i32229_4_lut (.I0(n9), .I1(n7_adj_3843), .I2(\deadband[2] ), 
            .I3(\PID_CONTROLLER.result [2]), .O(n47743));
    defparam i32229_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i32523_4_lut (.I0(n15), .I1(n13_adj_3845), .I2(n11_adj_3844), 
            .I3(n47743), .O(n48037));
    defparam i32523_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32215_4_lut (.I0(\deadband[9] ), .I1(n17_adj_3846), .I2(\PID_CONTROLLER.result [9]), 
            .I3(n48037), .O(n47729));
    defparam i32215_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i32769_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [11]), .I3(n47729), .O(n48283));
    defparam i32769_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i31591_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [12]), 
            .I2(\PID_CONTROLLER.result [13]), .I3(n48283), .O(n47105));
    defparam i31591_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 mult_14_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32507_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(n47105), .O(n48021));
    defparam i32507_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i32923_4_lut (.I0(\PID_CONTROLLER.result [17]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(\deadband[9] ), .I3(n48021), .O(n48437));
    defparam i32923_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 mult_14_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33070_4_lut (.I0(\PID_CONTROLLER.result [19]), .I1(\PID_CONTROLLER.result [18]), 
            .I2(\deadband[9] ), .I3(n48437), .O(n48584));
    defparam i33070_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i32655_3_lut (.I0(n6_adj_3850), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n48169));   // verilog/motorControl.v(37[10:27])
    defparam i32655_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32147_4_lut (.I0(\PID_CONTROLLER.result [22]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [9]), .O(n47661));
    defparam i32147_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i24_4_lut  (.I0(\PID_CONTROLLER.result [9]), 
            .I1(\PID_CONTROLLER.result [22]), .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [21]), 
            .O(n24_adj_3851));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i24_4_lut .LUT_INIT = 16'h8f0e;
    SB_LUT4 i31549_4_lut (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [12]), 
            .I2(\deadband[9] ), .I3(n47719), .O(n47063));
    defparam i31549_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i17_rep_164_2_lut (.I0(\PID_CONTROLLER.result [22]), .I1(\deadband[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n49657));   // verilog/TinyFPGA_B.v(85[22:30])
    defparam i17_rep_164_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32871_3_lut (.I0(n24_adj_3851), .I1(n8_adj_3852), .I2(n47661), 
            .I3(GND_net), .O(n48385));   // verilog/motorControl.v(37[10:27])
    defparam i32871_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31952_4_lut (.I0(n48169), .I1(\PID_CONTROLLER.result [12]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [11]), .O(n47466));   // verilog/motorControl.v(37[10:27])
    defparam i31952_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i4_4_lut  (.I0(\deadband[0] ), 
            .I1(\PID_CONTROLLER.result [1]), .I2(\deadband[1] ), .I3(\PID_CONTROLLER.result [0]), 
            .O(n4_adj_3853));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i4_4_lut .LUT_INIT = 16'h4d0c;
    SB_LUT4 i32653_3_lut (.I0(n4_adj_3853), .I1(\PID_CONTROLLER.result [13]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n48167));   // verilog/motorControl.v(37[10:27])
    defparam i32653_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31579_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [15]), 
            .I2(\PID_CONTROLLER.result [16]), .I3(n47705), .O(n47093));
    defparam i31579_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i19_rep_142_2_lut (.I0(\PID_CONTROLLER.result [17]), .I1(\deadband[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n49635));   // verilog/TinyFPGA_B.v(85[22:30])
    defparam i19_rep_142_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32989_3_lut (.I0(n30_adj_3849), .I1(n10_adj_3854), .I2(n47685), 
            .I3(GND_net), .O(n48503));   // verilog/motorControl.v(37[10:27])
    defparam i32989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31954_4_lut (.I0(n48167), .I1(\PID_CONTROLLER.result [15]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [14]), .O(n47468));   // verilog/motorControl.v(37[10:27])
    defparam i31954_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i33090_4_lut (.I0(n47468), .I1(n48503), .I2(n49635), .I3(n47093), 
            .O(n48604));   // verilog/motorControl.v(37[10:27])
    defparam i33090_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33091_3_lut (.I0(n48604), .I1(\PID_CONTROLLER.result [18]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n48605));   // verilog/motorControl.v(37[10:27])
    defparam i33091_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31553_4_lut (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [20]), 
            .I2(\deadband[9] ), .I3(n48584), .O(n47067));
    defparam i31553_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i33020_4_lut (.I0(n47466), .I1(n48385), .I2(n49657), .I3(n47063), 
            .O(n48534));   // verilog/motorControl.v(37[10:27])
    defparam i33020_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31960_4_lut (.I0(n48605), .I1(\PID_CONTROLLER.result [20]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [19]), .O(n47474));   // verilog/motorControl.v(37[10:27])
    defparam i31960_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i33086_4_lut (.I0(n47474), .I1(n48534), .I2(n49657), .I3(n47067), 
            .O(n48600));   // verilog/motorControl.v(37[10:27])
    defparam i33086_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33054_4_lut (.I0(n48600), .I1(\PID_CONTROLLER.result [24]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [23]), .O(n50_adj_3855));   // verilog/motorControl.v(37[10:27])
    defparam i33054_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 mult_12_i349_2_lut (.I0(\Kd[5] ), .I1(n67[11]), .I2(GND_net), 
            .I3(GND_net), .O(n519));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_816_i19_2_lut (.I0(\PID_CONTROLLER.result [9]), .I1(pwm_23__N_2951[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3856));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_23__I_816_i17_2_lut (.I0(\PID_CONTROLLER.result [8]), .I1(pwm_23__N_2951[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3857));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_23__I_816_i7_2_lut (.I0(\PID_CONTROLLER.result [3]), .I1(pwm_23__N_2951[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3858));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i13_2_lut (.I0(\PWMLimit[6] ), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_3859));   // verilog/motorControl.v(38[12:27])
    defparam LessThan_20_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32645_3_lut (.I0(n4_adj_3860), .I1(\PID_CONTROLLER.result[5] ), 
            .I2(n11), .I3(GND_net), .O(n48159));   // verilog/motorControl.v(38[12:27])
    defparam i32645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32646_3_lut (.I0(n48159), .I1(\PID_CONTROLLER.result [6]), 
            .I2(n13_adj_3859), .I3(GND_net), .O(n48160));   // verilog/motorControl.v(38[12:27])
    defparam i32646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32109_4_lut (.I0(n13_adj_3859), .I1(n11), .I2(n9_adj_10), 
            .I3(n46986), .O(n47623));
    defparam i32109_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_20_i8_3_lut (.I0(n6_adj_3863), .I1(\PID_CONTROLLER.result[4] ), 
            .I2(n9_adj_10), .I3(GND_net), .O(n8_adj_3864));   // verilog/motorControl.v(38[12:27])
    defparam LessThan_20_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31964_3_lut (.I0(n48160), .I1(\PID_CONTROLLER.result[7] ), 
            .I2(n15_adj_11), .I3(GND_net), .O(n47478));   // verilog/motorControl.v(38[12:27])
    defparam i31964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32673_4_lut (.I0(n47478), .I1(n8_adj_3864), .I2(n15_adj_11), 
            .I3(n47623), .O(n48187));   // verilog/motorControl.v(38[12:27])
    defparam i32673_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32674_3_lut (.I0(n48187), .I1(\PID_CONTROLLER.result [8]), 
            .I2(\PWMLimit[8] ), .I3(GND_net), .O(n18_adj_3866));   // verilog/motorControl.v(38[12:27])
    defparam i32674_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i3_4_lut (.I0(\PID_CONTROLLER.result [11]), .I1(n18_adj_3866), 
            .I2(\PID_CONTROLLER.result [9]), .I3(\PID_CONTROLLER.result [10]), 
            .O(n44105));   // verilog/motorControl.v(38[12:27])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n18_adj_3866), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [9]), .I3(\PID_CONTROLLER.result [11]), 
            .O(n43893));   // verilog/motorControl.v(38[12:27])
    defparam i2_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1388 (.I0(\PID_CONTROLLER.result [12]), .I1(\PWMLimit[9] ), 
            .I2(n43893), .I3(n44105), .O(n26_adj_3867));   // verilog/motorControl.v(38[12:27])
    defparam i1_4_lut_adj_1388.LUT_INIT = 16'hb3a2;
    SB_LUT4 i3_4_lut_adj_1389 (.I0(\PID_CONTROLLER.result [15]), .I1(n26_adj_3867), 
            .I2(\PID_CONTROLLER.result [13]), .I3(\PID_CONTROLLER.result [14]), 
            .O(n44113));   // verilog/motorControl.v(38[12:27])
    defparam i3_4_lut_adj_1389.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1390 (.I0(n26_adj_3867), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [13]), .I3(\PID_CONTROLLER.result [15]), 
            .O(n43892));   // verilog/motorControl.v(38[12:27])
    defparam i2_4_lut_adj_1390.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1391 (.I0(\PID_CONTROLLER.result [16]), .I1(\PWMLimit[9] ), 
            .I2(n43892), .I3(n44113), .O(n34_adj_3868));   // verilog/motorControl.v(38[12:27])
    defparam i1_4_lut_adj_1391.LUT_INIT = 16'hb3a2;
    SB_LUT4 i1_4_lut_adj_1392 (.I0(\PID_CONTROLLER.result [26]), .I1(n62_adj_3869), 
            .I2(n49_adj_3870), .I3(n34_adj_3868), .O(n42736));   // verilog/motorControl.v(38[12:27])
    defparam i1_4_lut_adj_1392.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(n42695), .I1(\PID_CONTROLLER.result [26]), .I2(n34_adj_3868), 
            .I3(GND_net), .O(n44333));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_adj_1393 (.I0(\PID_CONTROLLER.result [27]), .I1(\PWMLimit[9] ), 
            .I2(n44333), .I3(n42736), .O(n56_adj_3871));   // verilog/motorControl.v(38[12:27])
    defparam i1_4_lut_adj_1393.LUT_INIT = 16'hb3a2;
    SB_LUT4 i3_4_lut_adj_1394 (.I0(\PID_CONTROLLER.result [30]), .I1(n56_adj_3871), 
            .I2(\PID_CONTROLLER.result [28]), .I3(\PID_CONTROLLER.result [29]), 
            .O(n44118));   // verilog/motorControl.v(38[12:27])
    defparam i3_4_lut_adj_1394.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1395 (.I0(\PWMLimit[9] ), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n42629), .I3(n44118), .O(n387));   // verilog/motorControl.v(38[12:27])
    defparam i1_4_lut_adj_1395.LUT_INIT = 16'hb3a2;
    SB_LUT4 i6_3_lut (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [13]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n20_adj_3872));   // verilog/motorControl.v(37[31:51])
    defparam i6_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i2_3_lut_adj_1396 (.I0(\PID_CONTROLLER.result [10]), .I1(\PID_CONTROLLER.result [27]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n16_adj_3873));   // verilog/motorControl.v(37[31:51])
    defparam i2_3_lut_adj_1396.LUT_INIT = 16'h7e7e;
    SB_LUT4 i2_3_lut_adj_1397 (.I0(\PID_CONTROLLER.result [20]), .I1(\PID_CONTROLLER.result [15]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n10_adj_3874));   // verilog/motorControl.v(37[31:51])
    defparam i2_3_lut_adj_1397.LUT_INIT = 16'h7e7e;
    SB_LUT4 i4_3_lut (.I0(\PID_CONTROLLER.result [16]), .I1(\PID_CONTROLLER.result [19]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n12_adj_3875));   // verilog/motorControl.v(37[31:51])
    defparam i4_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i6_4_lut (.I0(\PID_CONTROLLER.result [12]), .I1(n12_adj_3875), 
            .I2(\PID_CONTROLLER.result [29]), .I3(pwm_23__N_2951[10]), .O(n14_adj_3876));   // verilog/motorControl.v(37[31:51])
    defparam i6_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i5_4_lut (.I0(\PID_CONTROLLER.result [17]), .I1(n10_adj_3874), 
            .I2(\PID_CONTROLLER.result [11]), .I3(pwm_23__N_2951[10]), .O(n13_adj_3877));   // verilog/motorControl.v(37[31:51])
    defparam i5_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i4_4_lut (.I0(\PID_CONTROLLER.result [24]), .I1(n13_adj_3877), 
            .I2(pwm_23__N_2951[10]), .I3(n14_adj_3876), .O(n18_adj_3878));   // verilog/motorControl.v(37[31:51])
    defparam i4_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 pwm_23__I_816_i5_2_lut (.I0(\PID_CONTROLLER.result [2]), .I1(pwm_23__N_2951[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3879));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31514_4_lut (.I0(n11_adj_12), .I1(n9_adj_13), .I2(n7_adj_3858), 
            .I3(n5_adj_3879), .O(n47028));
    defparam i31514_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 pwm_23__I_816_i8_3_lut (.I0(\pwm_23__N_2951[4] ), .I1(pwm_23__N_2951[8]), 
            .I2(n17_adj_3857), .I3(GND_net), .O(n8_adj_3882));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_23__I_816_i6_3_lut (.I0(pwm_23__N_2951[2]), .I1(pwm_23__N_2951[3]), 
            .I2(n7_adj_3858), .I3(GND_net), .O(n6_adj_3883));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_23__I_816_i16_3_lut (.I0(n8_adj_3882), .I1(pwm_23__N_2951[9]), 
            .I2(n19_adj_3856), .I3(GND_net), .O(n16_adj_3884));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31302_4_lut (.I0(n50_adj_3855), .I1(\PID_CONTROLLER.result [26]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [25]), .O(n46504));   // verilog/motorControl.v(37[10:27])
    defparam i31302_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 pwm_23__I_816_i4_3_lut (.I0(n46507), .I1(pwm_23__N_2951[1]), 
            .I2(\PID_CONTROLLER.result [1]), .I3(GND_net), .O(n4_adj_3885));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32649_3_lut (.I0(n4_adj_3885), .I1(\pwm_23__N_2951[5] ), .I2(n11_adj_12), 
            .I3(GND_net), .O(n48163));   // verilog/motorControl.v(37[31:51])
    defparam i32649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32650_3_lut (.I0(n48163), .I1(pwm_23__N_2951[6]), .I2(n13_adj_3842), 
            .I3(GND_net), .O(n48164));   // verilog/motorControl.v(37[31:51])
    defparam i32650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut (.I0(\PID_CONTROLLER.result [22]), .I1(n20_adj_3872), 
            .I2(\PID_CONTROLLER.result [30]), .I3(pwm_23__N_2951[10]), .O(n24_adj_3886));   // verilog/motorControl.v(37[31:51])
    defparam i10_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i8_4_lut (.I0(\PID_CONTROLLER.result [18]), .I1(n16_adj_3873), 
            .I2(\PID_CONTROLLER.result [26]), .I3(pwm_23__N_2951[10]), .O(n22_adj_3887));   // verilog/motorControl.v(37[31:51])
    defparam i8_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i9_4_lut (.I0(\PID_CONTROLLER.result [23]), .I1(n18_adj_3878), 
            .I2(\PID_CONTROLLER.result [14]), .I3(pwm_23__N_2951[10]), .O(n23_adj_3888));   // verilog/motorControl.v(37[31:51])
    defparam i9_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i7_3_lut (.I0(\PID_CONTROLLER.result [25]), .I1(\PID_CONTROLLER.result [28]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n21_adj_3889));   // verilog/motorControl.v(37[31:51])
    defparam i7_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i31504_4_lut (.I0(n17_adj_3857), .I1(n15_adj_14), .I2(n13_adj_3842), 
            .I3(n47028), .O(n47018));
    defparam i31504_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32951_4_lut (.I0(n16_adj_3884), .I1(n6_adj_3883), .I2(n19_adj_3856), 
            .I3(n47016), .O(n48465));   // verilog/motorControl.v(37[31:51])
    defparam i32951_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i31962_3_lut (.I0(n48164), .I1(\pwm_23__N_2951[7] ), .I2(n15_adj_14), 
            .I3(GND_net), .O(n47476));   // verilog/motorControl.v(37[31:51])
    defparam i31962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut (.I0(n21_adj_3889), .I1(n23_adj_3888), .I2(n22_adj_3887), 
            .I3(n24_adj_3886), .O(n44367));   // verilog/motorControl.v(37[31:51])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33084_4_lut (.I0(n47476), .I1(n48465), .I2(n19_adj_3856), 
            .I3(n47018), .O(n48598));   // verilog/motorControl.v(37[31:51])
    defparam i33084_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32141_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [29]), 
            .I2(\PID_CONTROLLER.result [30]), .I3(\PID_CONTROLLER.result [28]), 
            .O(n47655));
    defparam i32141_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 mult_12_i414_2_lut (.I0(\Kd[6] ), .I1(n67[11]), .I2(GND_net), 
            .I3(GND_net), .O(n616));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i56_3_lut  (.I0(n46504), .I1(\PID_CONTROLLER.result [27]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n56_adj_3891));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i56_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i60_4_lut  (.I0(\PID_CONTROLLER.result [28]), 
            .I1(\PID_CONTROLLER.result [30]), .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [29]), 
            .O(n60));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i60_4_lut .LUT_INIT = 16'h8f0e;
    SB_LUT4 i33056_4_lut (.I0(n48598), .I1(\PID_CONTROLLER.result [31]), 
            .I2(pwm_23__N_2951[10]), .I3(n44367), .O(pwm_23__N_2950));   // verilog/motorControl.v(37[31:51])
    defparam i33056_4_lut.LUT_INIT = 16'hcc8e;
    SB_LUT4 i32669_3_lut (.I0(n60), .I1(n56_adj_3891), .I2(n47655), .I3(GND_net), 
            .O(n48183));   // verilog/motorControl.v(37[10:27])
    defparam i32669_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_23__I_815_4_lut (.I0(n48183), .I1(pwm_23__N_2950), .I2(\deadband[9] ), 
            .I3(\PID_CONTROLLER.result [31]), .O(pwm_23__N_2948));   // verilog/motorControl.v(37[10:51])
    defparam pwm_23__I_815_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 LessThan_22_i17_2_lut (.I0(\PID_CONTROLLER.result [8]), .I1(n58[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3892));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1398 (.I0(\PID_CONTROLLER.result [28]), .I1(\PID_CONTROLLER.result [30]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(GND_net), .O(n42627));   // verilog/motorControl.v(38[12:27])
    defparam i2_3_lut_adj_1398.LUT_INIT = 16'h8080;
    SB_LUT4 i5_3_lut (.I0(\PID_CONTROLLER.result [20]), .I1(\PID_CONTROLLER.result [22]), 
            .I2(\PID_CONTROLLER.result [18]), .I3(GND_net), .O(n14_adj_3893));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6_4_lut_adj_1399 (.I0(\PID_CONTROLLER.result [23]), .I1(\PID_CONTROLLER.result [25]), 
            .I2(\PID_CONTROLLER.result [24]), .I3(\PID_CONTROLLER.result [19]), 
            .O(n15_adj_3894));
    defparam i6_4_lut_adj_1399.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1400 (.I0(n15_adj_3894), .I1(\PID_CONTROLLER.result [21]), 
            .I2(n14_adj_3893), .I3(\PID_CONTROLLER.result [17]), .O(n42695));
    defparam i8_4_lut_adj_1400.LUT_INIT = 16'h8000;
    SB_LUT4 i3_4_lut_adj_1401 (.I0(\PID_CONTROLLER.result [23]), .I1(\PID_CONTROLLER.result [24]), 
            .I2(\PID_CONTROLLER.result [22]), .I3(\PID_CONTROLLER.result [25]), 
            .O(n62_adj_3869));   // verilog/motorControl.v(31[14] 52[8])
    defparam i3_4_lut_adj_1401.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [19]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3895));   // verilog/motorControl.v(31[14] 52[8])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1402 (.I0(\PID_CONTROLLER.result [20]), .I1(\PID_CONTROLLER.result [17]), 
            .I2(\PID_CONTROLLER.result [18]), .I3(n6_adj_3895), .O(n49_adj_3870));   // verilog/motorControl.v(31[14] 52[8])
    defparam i4_4_lut_adj_1402.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_22_i13_2_lut (.I0(\PID_CONTROLLER.result [6]), .I1(n58[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_3896));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i7_2_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n58[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3897));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i19_2_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n58[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3898));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_2_lut (.I0(\PID_CONTROLLER.result [14]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_3899));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1403 (.I0(\PID_CONTROLLER.result [11]), .I1(\PID_CONTROLLER.result [27]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(\PID_CONTROLLER.result [10]), 
            .O(n24_adj_3900));
    defparam i10_4_lut_adj_1403.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_22_i5_2_lut (.I0(\PID_CONTROLLER.result [2]), .I1(n58[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3901));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31442_4_lut (.I0(n11_adj_15), .I1(n9_adj_16), .I2(n7_adj_3897), 
            .I3(n5_adj_3901), .O(n46955));
    defparam i31442_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_22_i4_4_lut (.I0(n58[0]), .I1(n58[1]), .I2(\PID_CONTROLLER.result [1]), 
            .I3(\PID_CONTROLLER.result [0]), .O(n4_adj_3904));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i32643_3_lut (.I0(n4_adj_3904), .I1(n415), .I2(n11_adj_15), 
            .I3(GND_net), .O(n48157));   // verilog/motorControl.v(40[21:37])
    defparam i32643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32644_3_lut (.I0(n48157), .I1(n58[6]), .I2(n13_adj_3896), 
            .I3(GND_net), .O(n48158));   // verilog/motorControl.v(40[21:37])
    defparam i32644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(\PID_CONTROLLER.result [27]), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(GND_net), .O(n10_adj_3905));   // verilog/motorControl.v(31[14] 52[8])
    defparam i1_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i8_4_lut_adj_1404 (.I0(\PID_CONTROLLER.result [30]), .I1(n49_adj_3870), 
            .I2(\PID_CONTROLLER.result [12]), .I3(\PID_CONTROLLER.result [28]), 
            .O(n22_adj_3906));
    defparam i8_4_lut_adj_1404.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(\PID_CONTROLLER.result [16]), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [11]), .I3(GND_net), .O(n12_adj_3907));   // verilog/motorControl.v(31[14] 52[8])
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7_4_lut (.I0(n58[10]), .I1(\PID_CONTROLLER.result [12]), .I2(\PID_CONTROLLER.result [26]), 
            .I3(n10_adj_3905), .O(n16_adj_3908));   // verilog/motorControl.v(31[14] 52[8])
    defparam i7_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i12_4_lut (.I0(\PID_CONTROLLER.result [29]), .I1(n24_adj_3900), 
            .I2(n18_adj_3899), .I3(n62_adj_3869), .O(n26_adj_3909));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31469_4_lut (.I0(n42695), .I1(n16_adj_3908), .I2(n12_adj_3907), 
            .I3(n42627), .O(n46613));   // verilog/motorControl.v(31[14] 52[8])
    defparam i31469_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(\PID_CONTROLLER.result [26]), .I1(n22_adj_3906), 
            .I2(n58[10]), .I3(GND_net), .O(n25_adj_3910));
    defparam i11_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 LessThan_22_i6_3_lut (.I0(n58[2]), .I1(n58[3]), .I2(n7_adj_3897), 
            .I3(GND_net), .O(n6_adj_3911));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32835_3_lut (.I0(n6_adj_3911), .I1(n416), .I2(n9_adj_16), 
            .I3(GND_net), .O(n48349));   // verilog/motorControl.v(40[21:37])
    defparam i32835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32836_3_lut (.I0(n48349), .I1(n58[8]), .I2(n17_adj_3892), 
            .I3(GND_net), .O(n48350));   // verilog/motorControl.v(40[21:37])
    defparam i32836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31434_4_lut (.I0(n17_adj_3892), .I1(n15_adj_17), .I2(n13_adj_3896), 
            .I3(n46955), .O(n46947));
    defparam i31434_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31972_3_lut (.I0(n48158), .I1(n413), .I2(n15_adj_17), .I3(GND_net), 
            .O(n47486));   // verilog/motorControl.v(40[21:37])
    defparam i31972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32626_3_lut (.I0(n48350), .I1(n58[9]), .I2(n19_adj_3898), 
            .I3(GND_net), .O(n48140));   // verilog/motorControl.v(40[21:37])
    defparam i32626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28_4_lut (.I0(n25_adj_3910), .I1(n46613), .I2(\PID_CONTROLLER.result [13]), 
            .I3(n26_adj_3909), .O(n20_adj_3913));   // verilog/motorControl.v(31[14] 52[8])
    defparam i28_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 i32677_4_lut (.I0(n48140), .I1(n47486), .I2(n19_adj_3898), 
            .I3(n46947), .O(n48191));   // verilog/motorControl.v(40[21:37])
    defparam i32677_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32418_4_lut (.I0(n48191), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n58[10]), .I3(n20_adj_3913), .O(n421));   // verilog/motorControl.v(40[21:37])
    defparam i32418_4_lut.LUT_INIT = 16'h8ecc;
    SB_LUT4 mux_24_i1_3_lut (.I0(\PID_CONTROLLER.result [0]), .I1(n58[0]), 
            .I2(n421), .I3(GND_net), .O(n471));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_12_i351_2_lut (.I0(\Kd[5] ), .I1(n67[12]), .I2(GND_net), 
            .I3(GND_net), .O(n522_adj_3834));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i416_2_lut (.I0(\Kd[6] ), .I1(n67[12]), .I2(GND_net), 
            .I3(GND_net), .O(n619_adj_3833));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i481_2_lut (.I0(\Kd[7] ), .I1(n67[12]), .I2(GND_net), 
            .I3(GND_net), .O(n716_adj_3832));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i93_2_lut (.I0(\Kd[1] ), .I1(n67[13]), .I2(GND_net), 
            .I3(GND_net), .O(n137_adj_3831));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i30_2_lut (.I0(\Kd[0] ), .I1(n67[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_3830));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i158_2_lut (.I0(\Kd[2] ), .I1(n67[13]), .I2(GND_net), 
            .I3(GND_net), .O(n234_adj_3829));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i223_2_lut (.I0(\Kd[3] ), .I1(n67[13]), .I2(GND_net), 
            .I3(GND_net), .O(n331_adj_3828));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i288_2_lut (.I0(\Kd[4] ), .I1(n67[13]), .I2(GND_net), 
            .I3(GND_net), .O(n428_adj_3827));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i288_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i353_2_lut (.I0(\Kd[5] ), .I1(n67[13]), .I2(GND_net), 
            .I3(GND_net), .O(n525_adj_3826));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i418_2_lut (.I0(\Kd[6] ), .I1(n67[13]), .I2(GND_net), 
            .I3(GND_net), .O(n622_adj_3825));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i483_2_lut (.I0(\Kd[7] ), .I1(n67[13]), .I2(GND_net), 
            .I3(GND_net), .O(n719_adj_3824));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i479_2_lut (.I0(\Kd[7] ), .I1(n67[11]), .I2(GND_net), 
            .I3(GND_net), .O(n713));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[22]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3823));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_3822));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_3821));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i95_2_lut (.I0(\Kd[1] ), .I1(n67[14]), .I2(GND_net), 
            .I3(GND_net), .O(n140_adj_3820));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i32_2_lut (.I0(\Kd[0] ), .I1(n67[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_3819));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i160_2_lut (.I0(\Kd[2] ), .I1(n67[14]), .I2(GND_net), 
            .I3(GND_net), .O(n237_adj_3818));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i225_2_lut (.I0(\Kd[3] ), .I1(n67[14]), .I2(GND_net), 
            .I3(GND_net), .O(n334_adj_3817));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i290_2_lut (.I0(\Kd[4] ), .I1(n67[14]), .I2(GND_net), 
            .I3(GND_net), .O(n431_adj_3816));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i355_2_lut (.I0(\Kd[5] ), .I1(n67[14]), .I2(GND_net), 
            .I3(GND_net), .O(n528_adj_3815));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i420_2_lut (.I0(\Kd[6] ), .I1(n67[14]), .I2(GND_net), 
            .I3(GND_net), .O(n625_adj_3814));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i485_2_lut (.I0(\Kd[7] ), .I1(n67[14]), .I2(GND_net), 
            .I3(GND_net), .O(n722_adj_3813));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i5_1_lut (.I0(\PWMLimit[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[4]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i6_1_lut (.I0(\PWMLimit[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[5]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i49_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n72));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i49_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[23]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i98_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n145_adj_3809));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i98_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i147_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n218_adj_3808));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i147_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 unary_minus_21_inv_0_i7_1_lut (.I0(\PWMLimit[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[6]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i196_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n291));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i196_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i245_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n364_adj_3806));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i245_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i294_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n437_adj_3805));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i294_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_12_i69_2_lut (.I0(\Kd[1] ), .I1(n67[1]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_3804));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i6_2_lut (.I0(\Kd[0] ), .I1(n67[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3803));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i343_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n510_adj_3802));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i343_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_12_i134_2_lut (.I0(\Kd[2] ), .I1(n67[1]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_3801));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i392_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n583_adj_3800));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i392_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 unary_minus_21_inv_0_i8_1_lut (.I0(\PWMLimit[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[7]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i199_2_lut (.I0(\Kd[3] ), .I1(n67[1]), .I2(GND_net), 
            .I3(GND_net), .O(n295_adj_3797));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i199_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n76[0]));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n282[0]));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3794));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3793));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i264_2_lut (.I0(\Kd[4] ), .I1(n67[1]), .I2(GND_net), 
            .I3(GND_net), .O(n392_adj_3792));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i264_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i97_2_lut (.I0(\Kd[1] ), .I1(n67[15]), .I2(GND_net), 
            .I3(GND_net), .O(n143_adj_3791));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i97_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i34_2_lut (.I0(\Kd[0] ), .I1(n67[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_3790));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i146_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n216_adj_3788));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i162_2_lut (.I0(\Kd[2] ), .I1(n67[15]), .I2(GND_net), 
            .I3(GND_net), .O(n240_adj_3787));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i329_2_lut (.I0(\Kd[5] ), .I1(n67[1]), .I2(GND_net), 
            .I3(GND_net), .O(n489_adj_3786));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i329_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i211_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n313_adj_3785));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i394_2_lut (.I0(\Kd[6] ), .I1(n67[1]), .I2(GND_net), 
            .I3(GND_net), .O(n586_adj_3784));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i227_2_lut (.I0(\Kd[3] ), .I1(n67[15]), .I2(GND_net), 
            .I3(GND_net), .O(n337_adj_3783));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i276_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n410_adj_3782));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i292_2_lut (.I0(\Kd[4] ), .I1(n67[15]), .I2(GND_net), 
            .I3(GND_net), .O(n434_adj_3781));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i341_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n507_adj_3780));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i459_2_lut (.I0(\Kd[7] ), .I1(n67[1]), .I2(GND_net), 
            .I3(GND_net), .O(n683_adj_3779));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33809_4_lut (.I0(n46608), .I1(n43470), .I2(n43441), .I3(n17_adj_3482), 
            .O(n42680));
    defparam i33809_4_lut.LUT_INIT = 16'hddfc;
    SB_LUT4 PHASES_5__I_0_i6_4_lut (.I0(PHASES_5__N_3039[4]), .I1(n22379), 
            .I2(n17_adj_3482), .I3(n878), .O(PHASES_5__N_2779[5]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i6_4_lut.LUT_INIT = 16'ha303;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n604_adj_3778));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i357_2_lut (.I0(\Kd[5] ), .I1(n67[15]), .I2(GND_net), 
            .I3(GND_net), .O(n531_adj_3777));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i1_1_lut (.I0(\PWMLimit[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[0]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n701_adj_3776));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i9_1_lut (.I0(\PWMLimit[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[8]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i2_1_lut (.I0(\PWMLimit[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[1]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i422_2_lut (.I0(\Kd[6] ), .I1(n67[15]), .I2(GND_net), 
            .I3(GND_net), .O(n628_adj_3774));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i487_2_lut (.I0(\Kd[7] ), .I1(n67[15]), .I2(GND_net), 
            .I3(GND_net), .O(n725_adj_3773));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3772));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i6_3_lut_3_lut (.I0(\PWMLimit[3] ), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(GND_net), .O(n6_adj_3863));   // verilog/motorControl.v(38[12:27])
    defparam LessThan_20_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i31473_3_lut_4_lut (.I0(\PWMLimit[3] ), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(\PWMLimit[2] ), .O(n46986));   // verilog/motorControl.v(38[12:27])
    defparam i31473_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_21_inv_0_i32_1_lut (.I0(\PWMLimit[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3771));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_3769));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_3767));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[5]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[18]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i27960_3_lut (.I0(hall2), .I1(hall1), .I2(hall3), .I3(GND_net), 
            .O(n43468));
    defparam i27960_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i27961_3_lut (.I0(hall2), .I1(hall3), .I2(hall1), .I3(GND_net), 
            .O(n43470));
    defparam i27961_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i33811_4_lut (.I0(n46609), .I1(n43470), .I2(n43468), .I3(n17_adj_3482), 
            .O(n42681));
    defparam i33811_4_lut.LUT_INIT = 16'hddfc;
    SB_LUT4 i10301_4_lut (.I0(n878), .I1(PHASES_5__N_3039[4]), .I2(n17_adj_3482), 
            .I3(n22379), .O(PHASES_5__N_2779[4]));   // verilog/motorControl.v(77[14] 98[8])
    defparam i10301_4_lut.LUT_INIT = 16'h0cac;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[6]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_adj_1405 (.I0(n881_adj_3481), .I1(n878), .I2(n934), 
            .I3(n19616), .O(n43907));
    defparam i3_4_lut_adj_1405.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_4_lut_adj_1406 (.I0(PHASES_5__N_3039[3]), .I1(n43907), .I2(n42708), 
            .I3(n880), .O(n23630));
    defparam i1_4_lut_adj_1406.LUT_INIT = 16'hccc8;
    SB_LUT4 mult_14_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 PHASES_5__I_0_i4_4_lut (.I0(PHASES_5__N_3039[2]), .I1(PHASES_5__N_3039[3]), 
            .I2(n17_adj_3482), .I3(n878), .O(PHASES_5__N_2779[3]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i4_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 mult_14_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6304_2_lut (.I0(hall1), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n19954));   // verilog/motorControl.v(87[7] 89[10])
    defparam i6304_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[7]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6499_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(PHASES_5__N_3039[3]));   // verilog/motorControl.v(87[7] 89[10])
    defparam i6499_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31_4_lut (.I0(n19954), .I1(n880), .I2(hall3), .I3(PHASES_5__N_3039[4]), 
            .O(n43507));
    defparam i31_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[8]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30_4_lut (.I0(n46611), .I1(n934), .I2(n17_adj_3482), .I3(n43507), 
            .O(n15_adj_3765));
    defparam i30_4_lut.LUT_INIT = 16'h5f5c;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[19]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 PHASES_5__I_0_i3_4_lut (.I0(PHASES_5__N_3039[3]), .I1(PHASES_5__N_3039[2]), 
            .I2(n17_adj_3482), .I3(n878), .O(PHASES_5__N_2779[2]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i3_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[9]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1407 (.I0(n20463), .I1(n17_adj_3482), .I2(n42708), 
            .I3(n4_adj_3914), .O(n23622));
    defparam i1_4_lut_adj_1407.LUT_INIT = 16'hfa32;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[10]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut (.I0(hall2), .I1(n19326), .I2(GND_net), .I3(GND_net), 
            .O(n902_adj_3915));   // verilog/motorControl.v(84[10:34])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[11]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut_adj_1408 (.I0(n880), .I1(PHASES_5__N_3039[4]), .I2(n902_adj_3915), 
            .I3(hall3), .O(n20463));   // verilog/motorControl.v(68[7] 70[10])
    defparam i2_4_lut_adj_1408.LUT_INIT = 16'hfafe;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[20]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i83_2_lut (.I0(\Kd[1] ), .I1(n67[8]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_3405));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i20_2_lut (.I0(\Kd[0] ), .I1(n67[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3404));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i73_3_lut (.I0(pwm[23]), .I1(n29), .I2(n30), .I3(GND_net), 
            .O(n878));   // verilog/motorControl.v(77[19:44])
    defparam i73_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i75_2_lut (.I0(hall1), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n880));   // verilog/motorControl.v(78[10:25])
    defparam i75_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i76_2_lut (.I0(n880), .I1(hall3), .I2(GND_net), .I3(GND_net), 
            .O(n881_adj_3481));   // verilog/motorControl.v(78[10:34])
    defparam i76_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1409 (.I0(hall1), .I1(hall3), .I2(GND_net), .I3(GND_net), 
            .O(n19326));   // verilog/motorControl.v(84[10:34])
    defparam i1_2_lut_adj_1409.LUT_INIT = 16'h2222;
    SB_LUT4 i6495_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(PHASES_5__N_3039[1]));   // verilog/motorControl.v(93[7] 95[10])
    defparam i6495_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_adj_1410 (.I0(hall2), .I1(PHASES_5__N_3039[1]), .I2(GND_net), 
            .I3(GND_net), .O(n934));   // verilog/motorControl.v(93[10:35])
    defparam i2_2_lut_adj_1410.LUT_INIT = 16'h4444;
    SB_LUT4 i88_2_lut (.I0(hall1), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(PHASES_5__N_3039[4]));   // verilog/motorControl.v(87[10:25])
    defparam i88_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5_4_lut_adj_1411 (.I0(n48193), .I1(pwm[21]), .I2(pwm[8]), 
            .I3(\pwm_count[8] ), .O(n20_adj_3918));
    defparam i5_4_lut_adj_1411.LUT_INIT = 16'hecfe;
    SB_LUT4 i11_4_lut (.I0(pwm[11]), .I1(pwm[17]), .I2(pwm[19]), .I3(pwm[12]), 
            .O(n26_adj_3919));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1412 (.I0(pwm[16]), .I1(pwm[10]), .I2(pwm[14]), 
            .I3(pwm[9]), .O(n24_adj_3920));
    defparam i9_4_lut_adj_1412.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1413 (.I0(pwm[13]), .I1(n26_adj_3919), .I2(n20_adj_3918), 
            .I3(pwm[22]), .O(n28_adj_3921));
    defparam i13_4_lut_adj_1413.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_3_lut (.I0(pwm[15]), .I1(pwm[18]), .I2(pwm[20]), .I3(GND_net), 
            .O(n23_adj_3922));
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1414 (.I0(pwm[23]), .I1(n23_adj_3922), .I2(n28_adj_3921), 
            .I3(n24_adj_3920), .O(n17_adj_3482));   // verilog/motorControl.v(58[9:32])
    defparam i1_4_lut_adj_1414.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_1415 (.I0(n43915), .I1(PHASES_5__N_3039[1]), .I2(n878), 
            .I3(n20463), .O(n23562));
    defparam i1_4_lut_adj_1415.LUT_INIT = 16'haa8a;
    SB_LUT4 i10317_4_lut (.I0(n46593), .I1(n16802), .I2(n17_adj_3482), 
            .I3(n19326), .O(PHASES_5__N_2779[0]));   // verilog/motorControl.v(77[14] 98[8])
    defparam i10317_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 mult_14_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_3764));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3403));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_3402));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31475_3_lut_3_lut (.I0(n58[10]), .I1(n421), .I2(\PID_CONTROLLER.result [17]), 
            .I3(GND_net), .O(n46604));   // verilog/motorControl.v(40[28:37])
    defparam i31475_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[12]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[21]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31792_3_lut_3_lut (.I0(n58[10]), .I1(n421), .I2(\PID_CONTROLLER.result [18]), 
            .I3(GND_net), .O(n46606));   // verilog/motorControl.v(40[28:37])
    defparam i31792_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 i31409_3_lut_3_lut (.I0(n58[10]), .I1(n421), .I2(\PID_CONTROLLER.result [19]), 
            .I3(GND_net), .O(n46565));   // verilog/motorControl.v(40[28:37])
    defparam i31409_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 mult_12_i148_2_lut (.I0(\Kd[2] ), .I1(n67[8]), .I2(GND_net), 
            .I3(GND_net), .O(n219_adj_3400));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31541_3_lut_3_lut (.I0(n58[10]), .I1(n421), .I2(\PID_CONTROLLER.result [20]), 
            .I3(GND_net), .O(n46567));   // verilog/motorControl.v(40[28:37])
    defparam i31541_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 mult_10_i150_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n222_adj_3399));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[13]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i213_2_lut (.I0(\Kd[3] ), .I1(n67[8]), .I2(GND_net), 
            .I3(GND_net), .O(n316_adj_3398));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i215_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n319_adj_3397));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i278_2_lut (.I0(\Kd[4] ), .I1(n67[8]), .I2(GND_net), 
            .I3(GND_net), .O(n413_adj_3396));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i280_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n416_adj_3395));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i343_2_lut (.I0(\Kd[5] ), .I1(n67[8]), .I2(GND_net), 
            .I3(GND_net), .O(n510_adj_3394));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n513_adj_3393));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[14]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[22]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31539_3_lut_3_lut (.I0(n58[10]), .I1(n421), .I2(\PID_CONTROLLER.result [23]), 
            .I3(GND_net), .O(n46573));   // verilog/motorControl.v(40[28:37])
    defparam i31539_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 i31544_3_lut_3_lut (.I0(n58[10]), .I1(n421), .I2(\PID_CONTROLLER.result [22]), 
            .I3(GND_net), .O(n46571));   // verilog/motorControl.v(40[28:37])
    defparam i31544_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 i31535_3_lut_3_lut (.I0(n58[10]), .I1(n421), .I2(\PID_CONTROLLER.result [21]), 
            .I3(GND_net), .O(n46569));   // verilog/motorControl.v(40[28:37])
    defparam i31535_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 mult_12_i408_2_lut (.I0(\Kd[6] ), .I1(n67[8]), .I2(GND_net), 
            .I3(GND_net), .O(n607_adj_3389));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n610_adj_3388));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[15]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i473_2_lut (.I0(\Kd[7] ), .I1(n67[8]), .I2(GND_net), 
            .I3(GND_net), .O(n704_adj_3386));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i475_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n707_adj_3385));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i99_2_lut (.I0(\Kd[1] ), .I1(n67[16]), .I2(GND_net), 
            .I3(GND_net), .O(n146_adj_3762));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i99_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i36_2_lut (.I0(\Kd[0] ), .I1(n67[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_3761));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1416 (.I0(Kd_delay_counter[5]), .I1(Kd_delay_counter[3]), 
            .I2(Kd_delay_counter[6]), .I3(Kd_delay_counter[4]), .O(n12_adj_3923));   // verilog/motorControl.v(49[10:29])
    defparam i5_4_lut_adj_1416.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[16]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1417 (.I0(Kd_delay_counter[1]), .I1(n12_adj_3923), 
            .I2(Kd_delay_counter[2]), .I3(Kd_delay_counter[0]), .O(n44066));   // verilog/motorControl.v(49[10:29])
    defparam i6_4_lut_adj_1417.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_14_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[17]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i164_2_lut (.I0(\Kd[2] ), .I1(n67[16]), .I2(GND_net), 
            .I3(GND_net), .O(n243_adj_3760));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i164_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n70[23]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i229_2_lut (.I0(\Kd[3] ), .I1(n67[16]), .I2(GND_net), 
            .I3(GND_net), .O(n340_adj_3758));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[18]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[19]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i294_2_lut (.I0(\Kd[4] ), .I1(n67[16]), .I2(GND_net), 
            .I3(GND_net), .O(n437_adj_3756));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i85_2_lut (.I0(\Kd[1] ), .I1(n67[9]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i22_2_lut (.I0(\Kd[0] ), .I1(n67[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_3375));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i107_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n158));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i44_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n65));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i150_2_lut (.I0(\Kd[2] ), .I1(n67[9]), .I2(GND_net), 
            .I3(GND_net), .O(n222));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i172_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n255));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3754));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i215_2_lut (.I0(\Kd[3] ), .I1(n67[9]), .I2(GND_net), 
            .I3(GND_net), .O(n319));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3753));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i237_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n352));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i280_2_lut (.I0(\Kd[4] ), .I1(n67[9]), .I2(GND_net), 
            .I3(GND_net), .O(n416_c));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n449_adj_3374));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i345_2_lut (.I0(\Kd[5] ), .I1(n67[9]), .I2(GND_net), 
            .I3(GND_net), .O(n513));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n546));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i410_2_lut (.I0(\Kd[6] ), .I1(n67[9]), .I2(GND_net), 
            .I3(GND_net), .O(n610));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i359_2_lut (.I0(\Kd[5] ), .I1(n67[16]), .I2(GND_net), 
            .I3(GND_net), .O(n534_adj_3752));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i432_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n643));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i144_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n213_adj_3750));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i209_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n310_adj_3747));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i274_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n407_adj_3745));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i339_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n504_adj_3743));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i339_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i475_2_lut (.I0(\Kd[7] ), .I1(n67[9]), .I2(GND_net), 
            .I3(GND_net), .O(n707));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n601_adj_3741));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i424_2_lut (.I0(\Kd[6] ), .I1(n67[16]), .I2(GND_net), 
            .I3(GND_net), .O(n631_adj_3740));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i489_2_lut (.I0(\Kd[7] ), .I1(n67[16]), .I2(GND_net), 
            .I3(GND_net), .O(n728_adj_3738));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n698_adj_3737));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i497_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_c));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i148_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n219));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i213_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n316));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i278_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n413_c));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i101_2_lut (.I0(\Kd[1] ), .I1(n67[17]), .I2(GND_net), 
            .I3(GND_net), .O(n149_adj_3733));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i343_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n510));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i38_2_lut (.I0(\Kd[0] ), .I1(n67[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_3732));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n607));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i473_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n704));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i166_2_lut (.I0(\Kd[2] ), .I1(n67[17]), .I2(GND_net), 
            .I3(GND_net), .O(n246_adj_3731));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[20]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i231_2_lut (.I0(\Kd[3] ), .I1(n67[17]), .I2(GND_net), 
            .I3(GND_net), .O(n343_adj_3730));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i87_2_lut (.I0(\Kd[1] ), .I1(n67[10]), .I2(GND_net), 
            .I3(GND_net), .O(n128));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i87_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i24_2_lut (.I0(\Kd[0] ), .I1(n67[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i152_2_lut (.I0(\Kd[2] ), .I1(n67[10]), .I2(GND_net), 
            .I3(GND_net), .O(n225));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i217_2_lut (.I0(\Kd[3] ), .I1(n67[10]), .I2(GND_net), 
            .I3(GND_net), .O(n322));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i282_2_lut (.I0(\Kd[4] ), .I1(n67[10]), .I2(GND_net), 
            .I3(GND_net), .O(n419_adj_3371));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i347_2_lut (.I0(\Kd[5] ), .I1(n67[10]), .I2(GND_net), 
            .I3(GND_net), .O(n516));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i296_2_lut (.I0(\Kd[4] ), .I1(n67[17]), .I2(GND_net), 
            .I3(GND_net), .O(n440_adj_3729));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i412_2_lut (.I0(\Kd[6] ), .I1(n67[10]), .I2(GND_net), 
            .I3(GND_net), .O(n613));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[21]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i477_2_lut (.I0(\Kd[7] ), .I1(n67[10]), .I2(GND_net), 
            .I3(GND_net), .O(n710));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i361_2_lut (.I0(\Kd[5] ), .I1(n67[17]), .I2(GND_net), 
            .I3(GND_net), .O(n537_adj_3728));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i426_2_lut (.I0(\Kd[6] ), .I1(n67[17]), .I2(GND_net), 
            .I3(GND_net), .O(n634_adj_3727));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i426_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i491_2_lut (.I0(\Kd[7] ), .I1(n67[17]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_3726));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i93_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n137_adj_3725));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i158_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n234_adj_3724));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3723));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3722));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i142_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n210_adj_3721));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i223_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n331));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i207_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n307_adj_3720));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i272_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n404_adj_3719));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i337_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n501_adj_3718));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i288_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n428));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i288_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n598_adj_3717));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n695_adj_3716));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n525_adj_3715));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n622));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i483_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n719));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i103_2_lut (.I0(\Kd[1] ), .I1(n67[18]), .I2(GND_net), 
            .I3(GND_net), .O(n152_adj_3714));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i40_2_lut (.I0(\Kd[0] ), .I1(n67[19]), .I2(GND_net), 
            .I3(GND_net), .O(n59_adj_3713));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i168_2_lut (.I0(\Kd[2] ), .I1(n67[18]), .I2(GND_net), 
            .I3(GND_net), .O(n249_adj_3712));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i168_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i233_2_lut (.I0(\Kd[3] ), .I1(n67[18]), .I2(GND_net), 
            .I3(GND_net), .O(n346_adj_3711));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3710));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i298_2_lut (.I0(\Kd[4] ), .I1(n67[18]), .I2(GND_net), 
            .I3(GND_net), .O(n443_adj_3709));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i363_2_lut (.I0(\Kd[5] ), .I1(n67[18]), .I2(GND_net), 
            .I3(GND_net), .O(n540_adj_3708));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_3707));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_3705));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_3703));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i428_2_lut (.I0(\Kd[6] ), .I1(n67[18]), .I2(GND_net), 
            .I3(GND_net), .O(n637_adj_3701));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i493_2_lut (.I0(\Kd[7] ), .I1(n67[18]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_3700));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i493_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3698));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3697));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i140_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n207_adj_3696));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i205_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n304_adj_3695));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i205_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i270_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n401_adj_3694));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i2_2_lut (.I0(\Kd[0] ), .I1(n67[0]), .I2(GND_net), 
            .I3(GND_net), .O(n191[0]));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i105_2_lut (.I0(\Kd[1] ), .I1(n67[19]), .I2(GND_net), 
            .I3(GND_net), .O(n155_adj_3693));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i42_2_lut (.I0(\Kd[0] ), .I1(n67[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_3692));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i335_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n498_adj_3690));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i335_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n595_adj_3688));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n692_adj_3687));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i170_2_lut (.I0(\Kd[2] ), .I1(n67[19]), .I2(GND_net), 
            .I3(GND_net), .O(n252_adj_3686));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i170_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i235_2_lut (.I0(\Kd[3] ), .I1(n67[19]), .I2(GND_net), 
            .I3(GND_net), .O(n349_adj_3685));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i300_2_lut (.I0(\Kd[4] ), .I1(n67[19]), .I2(GND_net), 
            .I3(GND_net), .O(n446_adj_3683));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i365_2_lut (.I0(\Kd[5] ), .I1(n67[19]), .I2(GND_net), 
            .I3(GND_net), .O(n543_adj_3682));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\Kd[3] ), .I1(n67[25]), .I2(n4_adj_3924), 
            .I3(n10115[1]), .O(n10850[2]));   // verilog/motorControl.v(36[26:45])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_12_i430_2_lut (.I0(\Kd[6] ), .I1(n67[19]), .I2(GND_net), 
            .I3(GND_net), .O(n640_adj_3681));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i430_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22529_3_lut_4_lut (.I0(n16641[2]), .I1(\Kp[4] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n6_adj_3925), .O(n8_adj_3926));   // verilog/motorControl.v(36[17:23])
    defparam i22529_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i2_3_lut_4_lut_adj_1418 (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(\Kp[4] ), .I3(n6_adj_3925), .O(n8_adj_3927));   // verilog/motorControl.v(36[17:23])
    defparam i2_3_lut_4_lut_adj_1418.LUT_INIT = 16'hb748;
    SB_LUT4 i22688_3_lut_4_lut (.I0(n16654[1]), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n4_adj_3928), .O(n6_adj_3925));   // verilog/motorControl.v(36[17:23])
    defparam i22688_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i22513_4_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n16641[0]), .I3(n36197), .O(n4_adj_3928));   // verilog/motorControl.v(36[17:23])
    defparam i22513_4_lut_4_lut.LUT_INIT = 16'hf8a0;
    SB_LUT4 i22899_2_lut_3_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(\Kp[1] ), .I3(GND_net), .O(n36197));   // verilog/motorControl.v(36[17:23])
    defparam i22899_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut (.I0(n16641[2]), .I1(\Kp[4] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n6_adj_3925), .O(n16641[3]));   // verilog/motorControl.v(36[17:23])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h956a;
    SB_LUT4 mult_12_i495_2_lut (.I0(\Kd[7] ), .I1(n67[19]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_3680));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n4_adj_3928), .I3(n38421), .O(n7_adj_3929));   // verilog/motorControl.v(36[17:23])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h78b4;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1419 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n4_adj_3928), .I3(n16654[1]), .O(n16641[2]));   // verilog/motorControl.v(36[17:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1419.LUT_INIT = 16'h8778;
    SB_LUT4 mult_12_i107_2_lut (.I0(\Kd[1] ), .I1(n67[20]), .I2(GND_net), 
            .I3(GND_net), .O(n158_adj_3679));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i44_2_lut (.I0(\Kd[0] ), .I1(n67[21]), .I2(GND_net), 
            .I3(GND_net), .O(n65_adj_3678));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i172_2_lut (.I0(\Kd[2] ), .I1(n67[20]), .I2(GND_net), 
            .I3(GND_net), .O(n255_adj_3677));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i237_2_lut (.I0(\Kd[3] ), .I1(n67[20]), .I2(GND_net), 
            .I3(GND_net), .O(n352_adj_3676));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i302_2_lut (.I0(\Kd[4] ), .I1(n67[20]), .I2(GND_net), 
            .I3(GND_net), .O(n449_adj_3675));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i367_2_lut (.I0(\Kd[5] ), .I1(n67[20]), .I2(GND_net), 
            .I3(GND_net), .O(n546_adj_3674));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i432_2_lut (.I0(\Kd[6] ), .I1(n67[20]), .I2(GND_net), 
            .I3(GND_net), .O(n643_adj_3673));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3672));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3671));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i497_2_lut (.I0(\Kd[7] ), .I1(n67[20]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_3670));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n204_adj_3669));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i203_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n301_adj_3668));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i268_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n398_adj_3667));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i333_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n495_adj_3666));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i333_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n592_adj_3665));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n689_adj_3664));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i109_2_lut (.I0(\Kd[1] ), .I1(n67[21]), .I2(GND_net), 
            .I3(GND_net), .O(n161_adj_3663));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i46_2_lut (.I0(\Kd[0] ), .I1(n67[22]), .I2(GND_net), 
            .I3(GND_net), .O(n68_adj_3662));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22836_3_lut_4_lut (.I0(n10850[2]), .I1(\Kd[4] ), .I2(n67[25]), 
            .I3(n6_adj_3930), .O(n8_adj_3931));   // verilog/motorControl.v(36[26:45])
    defparam i22836_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i2_3_lut_4_lut_adj_1420 (.I0(\Kd[5] ), .I1(n67[25]), .I2(\Kd[4] ), 
            .I3(n6_adj_3930), .O(n8_adj_3932));   // verilog/motorControl.v(36[26:45])
    defparam i2_3_lut_4_lut_adj_1420.LUT_INIT = 16'hb748;
    SB_LUT4 i22828_3_lut_4_lut (.I0(n10115[1]), .I1(\Kd[3] ), .I2(n67[25]), 
            .I3(n4_adj_3924), .O(n6_adj_3930));   // verilog/motorControl.v(36[26:45])
    defparam i22828_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i22732_2_lut_3_lut (.I0(\Kd[0] ), .I1(n67[25]), .I2(\Kd[1] ), 
            .I3(GND_net), .O(n36328));   // verilog/motorControl.v(36[26:45])
    defparam i22732_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut_adj_1421 (.I0(n10850[2]), .I1(\Kd[4] ), .I2(n67[25]), 
            .I3(n6_adj_3930), .O(n10115[3]));   // verilog/motorControl.v(36[26:45])
    defparam i1_3_lut_4_lut_adj_1421.LUT_INIT = 16'h956a;
    SB_LUT4 LessThan_4_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_3933));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i4_2_lut_adj_1422 (.I0(n19_c), .I1(n25), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_3934));   // verilog/motorControl.v(33[38:63])
    defparam i4_2_lut_adj_1422.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1423 (.I0(n33_adj_3383), .I1(n43), .I2(n27), 
            .I3(n35_adj_3382), .O(n24_adj_3935));   // verilog/motorControl.v(33[38:63])
    defparam i10_4_lut_adj_1423.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1424 (.I0(n41_adj_3372), .I1(n45), .I2(n31_adj_3387), 
            .I3(n23_adj_3407), .O(n22_adj_3936));   // verilog/motorControl.v(33[38:63])
    defparam i8_4_lut_adj_1424.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1425 (.I0(n29_adj_3391), .I1(n24_adj_3935), .I2(n18_adj_3934), 
            .I3(n37_adj_3378), .O(n26_adj_3937));   // verilog/motorControl.v(33[38:63])
    defparam i12_4_lut_adj_1425.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1426 (.I0(n21_c), .I1(n26_adj_3937), .I2(n22_adj_3936), 
            .I3(n39_adj_3376), .O(n44028));   // verilog/motorControl.v(33[38:63])
    defparam i13_4_lut_adj_1426.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_4_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(IntegralLimit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3938));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(IntegralLimit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3939));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(IntegralLimit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3940));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32321_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3940), 
            .I2(IntegralLimit[9]), .I3(n9_adj_3939), .O(n47835));
    defparam i32321_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32317_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[10]), 
            .I2(IntegralLimit[11]), .I3(n47835), .O(n47831));
    defparam i32317_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i31655_4_lut (.I0(n11_adj_3418), .I1(n9_adj_3420), .I2(n7_adj_3430), 
            .I3(n5_adj_3434), .O(n47169));
    defparam i31655_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_4_i13_rep_367_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n49860));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i13_rep_367_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32331_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n49860), 
            .I2(IntegralLimit[7]), .I3(n11_adj_3938), .O(n47845));
    defparam i32331_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32301_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n47845), .O(n47815));
    defparam i32301_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i31702_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n47216));
    defparam i31702_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_4_i35_rep_355_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n49848));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i35_rep_355_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_3941));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_4_i30_4_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[16]), .O(n30_adj_3942));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_4_i5_2_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(IntegralLimit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3943));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32341_4_lut (.I0(n9_adj_3939), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n5_adj_3943), .I3(IntegralLimit[3]), .O(n47855));
    defparam i32341_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i32337_4_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n11_adj_3938), 
            .I2(IntegralLimit[6]), .I3(n47855), .O(n47851));
    defparam i32337_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i31744_4_lut (.I0(n17_adj_3940), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n47851), .I3(IntegralLimit[7]), .O(n47258));
    defparam i31744_4_lut.LUT_INIT = 16'haeab;
    SB_LUT4 i32571_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[9]), 
            .I2(IntegralLimit[10]), .I3(n47258), .O(n48085));
    defparam i32571_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i32947_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[11]), 
            .I2(IntegralLimit[12]), .I3(n48085), .O(n48461));
    defparam i32947_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i32307_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n48461), .O(n47821));
    defparam i32307_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i32783_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n47821), .O(n48297));
    defparam i32783_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33018_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[17]), 
            .I2(IntegralLimit[18]), .I3(n48297), .O(n48532));
    defparam i33018_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33108_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[19]), 
            .I2(IntegralLimit[20]), .I3(n48532), .O(n48622));
    defparam i33108_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_4_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_3944));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31889_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(IntegralLimit[9]), .O(n47403));
    defparam i31889_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 LessThan_4_i24_4_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[21]), .O(n24_adj_3945));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i24_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i32663_3_lut (.I0(n6_adj_3944), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48177));   // verilog/motorControl.v(33[10:34])
    defparam i32663_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31671_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[12]), 
            .I2(IntegralLimit[21]), .I3(n47831), .O(n47185));
    defparam i31671_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_4_i45_rep_320_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n49813));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i45_rep_320_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32409_3_lut (.I0(n24_adj_3945), .I1(n8_adj_3933), .I2(n47403), 
            .I3(GND_net), .O(n47923));   // verilog/motorControl.v(33[10:34])
    defparam i32409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31938_4_lut (.I0(n48177), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[11]), .O(n47452));   // verilog/motorControl.v(33[10:34])
    defparam i31938_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_6_i4_4_lut (.I0(n63[0]), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3_adj_3437), .I3(\PID_CONTROLLER.integral [0]), .O(n4_adj_3946));   // verilog/motorControl.v(33[38:63])
    defparam LessThan_6_i4_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i32657_3_lut (.I0(n4_adj_3946), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n11_adj_3418), .I3(GND_net), .O(n48171));   // verilog/motorControl.v(33[38:63])
    defparam i32657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32658_3_lut (.I0(n48171), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n13_adj_3415), .I3(GND_net), .O(n48172));   // verilog/motorControl.v(33[38:63])
    defparam i32658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i8_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n17_adj_3411), .I3(GND_net), .O(n8_adj_3947));   // verilog/motorControl.v(33[38:63])
    defparam LessThan_6_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31641_2_lut (.I0(n17_adj_3411), .I1(n9_adj_3420), .I2(GND_net), 
            .I3(GND_net), .O(n47155));
    defparam i31641_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 LessThan_6_i6_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n7_adj_3430), .I3(GND_net), .O(n6_adj_3948));   // verilog/motorControl.v(33[38:63])
    defparam LessThan_6_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i16_3_lut (.I0(n8_adj_3947), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n44028), .I3(GND_net), .O(n16_adj_3949));   // verilog/motorControl.v(33[38:63])
    defparam LessThan_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31645_4_lut (.I0(n17_adj_3411), .I1(n15_adj_3414), .I2(n13_adj_3415), 
            .I3(n47169), .O(n47159));
    defparam i31645_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32739_4_lut (.I0(n16_adj_3949), .I1(n6_adj_3948), .I2(n44028), 
            .I3(n47155), .O(n48253));   // verilog/motorControl.v(33[38:63])
    defparam i32739_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i31948_3_lut (.I0(n48172), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n15_adj_3414), .I3(GND_net), .O(n47462));   // verilog/motorControl.v(33[38:63])
    defparam i31948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32995_4_lut (.I0(n47462), .I1(n48253), .I2(n44028), .I3(n47159), 
            .O(n48509));   // verilog/motorControl.v(33[38:63])
    defparam i32995_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_4_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(IntegralLimit[1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), .O(n4_adj_3950));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i32661_3_lut (.I0(n4_adj_3950), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48175));   // verilog/motorControl.v(33[10:34])
    defparam i32661_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31706_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n47815), .O(n47220));
    defparam i31706_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i32973_4_lut (.I0(n30_adj_3942), .I1(n10_adj_3941), .I2(n49848), 
            .I3(n47216), .O(n48487));   // verilog/motorControl.v(33[10:34])
    defparam i32973_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i31940_4_lut (.I0(n48175), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[14]), .O(n47454));   // verilog/motorControl.v(33[10:34])
    defparam i31940_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i33088_4_lut (.I0(n47454), .I1(n48487), .I2(n49848), .I3(n47220), 
            .O(n48602));   // verilog/motorControl.v(33[10:34])
    defparam i33088_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33089_3_lut (.I0(n48602), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48603));   // verilog/motorControl.v(33[10:34])
    defparam i33089_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32269_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(n48622), .O(n47783));
    defparam i32269_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i32873_4_lut (.I0(n47452), .I1(n47923), .I2(n49813), .I3(n47185), 
            .O(n48387));   // verilog/motorControl.v(33[10:34])
    defparam i32873_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31946_4_lut (.I0(n48603), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[19]), .O(n47460));   // verilog/motorControl.v(33[10:34])
    defparam i31946_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i32996_3_lut (.I0(n48509), .I1(n63[23]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48510));   // verilog/motorControl.v(33[38:63])
    defparam i32996_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32993_3_lut (.I0(n47460), .I1(n48387), .I2(n47783), .I3(GND_net), 
            .O(n48507));   // verilog/motorControl.v(33[10:34])
    defparam i32993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_1427 (.I0(n48507), .I1(n48510), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[23]), .O(n55_adj_3661));   // verilog/motorControl.v(33[10:63])
    defparam i8_4_lut_adj_1427.LUT_INIT = 16'h80c8;
    SB_LUT4 mult_12_i174_2_lut (.I0(\Kd[2] ), .I1(n67[21]), .I2(GND_net), 
            .I3(GND_net), .O(n258_adj_3660));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i239_2_lut (.I0(\Kd[3] ), .I1(n67[21]), .I2(GND_net), 
            .I3(GND_net), .O(n355_adj_3659));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i304_2_lut (.I0(\Kd[4] ), .I1(n67[21]), .I2(GND_net), 
            .I3(GND_net), .O(n452_adj_3658));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i369_2_lut (.I0(\Kd[5] ), .I1(n67[21]), .I2(GND_net), 
            .I3(GND_net), .O(n549_adj_3657));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i434_2_lut (.I0(\Kd[6] ), .I1(n67[21]), .I2(GND_net), 
            .I3(GND_net), .O(n646_adj_3656));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i499_2_lut (.I0(\Kd[7] ), .I1(n67[21]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_3655));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i111_2_lut (.I0(\Kd[1] ), .I1(n67[22]), .I2(GND_net), 
            .I3(GND_net), .O(n164_adj_3654));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i48_2_lut (.I0(\Kd[0] ), .I1(n67[23]), .I2(GND_net), 
            .I3(GND_net), .O(n71_adj_3653));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i48_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3652));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i176_2_lut (.I0(\Kd[2] ), .I1(n67[22]), .I2(GND_net), 
            .I3(GND_net), .O(n261_adj_3651));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i241_2_lut (.I0(\Kd[3] ), .I1(n67[22]), .I2(GND_net), 
            .I3(GND_net), .O(n358_adj_3650));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_3649));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i306_2_lut (.I0(\Kd[4] ), .I1(n67[22]), .I2(GND_net), 
            .I3(GND_net), .O(n455_adj_3647));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i371_2_lut (.I0(\Kd[5] ), .I1(n67[22]), .I2(GND_net), 
            .I3(GND_net), .O(n552_adj_3646));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i436_2_lut (.I0(\Kd[6] ), .I1(n67[22]), .I2(GND_net), 
            .I3(GND_net), .O(n649_adj_3645));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_3644));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i501_2_lut (.I0(\Kd[7] ), .I1(n67[22]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_3642));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3641));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3640));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i136_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n201_adj_3639));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i201_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n298_adj_3638));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i266_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n395_adj_3637));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i331_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n492_adj_3636));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n589_adj_3635));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i113_2_lut (.I0(\Kd[1] ), .I1(n67[23]), .I2(GND_net), 
            .I3(GND_net), .O(n167_adj_3634));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i50_2_lut (.I0(\Kd[0] ), .I1(n67[24]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_3633));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i50_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n686_adj_3632));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i117_2_lut (.I0(\Kd[1] ), .I1(n67[25]), .I2(GND_net), 
            .I3(GND_net), .O(n182_adj_3631));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i117_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i178_2_lut (.I0(\Kd[2] ), .I1(n67[23]), .I2(GND_net), 
            .I3(GND_net), .O(n264_adj_3630));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i182_2_lut (.I0(\Kd[2] ), .I1(n67[25]), .I2(GND_net), 
            .I3(GND_net), .O(n276_adj_3629));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i182_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i243_2_lut (.I0(\Kd[3] ), .I1(n67[23]), .I2(GND_net), 
            .I3(GND_net), .O(n361_adj_3628));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i308_2_lut (.I0(\Kd[4] ), .I1(n67[23]), .I2(GND_net), 
            .I3(GND_net), .O(n458_adj_3626));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i373_2_lut (.I0(\Kd[5] ), .I1(n67[23]), .I2(GND_net), 
            .I3(GND_net), .O(n555_adj_3623));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1428 (.I0(\Kd[2] ), .I1(\Kd[0] ), .I2(n67[25]), 
            .I3(\Kd[1] ), .O(n4_adj_3924));   // verilog/motorControl.v(36[26:45])
    defparam i2_4_lut_adj_1428.LUT_INIT = 16'ha080;
    SB_LUT4 mult_12_i247_2_lut (.I0(\Kd[3] ), .I1(n67[25]), .I2(GND_net), 
            .I3(GND_net), .O(n370_adj_3627));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22781_3_lut (.I0(n67[25]), .I1(n36328), .I2(n36343), .I3(GND_net), 
            .O(n10115[1]));   // verilog/motorControl.v(36[26:45])
    defparam i22781_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_12_i312_2_lut (.I0(\Kd[4] ), .I1(n67[25]), .I2(GND_net), 
            .I3(GND_net), .O(n464_adj_3624));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i379_2_lut (.I0(\Kd[5] ), .I1(n67[25]), .I2(GND_net), 
            .I3(GND_net), .O(n564));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i379_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i442_2_lut (.I0(\Kd[6] ), .I1(n67[25]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_3622));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i442_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1429 (.I0(n36328), .I1(n7_adj_3951), .I2(n8_adj_3931), 
            .I3(n8_adj_3932), .O(n44226));   // verilog/motorControl.v(36[26:45])
    defparam i5_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 mult_12_i438_2_lut (.I0(\Kd[6] ), .I1(n67[23]), .I2(GND_net), 
            .I3(GND_net), .O(n652_adj_3621));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i503_2_lut (.I0(\Kd[7] ), .I1(n67[23]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_3619));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i115_2_lut (.I0(\Kd[1] ), .I1(n67[24]), .I2(GND_net), 
            .I3(GND_net), .O(n170_adj_3618));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i52_2_lut (.I0(\Kd[0] ), .I1(n67[25]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_3617));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i52_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i180_2_lut (.I0(\Kd[2] ), .I1(n67[24]), .I2(GND_net), 
            .I3(GND_net), .O(n267));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i245_2_lut (.I0(\Kd[3] ), .I1(n67[24]), .I2(GND_net), 
            .I3(GND_net), .O(n364));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i310_2_lut (.I0(\Kd[4] ), .I1(n67[24]), .I2(GND_net), 
            .I3(GND_net), .O(n461_c));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3614));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i375_2_lut (.I0(\Kd[5] ), .I1(n67[24]), .I2(GND_net), 
            .I3(GND_net), .O(n558_adj_3613));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i199_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n295_adj_3612));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i199_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i264_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n392));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i264_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i440_2_lut (.I0(\Kd[6] ), .I1(n67[24]), .I2(GND_net), 
            .I3(GND_net), .O(n655));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i440_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i505_2_lut (.I0(\Kd[7] ), .I1(n67[24]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_3611));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i329_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n489));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i329_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n586));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n683));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15265_1_lut (.I0(pwm_count[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n28668));   // verilog/motorControl.v(99[18:29])
    defparam i15265_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i1_1_lut (.I0(pwm[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[0]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i2_1_lut (.I0(pwm[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[1]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i67_2_lut (.I0(\Kd[1] ), .I1(n67[0]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_3608));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i4_2_lut (.I0(\Kd[0] ), .I1(n67[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_3607));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i132_2_lut (.I0(\Kd[2] ), .I1(n67[0]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_3605));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i197_2_lut (.I0(\Kd[3] ), .I1(n67[0]), .I2(GND_net), 
            .I3(GND_net), .O(n292_adj_3604));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i262_2_lut (.I0(\Kd[4] ), .I1(n67[0]), .I2(GND_net), 
            .I3(GND_net), .O(n389_adj_3603));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i262_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i327_2_lut (.I0(\Kd[5] ), .I1(n67[0]), .I2(GND_net), 
            .I3(GND_net), .O(n486_adj_3601));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31804_2_lut_3_lut (.I0(hall3), .I1(hall1), .I2(n878), .I3(GND_net), 
            .O(n46593));   // verilog/motorControl.v(77[14] 98[8])
    defparam i31804_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 unary_minus_70_inv_0_i3_1_lut (.I0(pwm[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[2]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i4_1_lut (.I0(pwm[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[3]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i392_2_lut (.I0(\Kd[6] ), .I1(n67[0]), .I2(GND_net), 
            .I3(GND_net), .O(n583_adj_3598));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3660_2_lut_3_lut (.I0(hall1), .I1(hall2), .I2(PHASES_5__N_3039[1]), 
            .I3(GND_net), .O(n16802));   // verilog/motorControl.v(74[7] 76[10])
    defparam i3660_2_lut_3_lut.LUT_INIT = 16'h7474;
    SB_LUT4 mult_12_i457_2_lut (.I0(\Kd[7] ), .I1(n67[0]), .I2(GND_net), 
            .I3(GND_net), .O(n680_adj_3597));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i111_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i48_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n71));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i48_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i5_1_lut (.I0(pwm[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[4]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i176_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n261));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 PHASES_5__I_0_i2_4_lut_4_lut (.I0(n20375), .I1(hall3), .I2(hall1), 
            .I3(n17_adj_3482), .O(PHASES_5__N_2779[1]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i2_4_lut_4_lut.LUT_INIT = 16'h100c;
    SB_LUT4 i2_3_lut_4_lut_adj_1430 (.I0(hall1), .I1(hall2), .I2(n878), 
            .I3(PHASES_5__N_3039[1]), .O(n20375));   // verilog/motorControl.v(96[14] 98[8])
    defparam i2_3_lut_4_lut_adj_1430.LUT_INIT = 16'h7f4f;
    SB_LUT4 unary_minus_70_inv_0_i6_1_lut (.I0(pwm[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[5]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut (.I0(hall3), .I1(hall1), .I2(n17_adj_3482), 
            .I3(GND_net), .O(n42708));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 mult_10_i241_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n358));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i7_1_lut (.I0(pwm[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[6]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n455_adj_3588));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i8_1_lut (.I0(pwm[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[7]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i9_1_lut (.I0(pwm[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[8]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n552));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i10_1_lut (.I0(pwm[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n73[9]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i436_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n649));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i501_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3578));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i197_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n292));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i262_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n389));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i262_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i327_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n486));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i392_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n583));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n680));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i105_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n155));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i170_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n252));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i170_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i11_1_lut (.I0(pwm[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[10]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i91_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n134_adj_3564));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i91_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3563));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i235_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n349));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n446_adj_3559));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n543));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i156_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n231_adj_3558));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i95_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3557));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i46_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3556));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i430_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n640));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i430_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i221_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n328_adj_3553));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i144_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_3552));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i495_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i12_1_lut (.I0(pwm[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[11]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i286_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n425_adj_3549));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i71_2_lut (.I0(\Kd[1] ), .I1(n67[2]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i8_2_lut (.I0(\Kd[0] ), .I1(n67[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3548));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i136_2_lut (.I0(\Kd[2] ), .I1(n67[2]), .I2(GND_net), 
            .I3(GND_net), .O(n201));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i193_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i193_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n522_adj_3547));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i201_2_lut (.I0(\Kd[3] ), .I1(n67[2]), .I2(GND_net), 
            .I3(GND_net), .O(n298_adj_3545));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n619));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i266_2_lut (.I0(\Kd[4] ), .I1(n67[2]), .I2(GND_net), 
            .I3(GND_net), .O(n395));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i13_1_lut (.I0(pwm[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[12]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i242_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i242_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i481_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n716));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i331_2_lut (.I0(\Kd[5] ), .I1(n67[2]), .I2(GND_net), 
            .I3(GND_net), .O(n492));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i396_2_lut (.I0(\Kd[6] ), .I1(n67[2]), .I2(GND_net), 
            .I3(GND_net), .O(n589_adj_3541));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i103_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n152));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i40_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n59));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i461_2_lut (.I0(\Kd[7] ), .I1(n67[2]), .I2(GND_net), 
            .I3(GND_net), .O(n686));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i168_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n249));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i168_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i291_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i291_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31796_4_lut_4_lut (.I0(hall1), .I1(hall2), .I2(n878), .I3(hall3), 
            .O(n46611));
    defparam i31796_4_lut_4_lut.LUT_INIT = 16'h8010;
    SB_LUT4 i10292_2_lut_4_lut (.I0(PHASES_5__N_3039[4]), .I1(hall3), .I2(n19954), 
            .I3(n934), .O(PHASES_5__N_3039[2]));   // verilog/motorControl.v(74[7] 76[10])
    defparam i10292_2_lut_4_lut.LUT_INIT = 16'hff47;
    SB_LUT4 unary_minus_70_inv_0_i14_1_lut (.I0(pwm[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[13]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i233_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n346));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i15_1_lut (.I0(pwm[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[14]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n443_adj_3536));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i340_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i340_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n540));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i428_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n637));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i389_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i389_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i493_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i493_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i16_1_lut (.I0(pwm[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[15]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31801_2_lut_4_lut (.I0(PHASES_5__N_3039[4]), .I1(hall3), .I2(PHASES_5__N_3039[3]), 
            .I3(n878), .O(n46609));
    defparam i31801_2_lut_4_lut.LUT_INIT = 16'h0700;
    SB_LUT4 unary_minus_70_inv_0_i17_1_lut (.I0(pwm[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[16]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31794_2_lut_4_lut (.I0(hall2), .I1(hall1), .I2(hall3), .I3(n878), 
            .O(n46608));
    defparam i31794_2_lut_4_lut.LUT_INIT = 16'hd500;
    SB_LUT4 mult_10_i101_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n149));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i18_1_lut (.I0(pwm[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[17]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i166_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n246));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i19_1_lut (.I0(pwm[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[18]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i231_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n343));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i20_1_lut (.I0(pwm[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[19]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i21_1_lut (.I0(pwm[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[20]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i73_2_lut (.I0(\Kd[1] ), .I1(n67[3]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i10_2_lut (.I0(\Kd[0] ), .I1(n67[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_3525));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n440));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n537));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i22_1_lut (.I0(pwm[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[21]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i138_2_lut (.I0(\Kd[2] ), .I1(n67[3]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i203_2_lut (.I0(\Kd[3] ), .I1(n67[3]), .I2(GND_net), 
            .I3(GND_net), .O(n301_adj_3522));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i426_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n634));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i426_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i268_2_lut (.I0(\Kd[4] ), .I1(n67[3]), .I2(GND_net), 
            .I3(GND_net), .O(n398));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i23_1_lut (.I0(pwm[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n73[22]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i24_1_lut (.I0(pwm[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(PHASES_5__N_3046));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n131_adj_3518));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_3517));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i1_1_lut (.I0(\PID_CONTROLLER.err[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[0]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i491_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i2_1_lut (.I0(\PID_CONTROLLER.err[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[1]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i154_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n228_adj_3514));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i154_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i333_2_lut (.I0(\Kd[5] ), .I1(n67[3]), .I2(GND_net), 
            .I3(GND_net), .O(n495));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i333_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i3_1_lut (.I0(\PID_CONTROLLER.err[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[2]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i219_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n325_adj_3512));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i398_2_lut (.I0(\Kd[6] ), .I1(n67[3]), .I2(GND_net), 
            .I3(GND_net), .O(n592_adj_3511));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i4_1_lut (.I0(\PID_CONTROLLER.err[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[3]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i284_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n422_adj_3509));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i284_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i5_1_lut (.I0(\PID_CONTROLLER.err[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[4]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i463_2_lut (.I0(\Kd[7] ), .I1(n67[3]), .I2(GND_net), 
            .I3(GND_net), .O(n689));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n519_adj_3507));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i6_1_lut (.I0(\PID_CONTROLLER.err[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[5]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n616_adj_3505));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i7_1_lut (.I0(\PID_CONTROLLER.err[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[6]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i479_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n713_adj_3503));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i8_1_lut (.I0(\PID_CONTROLLER.err[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[7]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i9_1_lut (.I0(\PID_CONTROLLER.err[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[8]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31502_2_lut_4_lut (.I0(\PID_CONTROLLER.result [8]), .I1(pwm_23__N_2951[8]), 
            .I2(\pwm_23__N_2951[4] ), .I3(\PID_CONTROLLER.result[4] ), .O(n47016));
    defparam i31502_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut (.I0(\PID_CONTROLLER.result [28]), .I1(\PID_CONTROLLER.result [30]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(n56_adj_3871), .O(n42629));   // verilog/motorControl.v(38[12:27])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_12_i75_2_lut (.I0(\Kd[1] ), .I1(n67[4]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i12_2_lut (.I0(\Kd[0] ), .I1(n67[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3500));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i10_1_lut (.I0(\PID_CONTROLLER.err[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[9]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i140_2_lut (.I0(\Kd[2] ), .I1(n67[4]), .I2(GND_net), 
            .I3(GND_net), .O(n207));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i205_2_lut (.I0(\Kd[3] ), .I1(n67[4]), .I2(GND_net), 
            .I3(GND_net), .O(n304_adj_3498));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i205_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i270_2_lut (.I0(\Kd[4] ), .I1(n67[4]), .I2(GND_net), 
            .I3(GND_net), .O(n401));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i11_1_lut (.I0(\PID_CONTROLLER.err[10] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[10]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i505_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i12_1_lut (.I0(\PID_CONTROLLER.err[11] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[11]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i335_2_lut (.I0(\Kd[5] ), .I1(n67[4]), .I2(GND_net), 
            .I3(GND_net), .O(n498));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i335_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i400_2_lut (.I0(\Kd[6] ), .I1(n67[4]), .I2(GND_net), 
            .I3(GND_net), .O(n595_adj_3495));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i13_1_lut (.I0(\PID_CONTROLLER.err[12] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[12]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i465_2_lut (.I0(\Kd[7] ), .I1(n67[4]), .I2(GND_net), 
            .I3(GND_net), .O(n692));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i99_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n146));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i99_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3492));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i4_4_lut_4_lut (.I0(\PWMLimit[0] ), .I1(\PID_CONTROLLER.result [1]), 
            .I2(\PWMLimit[1] ), .I3(\PID_CONTROLLER.result [0]), .O(n4_adj_3860));   // verilog/motorControl.v(38[12:27])
    defparam LessThan_20_i4_4_lut_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_10_i164_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n243));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i164_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut  (.I0(\PID_CONTROLLER.result[4] ), 
            .I1(\PID_CONTROLLER.result [8]), .I2(\deadband[8] ), .I3(GND_net), 
            .O(n8_adj_3852));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [2]), 
            .I1(\PID_CONTROLLER.result [3]), .I2(\deadband[3] ), .I3(GND_net), 
            .O(n6_adj_3850));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut  (.I0(\PID_CONTROLLER.result[5] ), 
            .I1(\PID_CONTROLLER.result [6]), .I2(\deadband[6] ), .I3(GND_net), 
            .O(n10_adj_3854));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_11_inv_0_i14_1_lut (.I0(\PID_CONTROLLER.err[13] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[13]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i229_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n340));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i15_1_lut (.I0(\PID_CONTROLLER.err[14] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[14]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i16_1_lut (.I0(\PID_CONTROLLER.err[15] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[15]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i294_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n437));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i17_1_lut (.I0(\PID_CONTROLLER.err[16] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[16]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i18_1_lut (.I0(\PID_CONTROLLER.err[17] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[17]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n534));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n631));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i19_1_lut (.I0(\PID_CONTROLLER.err[18] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[18]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i489_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n728));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i20_1_lut (.I0(\PID_CONTROLLER.err[19] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[19]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i21_1_lut (.I0(\PID_CONTROLLER.err[20] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[20]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i22_1_lut (.I0(\PID_CONTROLLER.err[21] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[21]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i77_2_lut (.I0(\Kd[1] ), .I1(n67[5]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i14_2_lut (.I0(\Kd[0] ), .I1(n67[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_3480));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i142_2_lut (.I0(\Kd[2] ), .I1(n67[5]), .I2(GND_net), 
            .I3(GND_net), .O(n210));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i207_2_lut (.I0(\Kd[3] ), .I1(n67[5]), .I2(GND_net), 
            .I3(GND_net), .O(n307_adj_3479));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22506_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(GND_net), .O(n16641[0]));   // verilog/motorControl.v(36[17:23])
    defparam i22506_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 mult_12_i272_2_lut (.I0(\Kd[4] ), .I1(n67[5]), .I2(GND_net), 
            .I3(GND_net), .O(n404));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i23_1_lut (.I0(\PID_CONTROLLER.err[22] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[22]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22507_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n38421));   // verilog/motorControl.v(36[17:23])
    defparam i22507_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mult_12_i337_2_lut (.I0(\Kd[5] ), .I1(n67[5]), .I2(GND_net), 
            .I3(GND_net), .O(n501));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i402_2_lut (.I0(\Kd[6] ), .I1(n67[5]), .I2(GND_net), 
            .I3(GND_net), .O(n598_adj_3477));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i467_2_lut (.I0(\Kd[7] ), .I1(n67[5]), .I2(GND_net), 
            .I3(GND_net), .O(n695));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i24_1_lut (.I0(\PID_CONTROLLER.err[23] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[23]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i115_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n182));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15554_1_lut (.I0(\PID_CONTROLLER.result [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28960));   // verilog/motorControl.v(31[14] 52[8])
    defparam i15554_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i1_1_lut (.I0(\deadband[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[0]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i2_1_lut (.I0(\deadband[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[1]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i3_1_lut (.I0(\deadband[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n69[2]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i286_2_lut (.I0(\Kd[4] ), .I1(n67[12]), .I2(GND_net), 
            .I3(GND_net), .O(n425));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n558));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i180_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n276));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i245_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n370_adj_3471));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22508_3_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n36197), .I2(n38421), 
            .I3(GND_net), .O(n16654[1]));   // verilog/motorControl.v(36[17:23])
    defparam i22508_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n464));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i442_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i442_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1431 (.I0(n36197), .I1(n7_adj_3929), .I2(n8_adj_3926), 
            .I3(n8_adj_3927), .O(n43817));   // verilog/motorControl.v(36[17:23])
    defparam i5_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i97_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n143));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i97_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i162_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n240));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i227_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n337));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i292_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n434));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n531));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n628));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i487_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n725));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_556_i4_4_lut_4_lut (.I0(pwm_count[0]), .I1(pwm[0]), 
            .I2(\pwm_count[1] ), .I3(pwm[1]), .O(n4));   // verilog/motorControl.v(99[18:29])
    defparam LessThan_556_i4_4_lut_4_lut.LUT_INIT = 16'h4f04;
    SB_LUT4 i22813_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(\Kd[2] ), 
            .I3(GND_net), .O(n36343));   // verilog/motorControl.v(36[26:45])
    defparam i22813_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i22812_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(n67[25]), 
            .I3(GND_net), .O(n10115[0]));   // verilog/motorControl.v(36[26:45])
    defparam i22812_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i1_3_lut_4_lut_adj_1432 (.I0(n370_adj_3627), .I1(n4_adj_3924), 
            .I2(n36343), .I3(n67[25]), .O(n7_adj_3951));   // verilog/motorControl.v(36[26:45])
    defparam i1_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6966;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1433 (.I0(hall1), .I1(hall3), .I2(n880), 
            .I3(n20375), .O(n4_adj_3914));
    defparam i1_2_lut_3_lut_4_lut_adj_1433.LUT_INIT = 16'hffe2;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=47, LSE_LCOL=12, LSE_RCOL=39, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, n22513, GND_net, \Kd[7] , gearBoxRatio, rx_data, 
            IntegralLimit, n24320, \data_in[0] , n24319, n24318, \deadband[9] , 
            \deadband[8] , \deadband[7] , \deadband[6] , \deadband[5] , 
            \deadband[4] , \deadband[3] , \deadband[2] , n24482, VCC_net, 
            byte_transmit_counter, \deadband[1] , n24478, setpoint, 
            n24477, n24476, n24475, n24474, n24473, n24472, n24471, 
            n24470, n24469, n24468, n24467, n24466, n24465, n24464, 
            n24463, n24462, n24461, n24460, n24459, n24458, n24457, 
            n24456, n23891, n24306, \data_in[1] , n24305, \data_in[2] , 
            n24304, n24303, n24302, n24301, n24300, n24299, n24298, 
            n24297, \data_in[3] , n24296, n24295, n24294, n24293, 
            n24292, n24291, n24290, n24289, \data_out_frame[0][2] , 
            n24288, \data_out_frame[0][3] , n24287, \data_out_frame[0][4] , 
            n24284, \data_out_frame[5][2] , n24317, n24316, n24315, 
            n24314, rx_data_ready, n24313, n24312, \Kp[1] , \Kp[2] , 
            \FRAME_MATCHER.state[0] , n22525, n24158, \data_out_frame[22] , 
            \Kp[3] , \Kp[4] , \FRAME_MATCHER.state[2] , n22498, encoder0_position, 
            displacement, \Kp[5] , \FRAME_MATCHER.state[3] , n22528, 
            n23894, pwm, encoder1_position, control_mode, n23907, 
            n3840, n23904, n23901, n24311, \Kp[6] , n23898, n41946, 
            n23895, n23892, n23889, n2241, \PWMLimit[1] , \PWMLimit[2] , 
            \PWMLimit[3] , \PWMLimit[4] , \PWMLimit[5] , \PWMLimit[6] , 
            \PWMLimit[7] , \PWMLimit[8] , \PWMLimit[9] , n49493, \Kp[7] , 
            \Ki[1] , \Ki[2] , \Ki[3] , n24310, n24309, \Ki[4] , 
            n5025, n5023, n23616, n24308, n3362, n24307, \Ki[5] , 
            n23897, n23900, n23903, n23906, n23909, \Ki[6] , \Ki[7] , 
            \Kd[1] , \Kd[2] , \Kd[3] , \Kd[4] , \Kd[5] , \Kd[6] , 
            \deadband[0] , n23828, n42006, \PWMLimit[0] , n23808, 
            \Kd[0] , \Ki[0] , \Kp[0] , n3800, n3801, n3802, n3803, 
            n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, 
            n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, 
            n3820, n3821, n3823, n3822, n44107, n28694, n122, 
            n2854, n63, n5, n50013, n39599, \FRAME_MATCHER.state_31__N_1860[1] , 
            n43447, n22512, n43773, n2119, n3758, n737, n20156, 
            n3, n22511, n5_adj_3, n23847, n23850, n23853, n23856, 
            n23859, n23862, n23865, n23868, n23872, r_Bit_Index, 
            n23875, n23845, n23848, n23851, n23915, n23918, n23854, 
            n23857, n23860, n23863, n23866, n23913, tx_o, n23655, 
            n23785, n4038, n23914, tx_enable, n23878, r_Bit_Index_adj_9, 
            n23881, n24453, n29023, \r_SM_Main[1] , r_Rx_Data, LED_c, 
            n24391, \r_SM_Main[2] , n23888, n23887, n23886, n23885, 
            n23884, n23883, n23882, n23817, n46591, n22534, n4, 
            n28989, n28517, n4_adj_7, n4_adj_8, n23649, n23783, 
            n4016, n22539, n1, n46590) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    output n22513;
    input GND_net;
    output \Kd[7] ;
    output [23:0]gearBoxRatio;
    output [7:0]rx_data;
    output [23:0]IntegralLimit;
    input n24320;
    output [7:0]\data_in[0] ;
    input n24319;
    input n24318;
    output \deadband[9] ;
    output \deadband[8] ;
    output \deadband[7] ;
    output \deadband[6] ;
    output \deadband[5] ;
    output \deadband[4] ;
    output \deadband[3] ;
    output \deadband[2] ;
    input n24482;
    input VCC_net;
    output [7:0]byte_transmit_counter;
    output \deadband[1] ;
    input n24478;
    output [23:0]setpoint;
    input n24477;
    input n24476;
    input n24475;
    input n24474;
    input n24473;
    input n24472;
    input n24471;
    input n24470;
    input n24469;
    input n24468;
    input n24467;
    input n24466;
    input n24465;
    input n24464;
    input n24463;
    input n24462;
    input n24461;
    input n24460;
    input n24459;
    input n24458;
    input n24457;
    input n24456;
    input n23891;
    input n24306;
    output [7:0]\data_in[1] ;
    input n24305;
    output [7:0]\data_in[2] ;
    input n24304;
    input n24303;
    input n24302;
    input n24301;
    input n24300;
    input n24299;
    input n24298;
    input n24297;
    output [7:0]\data_in[3] ;
    input n24296;
    input n24295;
    input n24294;
    input n24293;
    input n24292;
    input n24291;
    input n24290;
    input n24289;
    output \data_out_frame[0][2] ;
    input n24288;
    output \data_out_frame[0][3] ;
    input n24287;
    output \data_out_frame[0][4] ;
    input n24284;
    output \data_out_frame[5][2] ;
    input n24317;
    input n24316;
    input n24315;
    input n24314;
    output rx_data_ready;
    input n24313;
    input n24312;
    output \Kp[1] ;
    output \Kp[2] ;
    output \FRAME_MATCHER.state[0] ;
    output n22525;
    input n24158;
    output [7:0]\data_out_frame[22] ;
    output \Kp[3] ;
    output \Kp[4] ;
    output \FRAME_MATCHER.state[2] ;
    output n22498;
    input [23:0]encoder0_position;
    input [23:0]displacement;
    output \Kp[5] ;
    output \FRAME_MATCHER.state[3] ;
    output n22528;
    input n23894;
    input [23:0]pwm;
    input [23:0]encoder1_position;
    output [7:0]control_mode;
    output n23907;
    output n3840;
    output n23904;
    output n23901;
    input n24311;
    output \Kp[6] ;
    output n23898;
    input n41946;
    output n23895;
    output n23892;
    output n23889;
    output n2241;
    output \PWMLimit[1] ;
    output \PWMLimit[2] ;
    output \PWMLimit[3] ;
    output \PWMLimit[4] ;
    output \PWMLimit[5] ;
    output \PWMLimit[6] ;
    output \PWMLimit[7] ;
    output \PWMLimit[8] ;
    output \PWMLimit[9] ;
    input n49493;
    output \Kp[7] ;
    output \Ki[1] ;
    output \Ki[2] ;
    output \Ki[3] ;
    input n24310;
    input n24309;
    output \Ki[4] ;
    output n5025;
    output n5023;
    output n23616;
    input n24308;
    output n3362;
    input n24307;
    output \Ki[5] ;
    input n23897;
    input n23900;
    input n23903;
    input n23906;
    input n23909;
    output \Ki[6] ;
    output \Ki[7] ;
    output \Kd[1] ;
    output \Kd[2] ;
    output \Kd[3] ;
    output \Kd[4] ;
    output \Kd[5] ;
    output \Kd[6] ;
    output \deadband[0] ;
    input n23828;
    input n42006;
    output \PWMLimit[0] ;
    input n23808;
    output \Kd[0] ;
    output \Ki[0] ;
    output \Kp[0] ;
    output n3800;
    output n3801;
    output n3802;
    output n3803;
    output n3804;
    output n3805;
    output n3806;
    output n3807;
    output n3808;
    output n3809;
    output n3810;
    output n3811;
    output n3812;
    output n3813;
    output n3814;
    output n3815;
    output n3816;
    output n3817;
    output n3818;
    output n3819;
    output n3820;
    output n3821;
    output n3823;
    output n3822;
    output n44107;
    output n28694;
    output n122;
    output n2854;
    output n63;
    output n5;
    output n50013;
    output n39599;
    output \FRAME_MATCHER.state_31__N_1860[1] ;
    output n43447;
    output n22512;
    input n43773;
    output n2119;
    output n3758;
    output n737;
    output n20156;
    output n3;
    output n22511;
    output n5_adj_3;
    input n23847;
    input n23850;
    input n23853;
    input n23856;
    input n23859;
    input n23862;
    input n23865;
    input n23868;
    input n23872;
    output [2:0]r_Bit_Index;
    input n23875;
    output n23845;
    output n23848;
    output n23851;
    input n23915;
    input n23918;
    output n23854;
    output n23857;
    output n23860;
    output n23863;
    output n23866;
    output n23913;
    output tx_o;
    output n23655;
    output n23785;
    output n4038;
    output n23914;
    output tx_enable;
    input n23878;
    output [2:0]r_Bit_Index_adj_9;
    input n23881;
    input n24453;
    input n29023;
    output \r_SM_Main[1] ;
    output r_Rx_Data;
    input LED_c;
    input n24391;
    output \r_SM_Main[2] ;
    input n23888;
    input n23887;
    input n23886;
    input n23885;
    input n23884;
    input n23883;
    input n23882;
    input n23817;
    output n46591;
    output n22534;
    output n4;
    output n28989;
    output n28517;
    output n4_adj_7;
    output n4_adj_8;
    output n23649;
    output n23783;
    output n4016;
    output n22539;
    output n1;
    output n46590;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n24271;
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(94[12:26])
    
    wire n24270;
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(94[12:26])
    
    wire n28588, n22520;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(112[11:12])
    
    wire n3_c, n24269, n24268, n3_adj_3110, n3_adj_3111;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(93[12:25])
    
    wire n23449, n23233, n43133, n3_adj_3112, n36460, n36461, n24267, 
        n3_adj_3113, n24344, n24343, n24342, n24341, n3_adj_3114, 
        n24266, n24340, n24339, n3_adj_3115, n24265, n3_adj_3116, 
        n3_adj_3117, n3_adj_3118, n3_adj_3119, n3_adj_3120, n23229, 
        n23168, n43102, n3_adj_3121, n3_adj_3122, n3_adj_3123, n43885;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(93[12:25])
    
    wire n14, n3_adj_3124, n8, n42698;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(93[12:25])
    
    wire n24023, n24338, n24024, n24025, n24026, n24264, n24337, 
        n24027, n24028, n24029, n23479, n14_adj_3125, n24336, n24335, 
        n24377, n2, n36459, n1508, n24030, n8_adj_3126, n24015, 
        n24016, n24334, n24333, n24332, n24331, n24263, n36472, 
        n36473, n24330, n24329, n24328, n24327, n24326, n24325, 
        n24324, n24323, n24017, n24322, n24321, n24018, n2_adj_3127, 
        n36471, n24262;
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(94[12:26])
    
    wire n24261, n24019, n24020, n2_adj_3128, n36470, n24021, n24022, 
        n2_adj_3129, n36458, n2_adj_3130, n36469;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(93[12:25])
    
    wire Kp_23__N_838, n43148, n23038;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(93[12:25])
    
    wire n39055, n8_adj_3131, n24007, n24490, n24008, n24489, n24488, 
        n24487, n24486, n24485, n24484, n24483, n24009, n24479;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(99[12:33])
    
    wire n24260, n24259, n24258, n24257, n24256, n24255, n24254;
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(94[12:26])
    
    wire n24253, n24252, n24251, n24250, n24249, n24248, n24247, 
        n24246;
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(94[12:26])
    
    wire n24286;
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(94[12:26])
    
    wire n24285, n24283, n24282, n24376, n24375, n24374, n24373, 
        n24372, n24371, n24370, n24245, n24244, n24243, n24242, 
        n24241, n24281, n24280, n24279, n24278, n24277, n24276, 
        n24240, n24239, n24275, n24010, n24274, n24238;
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(94[12:26])
    
    wire n24369, n24011, n24237, n24012, n24013, n24014, n8_adj_3132, 
        n23999, n24000, n24001, n24002, n24236, n24235, n24234, 
        n24233, n24003, n24232, n24231, n24230;
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(94[12:26])
    
    wire n24229, n24228, n24227, n24226, n24225, n24224, n24223, 
        n24222;
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(94[12:26])
    
    wire n24221, n24220, n24219, n24004, n24218, n24217, n24216, 
        n24215, n24005, n24214;
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(94[12:26])
    
    wire n24213, n24212, n24211, \FRAME_MATCHER.rx_data_ready_prev , 
        n24210, n24006, n24209, n24273, n24368, n8_adj_3133;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(93[12:25])
    
    wire n23991, n24208, n24207, n23992, n24206;
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(94[12:26])
    
    wire n24205, n24204, n24203, n24379, n24202, n24367, n23993, 
        n23994, n24366, n24365, n23995, n24364, Kp_23__N_785, n43313, 
        n23513, n23996, n24363, n23997, n43105, Kp_23__N_994, n24201, 
        n24200, n24199, n24198;
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(94[12:26])
    
    wire n24197, n24196, n24195, n24194, n24193, n24192, n24191, 
        n24190;
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(94[12:26])
    
    wire n24189, n24188, n39460, Kp_23__N_945, n39629, n23026, n23998, 
        n24187, n24186;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(109[11:16])
    
    wire n22524, n24185, n43142, n43139, n8_adj_3134, n24184, n8_adj_3135;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(93[12:25])
    
    wire n23983, n24183, n24182;
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(94[12:26])
    
    wire n24181, n23462, n6, n24180, n23984, n24179, n23985, n24178, 
        n24177, n24176, n24175, n24174;
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(94[12:26])
    
    wire n24378, n24173, n24172, n24171, n24170, n24169, n24168, 
        n24167, n24166;
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(94[12:26])
    
    wire n24165, n24164, n23986, n24163, n24162, n24161, n24160, 
        n24159, n22942, n10, n43172, n23987, n24157;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(93[12:25])
    
    wire n24156, n24155, n23988, n23989, n24154, n24153, n24152, 
        n24151, n24150;
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(93[12:25])
    
    wire n23990, n24149, n24148, n24147, n24146, n24145, n24362, 
        n24144, n24361, n24143, n24142;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(93[12:25])
    
    wire n24141, n24140, n24139, n24138, n24137, n24136, n24135, 
        n24134;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(93[12:25])
    
    wire n24133, n24132, n24131, n24130, n24129, n24128, n24127, 
        n24126;
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(93[12:25])
    
    wire n24125, n24124, n24123, n24122, n24121, n24120, n24119, 
        n24118;
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(93[12:25])
    
    wire n24117, n24116, n24115, n24114, n24113, n24112, n24111, 
        n24110;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(93[12:25])
    
    wire n2_adj_3136, n36468, n24109, n24360, n2_adj_3137, n36457, 
        n24108, n24387, n24107, n2_adj_3138, n36467;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(94[12:26])
    
    wire n19, n46842, n5_c;
    wire [7:0]\data_out_frame[22]_c ;   // verilog/coms.v(94[12:26])
    
    wire n44683, n49387, n44684, n44661, n24106, n24105, n44663, 
        n49471, n49477, n44662, n24104, n24103, n43193, n24102;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(93[12:25])
    
    wire n24101, n24100, n24099, n24098, n2_adj_3139, n36466, n24097, 
        n24096, n24095, n24094, n24093, n24092, n24091, n24090, 
        n24089, n24088, n42743, n39501, n42612, n24087, n42782, 
        n43238, n43030, n43310, n43231, n43077, n2_adj_3140, n36465, 
        n23017, Kp_23__N_776, n10_adj_3141, n39257, n43017, n24086;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(93[12:25])
    
    wire n43585, n43071, n43283, n43099, n10_adj_3142, n22891, n23266, 
        n23467, n43136, Kp_23__N_192, n24085, n10_adj_3143, n43228, 
        n43130, n21140, n14_adj_3144, n43225, n42904, n24084, n42995, 
        n24083, n43234, n43064, n2_adj_3145, n36456, n43011, n15, 
        n24082, n23208, n24386, n2_adj_3146, n36464, n39029, n43068, 
        n42969;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(93[12:25])
    
    wire n23018, n24272, n43295, n43322, n43005, n22801, n43059, 
        n43184, n43298, n15_adj_3147, n43084, n14_adj_3148, n44327, 
        n44318, n19_adj_3149, n46624, n49480, n17, n16, n49483, 
        n49474, n49468, n49462, n49465, n49456, n49459, n22682, 
        n43834, n22885;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(93[12:25])
    
    wire n6_adj_3150;
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(93[12:25])
    
    wire n42958, n42999, n10_adj_3151, n43221, n22858, n43056, n7, 
        n56, n42913, n55, n63_c, n43053, n43074, n42925, n60, 
        n42765, n22770, n58, n43262, n59, n43244, n43050, n57, 
        n62, n68, n42907, Kp_23__N_319, n61, n69, n43253, n43274, 
        n43181, n12, n43008, n15_adj_3152, n42919, n43026, n43090, 
        n12_adj_3153, n43241, n42901, n43196, n8_adj_3154, n42951, 
        n23470, n24385, n36492, Kp_23__N_458, n22826, n10_adj_3155, 
        n43271, n36491, n36490, n43042, n24081, n24080, n49450, 
        n24079, n49453, n24078, n24077, n49444, n24076, n49447, 
        n24075, n24074, n49438, n24073, n49441, n24072, n24071, 
        n49432, n24070, n49435, n24069, n24068, n49426, n24067, 
        n49429, n24066, n24065, n49420, n24064, n49423, n24063, 
        n24062, n49414, n24061, n48097, n24060, n24059, n49408, 
        n24058, n44739, n24057, n24056, n49402, n24055, n42840, 
        n22750, n12_adj_3156, n49405, n24054, n22815, n22781, n10_adj_3157, 
        n43316, n6_adj_3158, n22853, n42829, n23347, n23032, n10_adj_3159, 
        n10_adj_3160, n14_adj_3161, n24053, n24052, n24051, n24384, 
        n24359, n12_adj_3162, n24383, n7_adj_3163, n8_adj_3164, n36489, 
        n43256, n42755, n12_adj_3165, n43319, n39692, n22977, Kp_23__N_515, 
        n12_adj_3166, n42088, n42004, n42084, n41998, n42200, n41892, 
        n7_adj_3167, n8_adj_3168, n7_adj_3169, n28539, n42136, n28932, 
        n7_adj_3170, n8_adj_3171, n7_adj_3172, n8_adj_3173, n42124, 
        n41966, n42122, n42008, n7_adj_3174, n8_adj_3175, n42120, 
        n42010, n28495, n8_adj_3176, n42118, n42012, n7_adj_3177, 
        n8_adj_3178, n42116, n42014, n42114, n42016, n42112, n42018, 
        n42110, n42020, n42108, n42022, n42106, n42024, n42104, 
        n42026, n42102, n42028, n42100, n42030, n42044, n28920, 
        n28493, n28918, n42098, n41958, n41956, n42198, n49489, 
        n24050, n43081, n38953, n39049, n24049, n24048, n24047, 
        n24046, n24045, n24044, n24043, n24042, n24041, n24040, 
        n24039, n24038, n44064, n23610, n42769, n39661, n16_adj_3179, 
        n43033, n10_adj_3180, n14_adj_3181, n42984, n42924, n23309, 
        n43286, n23113, n6_adj_3182, n39672, n22958, n42897, n43063, 
        n23311, n43849, n44248, n44212, n44323, n43950, n43632, 
        n44218, n44444, n24037, n42849, n43259, n6_adj_3183, n42877, 
        n43162, n39331, n39675, n8_adj_3184, n43247, n23528, n4_c, 
        n24036, n36488, n42821, n6_adj_3185, n5_adj_3186, n39619, 
        n43014, n22979, n43054, n42832, n42817, n6_adj_3187, Kp_23__N_290, 
        n43145, n21084, n18, Kp_23__N_325, n20, n42772, n19_adj_3188, 
        n43117, n38906, n2_adj_3189, n23446, n5_adj_3190, n23164, 
        n12_adj_3191, n4_adj_3192, n10_adj_3193, n23519, n6_adj_3194, 
        n6_adj_3195, n39648, n14_adj_3196, n14_adj_3197, n13, n13_adj_3198, 
        n28473, n8_adj_3199, n44463, n10_adj_3200, n43842, n8_adj_3201, 
        n10_adj_3202, n2_adj_3203, n2_adj_3204, n2_adj_3205, n2_adj_3206, 
        n2_adj_3207, n2_adj_3208, n2_adj_3209, n2_adj_3210, n2_adj_3211, 
        n2_adj_3212, n2_adj_3213, n2_adj_3214, n2_adj_3215, n3_adj_3216, 
        n3_adj_3217, n3_adj_3218, n3_adj_3219, n3_adj_3220, n3_adj_3221, 
        n2_adj_3222, n3_adj_3223, n2_adj_3224, n3_adj_3225, n2_adj_3226, 
        n3_adj_3227, n2_adj_3228, n3_adj_3229, n3_adj_3230, n3_adj_3231, 
        n3_adj_3232, n3_adj_3233, n2_adj_3234, n3_adj_3235, n24035, 
        n43618, n10_adj_3236, n24034, n24033, n24032, n24031, n36487, 
        n36455, n43891, n49396, n44596, n36463, n36486, n10_adj_3237, 
        n11, tx_transmit_N_2639, n9, n49513, n12_adj_3238, n12_adj_3239, 
        n49399, n36485, n6_adj_3240, n43615, n36484, n8_adj_3241, 
        n44547, n36483, n43841, n44167, n42902, n13_adj_3242, n36482, 
        n44377, n12_adj_3243, n16_adj_3244, n43617, n31, n28496, 
        n36481, n23982, n23981, n23980, n23979, n23978, n23977, 
        n23976, n23975, n23974, n23973, n23972, n23971, n23970, 
        n28310, n23968, n23967, n36480, n2_adj_3245, n161, n36462, 
        n36479, n36478, n36477, n24358, n24357, n24356, n24355, 
        n49384, n24354, n28895;
    wire [31:0]\FRAME_MATCHER.state_31__N_1924 ;
    
    wire n36476, n24353, n46678;
    wire [2:0]r_SM_Main_2__N_2747;
    
    wire n43341, n24352, n36475, n24351, n24350, n24349, n24382, 
        n14_adj_3246, n49378, n49381, n36474, n13_adj_3247, n6_adj_3248, 
        n12_adj_3249, n14_adj_3250, n15_adj_3251, n29039, n22492, 
        n49497, n4_adj_3252, n24348, n24347, n24346, n24345, n23829, 
        n3_adj_3253, n24381, n24380, n23811, n23810, n23809, n23807, 
        n23806, n23805, n23804, n23803, n28475, n44681, n44680;
    wire [7:0]tx_data;   // verilog/coms.v(102[13:20])
    
    wire n44678, n44677, n44675, n44674, n44672, n44671, n49372, 
        n44666, n44665, n44669, n44668, n44689, n44688, n49375, 
        n5_adj_3254, n49366, n49369, n31_adj_3255, n49360, n19960, 
        n15_adj_3256, n28, n26, n27, n25, n20014, n6_adj_3257, 
        n29029, n29035, n4_adj_3258, n19_adj_3259, n47008, n5_adj_3260, 
        n44659, n49363, n44660, n46420, n44679, n19_adj_3261, n47001, 
        n5_adj_3262, n44656, n49357, n44657, n44676, n49333, n19_adj_3263, 
        n46994, n5_adj_3264, n44653, n49351, n44654, n44673, n49339, 
        n19_adj_3265, n44650, n49345, n44651, n46586, n6_adj_3266, 
        n5_adj_3267, n44670, n46583, n19_adj_3268, n6_adj_3269, n5_adj_3270, 
        n44695, n44696, n44667, n19_adj_3271, n46974, n5_adj_3272, 
        n44692, n44693, n44642, n44664, n38, n39, n37, n44638, 
        n46, n44640, n63_adj_3273, n63_adj_3274, n42916, n43175, 
        n10_adj_3277, n38965, n42813, n42863, n10_adj_3278, n43114, 
        n23356, n39622, n14_adj_3279, n44450, n38900, n38998, n43036, 
        n6_adj_3280, n39315, n43152, n42936, n43304, n1692, n43307, 
        n10_adj_3281, n42883, n23431, n4_adj_3282, n8_adj_3283, n1506, 
        n43111, n43127, n23371, n23546, n43205, n42955, n16_adj_3284, 
        n43187, n43289, n42868, n17_adj_3285, n15_adj_3286, n38926, 
        n42791, n43096, n43062, n12_adj_3287, n22703, n43268, n39004, 
        n23071, n23368, n23522, n44332, n49354, n43334, n42836, 
        n63_adj_3288;
    wire [31:0]\FRAME_MATCHER.state_31__N_1892 ;
    
    wire n6_adj_3289;
    wire [31:0]\FRAME_MATCHER.state_31__N_1988 ;
    
    wire n113, n11_adj_3290, n13_adj_3291, n34109, n10_adj_3292, n44037, 
        n42865, n23485, n42752, n22664, n42974, n42948, n43156, 
        n22187, n43292, n43199, n1512, n22700, n43280, n42789, 
        n22292, n1608, n42871, n10_adj_3293, n23335, n22712, n23128, 
        n43159, n42694, n20285, n22510, n43165, n44266, n22518, 
        n10_adj_3294, n22517, n22967, n16_adj_3295, n42786, n43020, 
        n6_adj_3296, n4_adj_3297, n29027, n39653, n43325, n10_adj_3298, 
        n22570, n42746, n35, n26_adj_3299, n36, n44306, n34, n40, 
        n38_adj_3300, n39_adj_3301, n37_adj_3302, n22636, n10_adj_3303, 
        n44634, n22422, n16_adj_3304, n17_adj_3305, n22501, n10_adj_3306, 
        n10_adj_3307, n14_adj_3308, n22544, n18_adj_3309, n20_adj_3310, 
        n15_adj_3311, n16_adj_3312, n17_adj_3313, n19202, n20_adj_3314, 
        n19_adj_3315, n49348, n44636, n43124, n22416, n4_adj_3316, 
        n44, n20211, n40_adj_3317, n23194, n43265, n6_adj_3318, 
        n10_adj_3319, n38682, n745, n48, n42874, n49342, n49336, 
        n2_adj_3321, n49330, n16_adj_3322, n38984, n43211, n42987, 
        n5_adj_3323, n42826, n43169, n42762, n23000, n42929, n1713, 
        n1592, n42714, n28467, n42723, n38679, n8_adj_3324, n22766, 
        n42886, n38980, n23326, n12_adj_3325, n39334, n42749, n44449, 
        n39432, n38994, n1661, n44381, n14_adj_3326, n43331, n42857, 
        n15_adj_3327, n39342, n39601, n42776, n28540, n22675, n23488, 
        n42889, n23243, n22639, n43250, n43087, n43215, n43023, 
        n22720, n12_adj_3328, n42880, n43190, n42945, n12_adj_3329, 
        n43301, n23317, n42977, n12_adj_3330, n44360, n20_adj_3331, 
        n38986, n23, n44199, n23096, n43277, n22, n26_adj_3332, 
        n44382, n42939, n38_adj_3333, n36_adj_3334, n43202, n37_adj_3335, 
        n40_adj_3336, n44_adj_3337, n39_adj_3338, n12_adj_3339, n43093, 
        n10_adj_3340, n6_adj_3341, n43108, n23329, n22_adj_3342, n20_adj_3343, 
        n24, n6_adj_3344, n23151, n42809, n42779, n42898, n10_adj_3345, 
        n14_adj_3346, n22738, n42799, n43218, n43002, n42860, n52, 
        n60_adj_3347, n58_adj_3348, n59_adj_3349, n57_adj_3350, n38_adj_3351, 
        n54, n56_adj_3352, n55_adj_3353, n66, n61_adj_3354, n43121, 
        n23313, n39012, n38931, n42964, n42932, n18_adj_3356, n20_adj_3357, 
        n12_adj_3358, n38920, n12_adj_3359, n7_adj_3360, n12_adj_3361;
    
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n24271));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n24270));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 select_278_Select_16_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [16]), .O(n3_c));
    defparam select_278_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n24269));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n24268));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 select_278_Select_17_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_3110));
    defparam select_278_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_18_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_3111));
    defparam select_278_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[8] [4]), .I1(n23449), .I2(\data_in_frame[8] [6]), 
            .I3(n23233), .O(n43133));   // verilog/coms.v(69[16:41])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_278_Select_19_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_3112));
    defparam select_278_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_CARRY add_41_8 (.CI(n36460), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n36461));
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n24267));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 select_278_Select_20_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_3113));
    defparam select_278_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFF Kd_i7 (.Q(\Kd[7] ), .C(clk32MHz), .D(n24344));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n24343));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n24342));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n24341));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 select_278_Select_21_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_3114));
    defparam select_278_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n24266));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n24340));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n24339));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 select_278_Select_22_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_3115));
    defparam select_278_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n24265));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 select_278_Select_23_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_3116));
    defparam select_278_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_24_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_3117));
    defparam select_278_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_25_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_3118));
    defparam select_278_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_26_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_3119));
    defparam select_278_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_27_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_3120));
    defparam select_278_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_4_lut_adj_829 (.I0(\data_in_frame[8] [4]), .I1(n23449), 
            .I2(n23229), .I3(n23168), .O(n43102));   // verilog/coms.v(69[16:41])
    defparam i2_3_lut_4_lut_adj_829.LUT_INIT = 16'h6996;
    SB_LUT4 select_278_Select_28_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_3121));
    defparam select_278_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_29_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_3122));
    defparam select_278_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_30_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_3123));
    defparam select_278_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i5_3_lut_4_lut (.I0(n43885), .I1(\data_in_frame[17] [0]), .I2(\data_in_frame[12] [5]), 
            .I3(\data_in_frame[19] [1]), .O(n14));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_278_Select_31_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_3124));
    defparam select_278_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i10605_3_lut_4_lut (.I0(n8), .I1(n42698), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n24023));
    defparam i10605_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n24338));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10606_3_lut_4_lut (.I0(n8), .I1(n42698), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n24024));
    defparam i10606_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10607_3_lut_4_lut (.I0(n8), .I1(n42698), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n24025));
    defparam i10607_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10608_3_lut_4_lut (.I0(n8), .I1(n42698), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n24026));
    defparam i10608_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n24264));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n24337));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10609_3_lut_4_lut (.I0(n8), .I1(n42698), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n24027));
    defparam i10609_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10610_3_lut_4_lut (.I0(n8), .I1(n42698), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n24028));
    defparam i10610_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10611_3_lut_4_lut (.I0(n8), .I1(n42698), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n24029));
    defparam i10611_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_830 (.I0(n43885), .I1(\data_in_frame[17] [0]), 
            .I2(\data_in_frame[17] [6]), .I3(n23479), .O(n14_adj_3125));
    defparam i5_3_lut_4_lut_adj_830.LUT_INIT = 16'h9669;
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n24336));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n24335));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n24377));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_7_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n36459), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10612_3_lut_4_lut (.I0(n8), .I1(n42698), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n24030));
    defparam i10612_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10597_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42698), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n24015));
    defparam i10597_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10598_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42698), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n24016));
    defparam i10598_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n24334));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n24333));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n24332));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n24331));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n24263));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_20 (.CI(n36472), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n36473));
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n24330));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n24329));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n24328));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n24327));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n24326));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n24325));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n24324));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n24323));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10599_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42698), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n24017));
    defparam i10599_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n24322));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n24321));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n24320));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n24319));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10600_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42698), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n24018));
    defparam i10600_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_41_19_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n36471), .O(n2_adj_3127)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_19_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n24318));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n24262));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n24261));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_7 (.CI(n36459), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n36460));
    SB_LUT4 i10601_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42698), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n24019));
    defparam i10601_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_41_19 (.CI(n36471), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n36472));
    SB_LUT4 i10602_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42698), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n24020));
    defparam i10602_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_41_18_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n36470), .O(n2_adj_3128)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_18 (.CI(n36470), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n36471));
    SB_LUT4 i10603_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42698), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n24021));
    defparam i10603_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10604_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42698), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n24022));
    defparam i10604_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_41_6_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n36458), .O(n2_adj_3129)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_41_17_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n36469), .O(n2_adj_3130)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_831 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[13] [4]), .I3(Kp_23__N_838), .O(n43148));   // verilog/coms.v(71[16:43])
    defparam i2_3_lut_4_lut_adj_831.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_832 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(n23038), .I3(\data_in_frame[18] [0]), .O(n39055));   // verilog/coms.v(71[16:43])
    defparam i2_3_lut_4_lut_adj_832.LUT_INIT = 16'h6996;
    SB_LUT4 i10589_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42698), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n24007));
    defparam i10589_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF deadband_i0_i9 (.Q(\deadband[9] ), .C(clk32MHz), .D(n24490));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10590_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42698), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n24008));
    defparam i10590_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF deadband_i0_i8 (.Q(\deadband[8] ), .C(clk32MHz), .D(n24489));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i7 (.Q(\deadband[7] ), .C(clk32MHz), .D(n24488));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i6 (.Q(\deadband[6] ), .C(clk32MHz), .D(n24487));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i5 (.Q(\deadband[5] ), .C(clk32MHz), .D(n24486));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i4 (.Q(\deadband[4] ), .C(clk32MHz), .D(n24485));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i3 (.Q(\deadband[3] ), .C(clk32MHz), .D(n24484));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i2 (.Q(\deadband[2] ), .C(clk32MHz), .D(n24483));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10591_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42698), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n24009));
    defparam i10591_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(VCC_net), .D(n24482));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i1 (.Q(\deadband[1] ), .C(clk32MHz), .D(n24479));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n24478));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n24477));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n24476));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n24475));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n24474));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n24473));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n24472));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n24471));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n24470));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n24469));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n24468));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n24467));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n24466));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n24465));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n24464));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n24463));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n24462));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n24461));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n24460));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n24459));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n24458));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n24457));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n24456));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter_c[1]), .C(clk32MHz), 
           .D(n23891));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n24260));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n24306));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n24259));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n24305));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n24258));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n24304));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n24257));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n24303));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n24256));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n24302));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n24255));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n24301));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n24254));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n24300));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n24253));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n24299));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n24252));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n24298));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n24251));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n24297));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n24250));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n24296));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n24249));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n24295));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n24248));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n24294));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n24247));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n24293));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n24246));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n24292));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n24291));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n24290));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk32MHz), 
           .D(n24289));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk32MHz), 
           .D(n24288));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk32MHz), 
           .D(n24287));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n24286));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n24285));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5][2] ), .C(clk32MHz), 
           .D(n24284));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n24283));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n24282));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n24376));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n24375));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n24374));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n24373));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n24372));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n24371));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n24370));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n24245));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n24244));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n24243));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n24242));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n24241));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n24281));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n24280));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n24279));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n24278));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n24277));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n24276));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n24240));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n24239));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n24275));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10592_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42698), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n24010));
    defparam i10592_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n24274));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n24238));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n24369));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10593_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42698), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n24011));
    defparam i10593_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n24237));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n24317));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10594_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42698), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n24012));
    defparam i10594_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10595_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42698), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n24013));
    defparam i10595_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10596_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42698), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n24014));
    defparam i10596_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10581_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42698), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n23999));
    defparam i10581_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10582_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42698), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n24000));
    defparam i10582_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10583_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42698), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n24001));
    defparam i10583_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10584_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42698), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n24002));
    defparam i10584_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n24236));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n24235));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n24234));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n24233));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10585_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42698), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n24003));
    defparam i10585_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n24232));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n24231));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n24230));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n24229));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n24228));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n24227));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n24316));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n24226));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n24225));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n24224));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n24223));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n24222));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n24221));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n24220));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_6 (.CI(n36458), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n36459));
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n24219));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n24315));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10586_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42698), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n24004));
    defparam i10586_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n24314));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n24218));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n24217));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n24216));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n24215));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10587_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42698), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n24005));
    defparam i10587_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n24214));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n24213));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n24212));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n24211));   // verilog/coms.v(125[12] 284[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3221  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n24210));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10588_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42698), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n24006));
    defparam i10588_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n24209));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n24273));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n24368));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10573_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42698), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n23991));
    defparam i10573_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n24208));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n24207));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10574_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42698), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n23992));
    defparam i10574_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n24206));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n24205));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n24313));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n24204));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n24312));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n24203));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n24379));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n24202));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n24367));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10575_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42698), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n23993));
    defparam i10575_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10576_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42698), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n23994));
    defparam i10576_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n24366));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n24365));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10577_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42698), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n23995));
    defparam i10577_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n24364));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_4_lut_adj_833 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[16] [7]), 
            .I2(Kp_23__N_785), .I3(n43313), .O(n23513));
    defparam i2_3_lut_4_lut_adj_833.LUT_INIT = 16'h6996;
    SB_LUT4 i10578_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42698), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n23996));
    defparam i10578_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n24363));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10579_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42698), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n23997));
    defparam i10579_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_834 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[16] [7]), 
            .I2(\data_in_frame[16] [5]), .I3(n43105), .O(Kp_23__N_994));
    defparam i2_3_lut_4_lut_adj_834.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n24201));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n24200));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n24199));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n24198));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n24197));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n24196));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n24195));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n24194));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n24193));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n24192));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n24191));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n24190));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n24189));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n24188));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_4_lut_adj_835 (.I0(n43885), .I1(n39460), .I2(Kp_23__N_945), 
            .I3(n39629), .O(n23026));
    defparam i2_3_lut_4_lut_adj_835.LUT_INIT = 16'h9669;
    SB_LUT4 i10580_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42698), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n23998));
    defparam i10580_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n24187));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n24186));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n22524), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n22525));   // verilog/coms.v(211[5:21])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i29087_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n22524), 
            .I2(n22520), .I3(\FRAME_MATCHER.state[0] ), .O(n28588));   // verilog/coms.v(211[5:21])
    defparam i29087_3_lut_4_lut.LUT_INIT = 16'he0ff;
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n24185));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(n43885), .I1(n39460), .I2(n43142), .I3(GND_net), 
            .O(n43139));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i3_3_lut_4_lut (.I0(n43885), .I1(n39460), .I2(n23513), .I3(\data_in_frame[19] [7]), 
            .O(n8_adj_3134));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n24184));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_17 (.CI(n36469), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n36470));
    SB_LUT4 i10565_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42698), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n23983));
    defparam i10565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n24183));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n24182));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n24181));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_3_lut_adj_836 (.I0(n23462), .I1(\data_in_frame[17] [5]), 
            .I2(n39055), .I3(GND_net), .O(n6));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_836.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n24180));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10566_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42698), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n23984));
    defparam i10566_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n24179));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10567_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42698), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n23985));
    defparam i10567_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n24178));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n24177));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n24176));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n24175));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n24174));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n24378));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n24173));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n24172));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n24171));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n24170));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n24169));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n24168));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n24167));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n24166));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n24165));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n24164));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10568_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42698), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n23986));
    defparam i10568_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n24163));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n24162));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n24161));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n24160));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n24159));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
           .D(n24158));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i5_3_lut_4_lut_adj_837 (.I0(n23462), .I1(\data_in_frame[17] [5]), 
            .I2(n22942), .I3(n10), .O(n43172));   // verilog/coms.v(73[16:43])
    defparam i5_3_lut_4_lut_adj_837.LUT_INIT = 16'h6996;
    SB_LUT4 i10569_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42698), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n23987));
    defparam i10569_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n24157));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n24156));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n24155));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10570_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42698), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n23988));
    defparam i10570_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10571_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42698), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n23989));
    defparam i10571_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n24154));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n24153));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n24152));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n24151));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n24150));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10572_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42698), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n23990));
    defparam i10572_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n24149));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n24148));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n24147));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n24146));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n24145));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n24362));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n24144));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n24361));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n24143));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n24142));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n24141));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n24140));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n24139));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n24138));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n24137));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n24136));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n24135));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n24134));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n24133));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n24132));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n24131));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n24130));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10846_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[14]), .I3(\data_out_frame[7] [6]), .O(n24264));
    defparam i10846_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n24129));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n24128));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n24127));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n24126));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10849_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[11]), .I3(\data_out_frame[7] [3]), .O(n24267));
    defparam i10849_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10742_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[6]), .I3(\data_out_frame[20] [6]), .O(n24160));
    defparam i10742_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n24125));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10859_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[17]), .I3(\data_out_frame[6] [1]), .O(n24277));
    defparam i10859_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n24124));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n24123));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n24122));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n24121));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n24120));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n24119));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n24118));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10804_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[8]), .I3(\data_out_frame[13] [0]), .O(n24222));
    defparam i10804_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n24117));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n24116));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n24115));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n24114));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n24113));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n24112));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n24111));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n24110));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_16_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n36468), .O(n2_adj_3136)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_16_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n24109));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10801_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[11]), .I3(\data_out_frame[13] [3]), .O(n24219));
    defparam i10801_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY add_41_16 (.CI(n36468), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n36469));
    SB_LUT4 i10803_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[9]), .I3(\data_out_frame[13] [1]), .O(n24221));
    defparam i10803_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n24360));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10802_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[10]), .I3(\data_out_frame[13] [2]), .O(n24220));
    defparam i10802_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10805_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[23]), .I3(\data_out_frame[12] [7]), .O(n24223));
    defparam i10805_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_838 (.I0(\FRAME_MATCHER.state[3] ), .I1(n22528), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(GND_net), .O(n22524));   // verilog/coms.v(147[5:27])
    defparam i1_2_lut_3_lut_adj_838.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_839 (.I0(\FRAME_MATCHER.state[3] ), .I1(n22528), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(GND_net), .O(n22520));   // verilog/coms.v(147[5:27])
    defparam i1_2_lut_3_lut_adj_839.LUT_INIT = 16'hfefe;
    SB_LUT4 i10806_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[22]), .I3(\data_out_frame[12] [6]), .O(n24224));
    defparam i10806_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10807_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[21]), .I3(\data_out_frame[12] [5]), .O(n24225));
    defparam i10807_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter_c[2]), .C(clk32MHz), 
           .D(n23894));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_5_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n36457), .O(n2_adj_3137)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n24108));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_5 (.CI(n36457), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n36458));
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n24387));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10808_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[20]), .I3(\data_out_frame[12] [4]), .O(n24226));
    defparam i10808_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n24107));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_15_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n36467), .O(n2_adj_3138)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31329_4_lut (.I0(byte_transmit_counter[0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter_c[2]), 
            .O(n46842));   // verilog/coms.v(103[34:55])
    defparam i31329_4_lut.LUT_INIT = 16'h880a;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29171_4_lut (.I0(n19), .I1(\data_out_frame[22]_c [0]), .I2(byte_transmit_counter_c[1]), 
            .I3(byte_transmit_counter[0]), .O(n44683));
    defparam i29171_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29172_3_lut (.I0(n49387), .I1(n44683), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44684));
    defparam i29172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29149_4_lut (.I0(n5_c), .I1(n46842), .I2(byte_transmit_counter_c[2]), 
            .I3(byte_transmit_counter_c[1]), .O(n44661));
    defparam i29149_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i10783_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[21]), .I3(\data_out_frame[15] [5]), .O(n24201));
    defparam i10783_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY add_41_15 (.CI(n36467), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n36468));
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n24106));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n24105));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i29151_4_lut (.I0(n44661), .I1(n44684), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44663));
    defparam i29151_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29150_3_lut (.I0(n49471), .I1(n49477), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44662));
    defparam i29150_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n24104));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n24103));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[9] [7]), .O(n43193));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10810_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[18]), .I3(\data_out_frame[12] [2]), .O(n24228));
    defparam i10810_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10811_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[17]), .I3(\data_out_frame[12] [1]), .O(n24229));
    defparam i10811_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10812_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[16]), .I3(\data_out_frame[12] [0]), .O(n24230));
    defparam i10812_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10813_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[7]), .I3(\data_out_frame[11] [7]), .O(n24231));
    defparam i10813_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10814_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[6]), .I3(\data_out_frame[11] [6]), .O(n24232));
    defparam i10814_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n24102));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n24101));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n24100));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n24099));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n24098));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10815_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[5]), .I3(\data_out_frame[11] [5]), .O(n24233));
    defparam i10815_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10816_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[4]), .I3(\data_out_frame[11] [4]), .O(n24234));
    defparam i10816_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_41_14_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n36466), .O(n2_adj_3139)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_14_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n24097));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10817_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[3]), .I3(\data_out_frame[11] [3]), .O(n24235));
    defparam i10817_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n24096));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n24095));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n24094));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n24093));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n24092));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10819_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[1]), .I3(\data_out_frame[11] [1]), .O(n24237));
    defparam i10819_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10820_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[0]), .I3(\data_out_frame[11] [0]), .O(n24238));
    defparam i10820_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n24091));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n24090));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n24089));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10856_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[20]), .I3(\data_out_frame[6] [4]), .O(n24274));
    defparam i10856_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10857_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[19]), .I3(\data_out_frame[6] [3]), .O(n24275));
    defparam i10857_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10858_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[18]), .I3(\data_out_frame[6] [2]), .O(n24276));
    defparam i10858_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10861_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(control_mode[7]), .I3(\data_out_frame[5] [7]), .O(n24279));
    defparam i10861_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10860_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[16]), .I3(\data_out_frame[6] [0]), .O(n24278));
    defparam i10860_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10825_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[11]), .I3(\data_out_frame[10] [3]), .O(n24243));
    defparam i10825_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10823_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[13]), .I3(\data_out_frame[10] [5]), .O(n24241));
    defparam i10823_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10824_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[12]), .I3(\data_out_frame[10] [4]), .O(n24242));
    defparam i10824_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n24088));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10826_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[10]), .I3(\data_out_frame[10] [2]), .O(n24244));
    defparam i10826_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10868_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(control_mode[0]), .I3(\data_out_frame[5] [0]), .O(n24286));
    defparam i10868_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut (.I0(n42743), .I1(n39501), .I2(n42612), .I3(GND_net), 
            .O(n22528));   // verilog/coms.v(147[5:27])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_41_14 (.CI(n36466), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n36467));
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n24087));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10827_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[9]), .I3(\data_out_frame[10] [1]), .O(n24245));
    defparam i10827_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_840 (.I0(\data_in_frame[17] [6]), .I1(n42782), 
            .I2(n39055), .I3(GND_net), .O(n43238));
    defparam i2_3_lut_adj_840.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut (.I0(n43030), .I1(n43310), .I2(n43231), .I3(n43077), 
            .O(n39629));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_13_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n36465), .O(n2_adj_3140)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut (.I0(n23017), .I1(Kp_23__N_776), .I2(\data_in_frame[18] [1]), 
            .I3(Kp_23__N_994), .O(n10_adj_3141));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n39257), .I1(n10_adj_3141), .I2(n23026), .I3(GND_net), 
            .O(n43017));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n24086));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10864_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(control_mode[4]), .I3(\data_out_frame[5] [4]), .O(n24282));
    defparam i10864_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_841 (.I0(n43585), .I1(n8_adj_3134), .I2(n23513), 
            .I3(n43139), .O(n43071));
    defparam i4_4_lut_adj_841.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_842 (.I0(n43283), .I1(n43099), .I2(\data_in_frame[6] [6]), 
            .I3(n43133), .O(n10_adj_3142));   // verilog/coms.v(69[16:41])
    defparam i4_4_lut_adj_842.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_843 (.I0(n22891), .I1(n23266), .I2(\data_in_frame[15] [4]), 
            .I3(GND_net), .O(n23467));   // verilog/coms.v(71[16:43])
    defparam i2_3_lut_adj_843.LUT_INIT = 16'h9696;
    SB_LUT4 i10865_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(control_mode[3]), .I3(\data_out_frame[5] [3]), .O(n24283));
    defparam i10865_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_844 (.I0(\data_in_frame[19] [6]), .I1(n43136), 
            .I2(Kp_23__N_192), .I3(\data_in_frame[17] [4]), .O(n10));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_844.LUT_INIT = 16'h6996;
    SB_LUT4 i10867_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(control_mode[1]), .I3(\data_out_frame[5] [1]), .O(n24285));
    defparam i10867_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n24085));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_13 (.CI(n36465), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n36466));
    SB_LUT4 i10828_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[8]), .I3(\data_out_frame[10] [0]), .O(n24246));
    defparam i10828_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_2_lut (.I0(\data_in_frame[12] [5]), .I1(n23462), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3143));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10829_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[23]), .I3(\data_out_frame[9] [7]), .O(n24247));
    defparam i10829_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i6_4_lut (.I0(n43228), .I1(n22891), .I2(n43130), .I3(n21140), 
            .O(n14_adj_3144));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10830_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[22]), .I3(\data_out_frame[9] [6]), .O(n24248));
    defparam i10830_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7_4_lut (.I0(\data_in_frame[19] [5]), .I1(n14_adj_3144), .I2(n10_adj_3143), 
            .I3(n43225), .O(n42904));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_18__7__I_0_3244_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_785));   // verilog/coms.v(75[16:27])
    defparam data_in_frame_18__7__I_0_3244_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10832_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[20]), .I3(\data_out_frame[9] [4]), .O(n24250));
    defparam i10832_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n24084));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10837_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[7]), .I3(\data_out_frame[8] [7]), .O(n24255));
    defparam i10837_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10834_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[18]), .I3(\data_out_frame[9] [2]), .O(n24252));
    defparam i10834_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42995));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10835_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[17]), .I3(\data_out_frame[9] [1]), .O(n24253));
    defparam i10835_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n24083));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i3_4_lut_adj_845 (.I0(\data_in_frame[18] [1]), .I1(n43234), 
            .I2(n43064), .I3(n42995), .O(n43313));
    defparam i3_4_lut_adj_845.LUT_INIT = 16'h6996;
    SB_LUT4 i10836_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[16]), .I3(\data_out_frame[9] [0]), .O(n24254));
    defparam i10836_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10838_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[6]), .I3(\data_out_frame[8] [6]), .O(n24256));
    defparam i10838_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10839_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[5]), .I3(\data_out_frame[8] [5]), .O(n24257));
    defparam i10839_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10840_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[4]), .I3(\data_out_frame[8] [4]), .O(n24258));
    defparam i10840_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_41_4_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n36456), .O(n2_adj_3145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_846 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43225));
    defparam i1_2_lut_adj_846.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_847 (.I0(n43225), .I1(\data_in_frame[16] [5]), 
            .I2(\data_in_frame[17] [7]), .I3(n43011), .O(n15));
    defparam i6_4_lut_adj_847.LUT_INIT = 16'h6996;
    SB_LUT4 i10841_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[3]), .I3(\data_out_frame[8] [3]), .O(n24259));
    defparam i10841_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(Kp_23__N_776), .I2(n14_adj_3125), 
            .I3(\data_in_frame[17] [5]), .O(n43585));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n24082));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10842_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[2]), .I3(\data_out_frame[8] [2]), .O(n24260));
    defparam i10842_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10843_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[1]), .I3(\data_out_frame[8] [1]), .O(n24261));
    defparam i10843_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10844_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[0]), .I3(\data_out_frame[8] [0]), .O(n24262));
    defparam i10844_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_848 (.I0(\data_in_frame[15] [3]), .I1(n43585), 
            .I2(n23208), .I3(n6), .O(n43142));
    defparam i4_4_lut_adj_848.LUT_INIT = 16'h9669;
    SB_LUT4 i10845_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[15]), .I3(\data_out_frame[7] [7]), .O(n24263));
    defparam i10845_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10847_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[13]), .I3(\data_out_frame[7] [5]), .O(n24265));
    defparam i10847_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n24386));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_12_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n36464), .O(n2_adj_3146)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10743_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[5]), .I3(\data_out_frame[20] [5]), .O(n24161));
    defparam i10743_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_849 (.I0(n39029), .I1(n43068), .I2(Kp_23__N_994), 
            .I3(GND_net), .O(n43885));
    defparam i2_3_lut_adj_849.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_850 (.I0(n42969), .I1(\data_in_frame[14] [5]), 
            .I2(n23018), .I3(GND_net), .O(n39029));
    defparam i2_3_lut_adj_850.LUT_INIT = 16'h9696;
    SB_LUT4 i10854_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[22]), .I3(\data_out_frame[6] [6]), .O(n24272));
    defparam i10854_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_851 (.I0(n43295), .I1(n43322), .I2(n43005), .I3(GND_net), 
            .O(n22942));   // verilog/coms.v(82[17:28])
    defparam i2_3_lut_adj_851.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_852 (.I0(Kp_23__N_945), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n22801));
    defparam i1_2_lut_adj_852.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_853 (.I0(n43059), .I1(\data_in_frame[9] [6]), .I2(n43184), 
            .I3(n43298), .O(n15_adj_3147));
    defparam i6_4_lut_adj_853.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_854 (.I0(n15_adj_3147), .I1(n43084), .I2(n14_adj_3148), 
            .I3(\data_in_frame[7] [4]), .O(n44327));
    defparam i8_4_lut_adj_854.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_855 (.I0(n44318), .I1(n44327), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_776));
    defparam i1_2_lut_adj_855.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter_c[1]), 
            .I1(n19_adj_3149), .I2(n46624), .I3(byte_transmit_counter_c[2]), 
            .O(n49480));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49480_bdd_4_lut (.I0(n49480), .I1(n17), .I2(n16), .I3(byte_transmit_counter_c[2]), 
            .O(n49483));
    defparam n49480_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n49474));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49474_bdd_4_lut (.I0(n49474), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n49477));
    defparam n49474_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33938 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n49468));
    defparam byte_transmit_counter_0__bdd_4_lut_33938.LUT_INIT = 16'he4aa;
    SB_LUT4 n49468_bdd_4_lut (.I0(n49468), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n49471));
    defparam n49468_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33933 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter_c[1]), .O(n49462));
    defparam byte_transmit_counter_0__bdd_4_lut_33933.LUT_INIT = 16'he4aa;
    SB_LUT4 n49462_bdd_4_lut (.I0(n49462), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter_c[1]), 
            .O(n49465));
    defparam n49462_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33928 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter_c[1]), .O(n49456));
    defparam byte_transmit_counter_0__bdd_4_lut_33928.LUT_INIT = 16'he4aa;
    SB_LUT4 n49456_bdd_4_lut (.I0(n49456), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter_c[1]), 
            .O(n49459));
    defparam n49456_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_856 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n22682));
    defparam i1_2_lut_adj_856.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_857 (.I0(n43834), .I1(\data_in_frame[13] [4]), 
            .I2(n22885), .I3(GND_net), .O(n42782));   // verilog/coms.v(71[16:43])
    defparam i2_3_lut_adj_857.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_858 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3150));   // verilog/coms.v(69[16:41])
    defparam i1_2_lut_adj_858.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_859 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[9] [0]), .I3(n6_adj_3150), .O(n43099));   // verilog/coms.v(69[16:41])
    defparam i4_4_lut_adj_859.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_860 (.I0(n42958), .I1(\data_in_frame[11] [1]), 
            .I2(\data_in_frame[13] [3]), .I3(n42999), .O(n10_adj_3151));   // verilog/coms.v(71[16:43])
    defparam i4_4_lut_adj_860.LUT_INIT = 16'h6996;
    SB_LUT4 i10741_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[7]), .I3(\data_out_frame[20] [7]), .O(n24159));
    defparam i10741_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_861 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43221));   // verilog/coms.v(82[17:28])
    defparam i1_2_lut_adj_861.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_862 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43130));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_862.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_863 (.I0(\data_in_frame[8] [7]), .I1(n22858), .I2(GND_net), 
            .I3(GND_net), .O(n43283));   // verilog/coms.v(69[16:41])
    defparam i1_2_lut_adj_863.LUT_INIT = 16'h6666;
    SB_LUT4 i10744_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[4]), .I3(\data_out_frame[20] [4]), .O(n24162));
    defparam i10744_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 data_in_frame_12__7__I_0_3240_2_lut (.I0(\data_in_frame[12] [7]), 
            .I1(\data_in_frame[12] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_192));   // verilog/coms.v(68[16:27])
    defparam data_in_frame_12__7__I_0_3240_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_864 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n23208));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_864.LUT_INIT = 16'h6666;
    SB_LUT4 i20_4_lut (.I0(n23208), .I1(\data_in_frame[8] [4]), .I2(n43056), 
            .I3(n7), .O(n56));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(Kp_23__N_192), .I1(n43148), .I2(n42913), .I3(n43834), 
            .O(n55));
    defparam i19_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i27_4_lut (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[14] [2]), 
            .I2(\data_in_frame[10] [5]), .I3(\data_in_frame[15] [2]), .O(n63_c));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(n43130), .I1(n43053), .I2(n43074), .I3(n42925), 
            .O(n60));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n42765), .I1(\data_in_frame[7] [0]), .I2(n22770), 
            .I3(\data_in_frame[11] [4]), .O(n58));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10745_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[3]), .I3(\data_out_frame[20] [3]), .O(n24163));
    defparam i10745_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10747_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[1]), .I3(\data_out_frame[20] [1]), .O(n24165));
    defparam i10747_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i23_4_lut (.I0(\data_in_frame[13] [0]), .I1(n43262), .I2(\data_in_frame[14] [4]), 
            .I3(n43221), .O(n59));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(\data_in_frame[14] [3]), .I1(n43099), .I2(n43244), 
            .I3(n43050), .O(n57));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[9] [6]), .I3(\data_in_frame[12] [5]), .O(n62));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i32_3_lut (.I0(n63_c), .I1(n55), .I2(n56), .I3(GND_net), 
            .O(n68));
    defparam i32_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i25_4_lut (.I0(n42907), .I1(Kp_23__N_319), .I2(\data_in_frame[14] [1]), 
            .I3(n23266), .O(n61));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut (.I0(n57), .I1(n59), .I2(n58), .I3(n60), .O(n69));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10748_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[0]), .I3(\data_out_frame[20] [0]), .O(n24166));
    defparam i10748_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i35_4_lut (.I0(n69), .I1(n61), .I2(n68), .I3(n62), .O(n39460));
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10749_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[15]), .I3(\data_out_frame[19] [7]), .O(n24167));
    defparam i10749_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10750_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[14]), .I3(\data_out_frame[19] [6]), .O(n24168));
    defparam i10750_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_865 (.I0(n23266), .I1(n42782), .I2(\data_in_frame[15] [5]), 
            .I3(GND_net), .O(n23479));
    defparam i2_3_lut_adj_865.LUT_INIT = 16'h9696;
    SB_LUT4 i10751_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[13]), .I3(\data_out_frame[19] [5]), .O(n24169));
    defparam i10751_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_866 (.I0(n23479), .I1(n39460), .I2(\data_in_frame[16] [0]), 
            .I3(GND_net), .O(n43068));
    defparam i2_3_lut_adj_866.LUT_INIT = 16'h9696;
    SB_LUT4 i10752_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[12]), .I3(\data_out_frame[19] [4]), .O(n24170));
    defparam i10752_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i5_4_lut (.I0(n43253), .I1(n43274), .I2(\data_in_frame[8] [1]), 
            .I3(n43181), .O(n12));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_867 (.I0(\data_in_frame[7] [7]), .I1(n12), .I2(n43322), 
            .I3(n43008), .O(n21140));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_867.LUT_INIT = 16'h6996;
    SB_LUT4 i10753_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[11]), .I3(\data_out_frame[19] [3]), .O(n24171));
    defparam i10753_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i6_4_lut_adj_868 (.I0(n21140), .I1(\data_in_frame[14] [6]), 
            .I2(n43068), .I3(n43105), .O(n15_adj_3152));
    defparam i6_4_lut_adj_868.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_869 (.I0(n15_adj_3152), .I1(n42919), .I2(n14), 
            .I3(n23018), .O(n43026));
    defparam i8_4_lut_adj_869.LUT_INIT = 16'h6996;
    SB_LUT4 i10754_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[10]), .I3(\data_out_frame[19] [2]), .O(n24172));
    defparam i10754_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i5_4_lut_adj_870 (.I0(n22801), .I1(n43090), .I2(\data_in_frame[12] [6]), 
            .I3(n22942), .O(n12_adj_3153));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_871 (.I0(\data_in_frame[17] [0]), .I1(n12_adj_3153), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[17] [1]), .O(n43241));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_872 (.I0(n42904), .I1(n43172), .I2(n23467), .I3(GND_net), 
            .O(n42901));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_adj_872.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_873 (.I0(n43196), .I1(n42901), .I2(n43241), .I3(n43026), 
            .O(n8_adj_3154));
    defparam i3_4_lut_adj_873.LUT_INIT = 16'h6996;
    SB_LUT4 i4_3_lut (.I0(\data_in_frame[19] [7]), .I1(n8_adj_3154), .I2(n42951), 
            .I3(GND_net), .O(n23470));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i10756_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[8]), .I3(\data_out_frame[19] [0]), .O(n24174));
    defparam i10756_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10757_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[23]), .I3(\data_out_frame[18] [7]), .O(n24175));
    defparam i10757_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n24385));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_564_9_lut (.I0(byte_transmit_counter_c[7]), .I1(byte_transmit_counter_c[7]), 
            .I2(n3840), .I3(n36492), .O(n23907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_564_9_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i3_4_lut_adj_874 (.I0(\data_in_frame[5] [6]), .I1(n23449), .I2(\data_in_frame[8] [2]), 
            .I3(Kp_23__N_458), .O(n43295));   // verilog/coms.v(69[16:41])
    defparam i3_4_lut_adj_874.LUT_INIT = 16'h6996;
    SB_LUT4 i10758_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[22]), .I3(\data_out_frame[18] [6]), .O(n24176));
    defparam i10758_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_875 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43181));
    defparam i1_2_lut_adj_875.LUT_INIT = 16'h6666;
    SB_LUT4 i10759_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[21]), .I3(\data_out_frame[18] [5]), .O(n24177));
    defparam i10759_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10760_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[20]), .I3(\data_out_frame[18] [4]), .O(n24178));
    defparam i10760_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_876 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[14] [7]), .I3(GND_net), .O(n42765));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_876.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_877 (.I0(n43181), .I1(n22826), .I2(\data_in_frame[12] [4]), 
            .I3(n43295), .O(n10_adj_3155));
    defparam i4_4_lut_adj_877.LUT_INIT = 16'h6996;
    SB_LUT4 i10761_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[19]), .I3(\data_out_frame[18] [3]), .O(n24179));
    defparam i10761_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_878 (.I0(n23018), .I1(n43102), .I2(n42765), .I3(n43271), 
            .O(n43090));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_878.LUT_INIT = 16'h6996;
    SB_LUT4 add_564_8_lut (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[6]), 
            .I2(n3840), .I3(n36491), .O(n23904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_564_8_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_564_8 (.CI(n36491), .I0(byte_transmit_counter_c[6]), .I1(n3840), 
            .CO(n36492));
    SB_LUT4 add_564_7_lut (.I0(byte_transmit_counter_c[5]), .I1(byte_transmit_counter_c[5]), 
            .I2(n3840), .I3(n36490), .O(n23901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_564_7_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i3_4_lut_adj_879 (.I0(\data_in_frame[4] [0]), .I1(n43042), .I2(\data_in_frame[1] [6]), 
            .I3(\data_in_frame[1] [4]), .O(n23449));   // verilog/coms.v(82[17:28])
    defparam i3_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n24081));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10763_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[17]), .I3(\data_out_frame[18] [1]), .O(n24181));
    defparam i10763_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10762_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[18]), .I3(\data_out_frame[18] [2]), .O(n24180));
    defparam i10762_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n24080));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33923 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter_c[1]), .O(n49450));
    defparam byte_transmit_counter_0__bdd_4_lut_33923.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n24079));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49450_bdd_4_lut (.I0(n49450), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n49453));
    defparam n49450_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n24078));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n24077));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10764_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[16]), .I3(\data_out_frame[18] [0]), .O(n24182));
    defparam i10764_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33918 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter_c[1]), .O(n49444));
    defparam byte_transmit_counter_0__bdd_4_lut_33918.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n24076));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49444_bdd_4_lut (.I0(n49444), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n49447));
    defparam n49444_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n24075));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n24074));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33913 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter_c[1]), .O(n49438));
    defparam byte_transmit_counter_0__bdd_4_lut_33913.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n24073));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49438_bdd_4_lut (.I0(n49438), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n49441));
    defparam n49438_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n24072));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n24071));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33908 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n49432));
    defparam byte_transmit_counter_0__bdd_4_lut_33908.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n24070));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49432_bdd_4_lut (.I0(n49432), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n49435));
    defparam n49432_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n24069));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n24068));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33903 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n49426));
    defparam byte_transmit_counter_0__bdd_4_lut_33903.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n24067));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49426_bdd_4_lut (.I0(n49426), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n49429));
    defparam n49426_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n24066));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n24065));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33898 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n49420));
    defparam byte_transmit_counter_0__bdd_4_lut_33898.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n24064));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49420_bdd_4_lut (.I0(n49420), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n49423));
    defparam n49420_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n24063));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n24062));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_adj_880 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n23168));   // verilog/coms.v(70[16:42])
    defparam i1_2_lut_adj_880.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33893 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n49414));
    defparam byte_transmit_counter_0__bdd_4_lut_33893.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n24061));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49414_bdd_4_lut (.I0(n49414), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n48097));
    defparam n49414_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n24060));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n24059));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33888 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n49408));
    defparam byte_transmit_counter_0__bdd_4_lut_33888.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n24058));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49408_bdd_4_lut (.I0(n49408), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n44739));
    defparam n49408_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n24057));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n24056));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33883 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter_c[1]), .O(n49402));
    defparam byte_transmit_counter_0__bdd_4_lut_33883.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n24055));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i5_4_lut_adj_881 (.I0(n23168), .I1(n42840), .I2(\data_in_frame[13] [1]), 
            .I3(n22750), .O(n12_adj_3156));   // verilog/coms.v(72[16:43])
    defparam i5_4_lut_adj_881.LUT_INIT = 16'h6996;
    SB_LUT4 n49402_bdd_4_lut (.I0(n49402), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n49405));
    defparam n49402_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n24054));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i6_4_lut_adj_882 (.I0(\data_in_frame[11] [0]), .I1(n12_adj_3156), 
            .I2(n43133), .I3(\data_in_frame[10] [7]), .O(n23462));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_883 (.I0(n22815), .I1(n22781), .I2(\data_in_frame[15] [2]), 
            .I3(n43102), .O(n43136));   // verilog/coms.v(70[16:42])
    defparam i3_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_884 (.I0(\data_in_frame[1] [7]), .I1(n43008), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3157));   // verilog/coms.v(225[9:81])
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_LUT4 i10765_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[7]), .I3(\data_out_frame[17] [7]), .O(n24183));
    defparam i10765_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_885 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43316));   // verilog/coms.v(225[9:81])
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_886 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43042));   // verilog/coms.v(82[17:28])
    defparam i1_2_lut_adj_886.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_887 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3158));   // verilog/coms.v(225[9:81])
    defparam i1_2_lut_adj_887.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_888 (.I0(n43253), .I1(n43042), .I2(n43316), .I3(n6_adj_3158), 
            .O(n43005));   // verilog/coms.v(225[9:81])
    defparam i4_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_889 (.I0(n22853), .I1(n42958), .I2(\data_in_frame[6] [4]), 
            .I3(GND_net), .O(n22781));   // verilog/coms.v(71[16:43])
    defparam i2_3_lut_adj_889.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_890 (.I0(\data_in_frame[6] [1]), .I1(n43005), .I2(\data_in_frame[8] [3]), 
            .I3(\data_in_frame[10] [5]), .O(n43271));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_891 (.I0(\data_in_frame[12] [7]), .I1(n43271), 
            .I2(n22781), .I3(GND_net), .O(n42840));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_adj_891.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n24311));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10766_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[6]), .I3(\data_out_frame[17] [6]), .O(n24184));
    defparam i10766_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_892 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n22815));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_892.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_893 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43059));
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_894 (.I0(\data_in_frame[5] [7]), .I1(n42829), .I2(\data_in_frame[1] [3]), 
            .I3(GND_net), .O(n23347));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_894.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_895 (.I0(n23347), .I1(n23032), .I2(\data_in_frame[8] [1]), 
            .I3(GND_net), .O(n43184));
    defparam i2_3_lut_adj_895.LUT_INIT = 16'h9696;
    SB_LUT4 i10767_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[5]), .I3(\data_out_frame[17] [5]), .O(n24185));
    defparam i10767_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10769_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[3]), .I3(\data_out_frame[17] [3]), .O(n24187));
    defparam i10769_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_896 (.I0(\data_in_frame[12] [3]), .I1(n43184), 
            .I2(\data_in_frame[10] [1]), .I3(\data_in_frame[9] [7]), .O(n10_adj_3159));
    defparam i4_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_897 (.I0(n42925), .I1(n10_adj_3159), .I2(\data_in_frame[7] [5]), 
            .I3(GND_net), .O(n42969));
    defparam i5_3_lut_adj_897.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_898 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43011));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h6666;
    SB_LUT4 i10770_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[2]), .I3(\data_out_frame[17] [2]), .O(n24188));
    defparam i10770_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_2_lut_adj_899 (.I0(\data_in_frame[15] [1]), .I1(n42969), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3160));   // verilog/coms.v(75[16:27])
    defparam i2_2_lut_adj_899.LUT_INIT = 16'h6666;
    SB_LUT4 i10771_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[1]), .I3(\data_out_frame[17] [1]), .O(n24189));
    defparam i10771_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i6_4_lut_adj_900 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[14] [6]), 
            .I2(n43011), .I3(\data_in_frame[16] [7]), .O(n14_adj_3161));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_901 (.I0(\data_in_frame[19] [3]), .I1(n14_adj_3161), 
            .I2(n10_adj_3160), .I3(n43228), .O(n43196));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n24053));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n24052));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_4 (.CI(n36456), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n36457));
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n24051));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n24384));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n24359));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10773_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[15]), .I3(\data_out_frame[16] [7]), .O(n24191));
    defparam i10773_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10775_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[13]), .I3(\data_out_frame[16] [5]), .O(n24193));
    defparam i10775_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i5_4_lut_adj_902 (.I0(\data_in_frame[17] [2]), .I1(n43136), 
            .I2(n23462), .I3(\data_in_frame[17] [3]), .O(n12_adj_3162));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_CARRY add_564_7 (.CI(n36490), .I0(byte_transmit_counter_c[5]), .I1(n3840), 
            .CO(n36491));
    SB_LUT4 i6_4_lut_adj_903 (.I0(\data_in_frame[12] [7]), .I1(n12_adj_3162), 
            .I2(\data_in_frame[19] [4]), .I3(n43090), .O(n42951));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 equal_1045_i7_2_lut (.I0(Kp_23__N_458), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/coms.v(225[9:81])
    defparam equal_1045_i7_2_lut.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n24383));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n7_adj_3163), .S(n8_adj_3164));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10776_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[12]), .I3(\data_out_frame[16] [4]), .O(n24194));
    defparam i10776_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_564_6_lut (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter_c[4]), 
            .I2(n3840), .I3(n36489), .O(n23898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_564_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_904 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43084));
    defparam i1_2_lut_adj_904.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_905 (.I0(\data_in_frame[1] [3]), .I1(n43274), .I2(GND_net), 
            .I3(GND_net), .O(n22770));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_adj_905.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_906 (.I0(n43084), .I1(n43256), .I2(\data_in_frame[11] [7]), 
            .I3(n42755), .O(n12_adj_3165));
    defparam i5_4_lut_adj_906.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_907 (.I0(\data_in_frame[7] [6]), .I1(n12_adj_3165), 
            .I2(n43319), .I3(n22770), .O(n39692));
    defparam i6_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_908 (.I0(\data_in_frame[12] [2]), .I1(n22977), 
            .I2(GND_net), .I3(GND_net), .O(n43298));
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_7__7__I_0_2_lut (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_515));   // verilog/coms.v(82[17:28])
    defparam data_in_frame_7__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_909 (.I0(\data_in_frame[14] [2]), .I1(n39692), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n43030));
    defparam i2_3_lut_adj_909.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_910 (.I0(n43077), .I1(\data_in_frame[12] [0]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n43244));
    defparam i2_3_lut_adj_910.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_911 (.I0(n22826), .I1(n43262), .I2(Kp_23__N_515), 
            .I3(\data_in_frame[10] [1]), .O(n12_adj_3166));
    defparam i5_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n42088), .S(n42004));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n42084), .S(n41998));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n42200), .S(n41892));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n7_adj_3167), .S(n8_adj_3168));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n7_adj_3169), .S(n28539));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n42136), .S(n28932));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n7_adj_3170), .S(n8_adj_3171));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n7_adj_3172), .S(n8_adj_3173));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n42124), .S(n41966));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n42122), .S(n42008));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n7_adj_3174), .S(n8_adj_3175));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n42120), .S(n42010));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n28495), .S(n8_adj_3176));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n42118), .S(n42012));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n7_adj_3177), .S(n8_adj_3178));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n42116), .S(n42014));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n42114), .S(n42016));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n42112), .S(n42018));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n42110), .S(n42020));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n42108), .S(n42022));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n42106), .S(n42024));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n42104), .S(n42026));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n42102), .S(n42028));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n42100), .S(n42030));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n42044), .S(n28920));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n28493), .S(n28918));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n42098), .S(n41958));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk32MHz), 
            .D(n41956), .S(n42198));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
            .D(n41946), .S(n49489));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n24050));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i6_4_lut_adj_912 (.I0(n39692), .I1(n12_adj_3166), .I2(\data_in_frame[14] [3]), 
            .I3(n43081), .O(n44318));
    defparam i6_4_lut_adj_912.LUT_INIT = 16'h6996;
    SB_LUT4 i10777_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[11]), .I3(\data_out_frame[16] [3]), .O(n24195));
    defparam i10777_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_913 (.I0(n44318), .I1(n43244), .I2(n43030), .I3(n38953), 
            .O(n23017));
    defparam i3_4_lut_adj_913.LUT_INIT = 16'h9669;
    SB_LUT4 i10778_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[10]), .I3(\data_out_frame[16] [2]), .O(n24196));
    defparam i10778_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_914 (.I0(\data_in_frame[16] [4]), .I1(n23017), 
            .I2(GND_net), .I3(GND_net), .O(n39049));
    defparam i1_2_lut_adj_914.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n24049));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n24048));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n24047));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n24046));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n24045));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10779_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[9]), .I3(\data_out_frame[16] [1]), .O(n24197));
    defparam i10779_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n24044));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n24043));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n24042));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n24041));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n24040));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n24039));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n24038));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22]_c [7]), .C(clk32MHz), 
            .E(n23610), .D(n44064));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i3_4_lut_adj_915 (.I0(\data_in_frame[4] [3]), .I1(n42769), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[2] [1]), .O(n22853));   // verilog/coms.v(225[9:81])
    defparam i3_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i10780_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[8]), .I3(\data_out_frame[16] [0]), .O(n24198));
    defparam i10780_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_916 (.I0(\data_in_frame[4] [7]), .I1(n39661), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_3179));
    defparam i1_2_lut_adj_916.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_917 (.I0(n43033), .I1(\data_in_frame[9] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3180));
    defparam i2_2_lut_adj_917.LUT_INIT = 16'h6666;
    SB_CARRY add_564_6 (.CI(n36489), .I0(byte_transmit_counter_c[4]), .I1(n3840), 
            .CO(n36490));
    SB_LUT4 i6_4_lut_adj_918 (.I0(n16_adj_3179), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[7] [1]), .I3(\data_in_frame[8] [7]), .O(n14_adj_3181));
    defparam i6_4_lut_adj_918.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_919 (.I0(\data_in_frame[11] [3]), .I1(n14_adj_3181), 
            .I2(n10_adj_3180), .I3(n22853), .O(n43834));
    defparam i7_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_920 (.I0(n43834), .I1(n42984), .I2(GND_net), 
            .I3(GND_net), .O(n23038));
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h9999;
    SB_LUT4 i10781_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[23]), .I3(\data_out_frame[15] [7]), .O(n24199));
    defparam i10781_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22]_c [6]), .C(clk32MHz), 
            .E(n23610), .D(n42924));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22]_c [5]), .C(clk32MHz), 
            .E(n23610), .D(n23309));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_adj_921 (.I0(n43286), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[16] [1]), .I3(GND_net), .O(n43234));   // verilog/coms.v(71[16:43])
    defparam i2_3_lut_adj_921.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_922 (.I0(n23113), .I1(n23038), .I2(\data_in_frame[13] [5]), 
            .I3(n6_adj_3182), .O(n39672));
    defparam i4_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22]_c [4]), .C(clk32MHz), 
            .E(n23610), .D(n22958));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22]_c [3]), .C(clk32MHz), 
            .E(n23610), .D(n42897));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22]_c [2]), .C(clk32MHz), 
            .E(n23610), .D(n43063));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22]_c [0]), .C(clk32MHz), 
            .E(n23610), .D(n23311));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n23610), .D(n43849));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n23610), .D(n44248));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n23610), .D(n44212));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n23610), .D(n44323));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n23610), .D(n43950));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n23610), .D(n43632));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n23610), .D(n44218));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n23610), .D(n44444));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n24037));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i3_4_lut_adj_923 (.I0(\data_in_frame[4] [2]), .I1(n42849), .I2(\data_in_frame[0] [0]), 
            .I3(\data_in_frame[1] [6]), .O(n23229));   // verilog/coms.v(67[16:27])
    defparam i3_4_lut_adj_923.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_924 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[6] [7]), 
            .I2(\data_in_frame[11] [2]), .I3(n23229), .O(n42999));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_924.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_925 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n22750));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_adj_925.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_926 (.I0(n43259), .I1(\data_in_frame[4] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3183));
    defparam i2_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[9] [4]), 
            .I2(n6_adj_3183), .I3(n43074), .O(n43077));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i10782_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[22]), .I3(\data_out_frame[15] [6]), .O(n24200));
    defparam i10782_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_927 (.I0(\data_in_frame[7] [3]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43319));
    defparam i1_2_lut_adj_927.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_928 (.I0(n42877), .I1(n43162), .I2(\data_in_frame[5] [3]), 
            .I3(GND_net), .O(n23032));   // verilog/coms.v(82[17:28])
    defparam i2_3_lut_adj_928.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_929 (.I0(n39661), .I1(n39331), .I2(\data_in_frame[4] [7]), 
            .I3(GND_net), .O(n43256));
    defparam i2_3_lut_adj_929.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_930 (.I0(\data_in_frame[7] [3]), .I1(n22977), .I2(n39675), 
            .I3(\data_in_frame[5] [0]), .O(n43259));
    defparam i3_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_931 (.I0(\data_in_frame[7] [1]), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43056));
    defparam i1_2_lut_adj_931.LUT_INIT = 16'h6666;
    SB_LUT4 i10784_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[20]), .I3(\data_out_frame[15] [4]), .O(n24202));
    defparam i10784_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_4_lut_adj_932 (.I0(\data_in_frame[11] [5]), .I1(n22858), 
            .I2(n8_adj_3184), .I3(n43247), .O(n43310));
    defparam i1_4_lut_adj_932.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_933 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42755));
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_934 (.I0(\data_in_frame[5] [2]), .I1(n23528), .I2(n4_c), 
            .I3(\data_in_frame[3] [1]), .O(n22977));
    defparam i1_4_lut_adj_934.LUT_INIT = 16'h6996;
    SB_LUT4 i10785_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[19]), .I3(\data_out_frame[15] [3]), .O(n24203));
    defparam i10785_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n24036));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_564_5_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[3]), 
            .I2(n3840), .I3(n36488), .O(n23895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_564_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i4_4_lut_adj_935 (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[3] [2]), 
            .I2(n42821), .I3(n6_adj_3185), .O(n5_adj_3186));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_936 (.I0(n43050), .I1(n43256), .I2(n23032), .I3(GND_net), 
            .O(n39619));
    defparam i2_3_lut_adj_936.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_937 (.I0(n39619), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[14] [1]), .I3(GND_net), .O(n43231));
    defparam i2_3_lut_adj_937.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_938 (.I0(n5_adj_3186), .I1(n43081), .I2(n22977), 
            .I3(GND_net), .O(n38953));
    defparam i2_3_lut_adj_938.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_939 (.I0(\data_in_frame[14] [0]), .I1(n43310), 
            .I2(GND_net), .I3(GND_net), .O(n43014));
    defparam i1_2_lut_adj_939.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_940 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n4_c));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_940.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_941 (.I0(\data_in_frame[5] [0]), .I1(n39675), .I2(GND_net), 
            .I3(GND_net), .O(n22979));
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_942 (.I0(\data_in_frame[6] [7]), .I1(n22979), .I2(\data_in_frame[6] [6]), 
            .I3(\data_in_frame[9] [2]), .O(n43033));
    defparam i3_4_lut_adj_942.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_943 (.I0(n39661), .I1(n43053), .I2(GND_net), 
            .I3(GND_net), .O(n43054));
    defparam i1_2_lut_adj_943.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_944 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42821));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_945 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n42829));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_945.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_946 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42849));   // verilog/coms.v(67[16:27])
    defparam i1_2_lut_adj_946.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_947 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43162));   // verilog/coms.v(82[17:28])
    defparam i1_2_lut_adj_947.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_948 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42832));   // verilog/coms.v(68[16:69])
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_949 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42817));   // verilog/coms.v(225[9:81])
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_950 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [6]), 
            .I2(n42817), .I3(n6_adj_3187), .O(Kp_23__N_290));   // verilog/coms.v(70[16:34])
    defparam i4_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_951 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(Kp_23__N_290), .I3(\data_in_frame[1] [0]), .O(n43145));   // verilog/coms.v(67[16:69])
    defparam i3_4_lut_adj_951.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_952 (.I0(n43145), .I1(Kp_23__N_290), .I2(n21084), 
            .I3(\data_in_frame[0] [7]), .O(n42877));   // verilog/coms.v(68[16:69])
    defparam i3_4_lut_adj_952.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_953 (.I0(\data_in_frame[3] [7]), .I1(n43145), .I2(\data_in_frame[0] [3]), 
            .I3(\data_in_frame[2] [6]), .O(n18));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n42832), .I1(n18), .I2(n43162), .I3(Kp_23__N_325), 
            .O(n20));   // verilog/coms.v(75[16:27])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_954 (.I0(n42772), .I1(Kp_23__N_319), .I2(n42849), 
            .I3(\data_in_frame[1] [5]), .O(n19_adj_3188));   // verilog/coms.v(75[16:27])
    defparam i8_4_lut_adj_954.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(n43117), .I1(n42829), .I2(n19_adj_3188), .I3(n20), 
            .O(n38906));   // verilog/coms.v(70[16:34])
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_955 (.I0(n38906), .I1(n42877), .I2(\data_in_frame[5] [1]), 
            .I3(GND_net), .O(n39331));
    defparam i2_3_lut_adj_955.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3189), .S(n3_adj_3124));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_adj_956 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42772));   // verilog/coms.v(161[9:87])
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42769));   // verilog/coms.v(161[9:87])
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_958 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n23446));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_958.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_959 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n5_adj_3190));   // verilog/coms.v(161[9:87])
    defparam i2_3_lut_adj_959.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_960 (.I0(n5_adj_3190), .I1(n23446), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_325));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h6666;
    SB_LUT4 equal_1045_i13_2_lut (.I0(Kp_23__N_319), .I1(\data_in_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n23233));   // verilog/coms.v(225[9:81])
    defparam equal_1045_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10786_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[18]), .I3(\data_out_frame[15] [2]), .O(n24204));
    defparam i10786_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_961 (.I0(n39331), .I1(\data_in_frame[9] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n43247));
    defparam i1_2_lut_adj_961.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_838));   // verilog/coms.v(67[16:27])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_962 (.I0(n39661), .I1(n43247), .I2(n23233), .I3(n23164), 
            .O(n12_adj_3191));
    defparam i5_4_lut_adj_962.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_963 (.I0(n43054), .I1(n12_adj_3191), .I2(\data_in_frame[11] [4]), 
            .I3(n43033), .O(n42984));
    defparam i6_4_lut_adj_963.LUT_INIT = 16'h9669;
    SB_LUT4 i10787_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[17]), .I3(\data_out_frame[15] [1]), .O(n24205));
    defparam i10787_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10788_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[16]), .I3(\data_out_frame[15] [0]), .O(n24206));
    defparam i10788_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10789_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[7]), .I3(\data_out_frame[14] [7]), .O(n24207));
    defparam i10789_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_964 (.I0(n42984), .I1(Kp_23__N_838), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3192));
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_965 (.I0(n43014), .I1(n38953), .I2(\data_in_frame[12] [0]), 
            .I3(n43231), .O(n10_adj_3193));
    defparam i4_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_966 (.I0(\data_in_frame[11] [7]), .I1(n10_adj_3193), 
            .I2(n23113), .I3(n4_adj_3192), .O(n39257));
    defparam i5_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_967 (.I0(n23519), .I1(\data_in_frame[9] [0]), .I2(\data_in_frame[6] [6]), 
            .I3(n6_adj_3194), .O(n22885));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_967.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_968 (.I0(n23113), .I1(n43148), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3195));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_969 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[16] [0]), 
            .I2(n22885), .I3(n6_adj_3195), .O(n43286));
    defparam i4_4_lut_adj_969.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\data_in_frame[16] [2]), .I1(n39257), 
            .I2(GND_net), .I3(GND_net), .O(n39648));
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_971 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3196));
    defparam i6_4_lut_adj_971.LUT_INIT = 16'h8000;
    SB_LUT4 i10790_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[6]), .I3(\data_out_frame[14] [6]), .O(n24208));
    defparam i10790_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i6_4_lut_adj_972 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3197));   // verilog/coms.v(227[13:35])
    defparam i6_4_lut_adj_972.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_973 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13));
    defparam i5_4_lut_adj_973.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_974 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_adj_3198));   // verilog/coms.v(227[13:35])
    defparam i5_4_lut_adj_974.LUT_INIT = 16'hfffe;
    SB_LUT4 i15076_4_lut (.I0(n13_adj_3198), .I1(n13), .I2(n14_adj_3197), 
            .I3(n14_adj_3196), .O(n28473));
    defparam i15076_4_lut.LUT_INIT = 16'h32fa;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[17] [7]), .I1(n39672), .I2(n43234), 
            .I3(GND_net), .O(n8_adj_3199));
    defparam i3_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_975 (.I0(n42951), .I1(n43196), .I2(\data_in_frame[21] [5]), 
            .I3(GND_net), .O(n44463));
    defparam i2_3_lut_adj_975.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_976 (.I0(n39648), .I1(\data_in_frame[20] [4]), 
            .I2(\data_in_frame[18] [3]), .I3(n43286), .O(n10_adj_3200));
    defparam i4_4_lut_adj_976.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_977 (.I0(\data_in_frame[18] [4]), .I1(n43064), 
            .I2(\data_in_frame[20] [6]), .I3(n39049), .O(n43842));
    defparam i3_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_978 (.I0(n23513), .I1(\data_in_frame[19] [0]), 
            .I2(n43139), .I3(n23470), .O(n8_adj_3201));   // verilog/coms.v(72[16:43])
    defparam i2_4_lut_adj_978.LUT_INIT = 16'h6996;
    SB_LUT4 i4_3_lut_adj_979 (.I0(n42919), .I1(n8_adj_3201), .I2(\data_in_frame[18] [5]), 
            .I3(GND_net), .O(n10_adj_3202));   // verilog/coms.v(72[16:43])
    defparam i4_3_lut_adj_979.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3203), .S(n3_adj_3123));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3204), .S(n3_adj_3122));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3205), .S(n3_adj_3121));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3206), .S(n3_adj_3120));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3207), .S(n3_adj_3119));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3208), .S(n3_adj_3118));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3209), .S(n3_adj_3117));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_3210), .S(n3_adj_3116));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_3211), .S(n3_adj_3115));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_3212), .S(n3_adj_3114));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_3213), .S(n3_adj_3113));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3214), .S(n3_adj_3112));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3215), .S(n3_adj_3111));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_3127), .S(n3_adj_3110));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3128), .S(n3_c));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3130), .S(n3_adj_3216));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3136), .S(n3_adj_3217));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3138), .S(n3_adj_3218));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3139), .S(n3_adj_3219));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3140), .S(n3_adj_3220));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3146), .S(n3_adj_3221));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3222), .S(n3_adj_3223));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3224), .S(n3_adj_3225));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3226), .S(n3_adj_3227));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3228), .S(n3_adj_3229));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_3230));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3129), .S(n3_adj_3231));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3137), .S(n3_adj_3232));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3145), .S(n3_adj_3233));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3234), .S(n3_adj_3235));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n24035));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_adj_980 (.I0(n43026), .I1(n43241), .I2(\data_in_frame[21] [3]), 
            .I3(GND_net), .O(n43618));
    defparam i2_3_lut_adj_980.LUT_INIT = 16'h9696;
    SB_LUT4 i10855_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[21]), .I3(\data_out_frame[6] [5]), .O(n24273));
    defparam i10855_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_981 (.I0(n22801), .I1(\data_in_frame[19] [0]), 
            .I2(n39049), .I3(n43026), .O(n10_adj_3236));
    defparam i4_4_lut_adj_981.LUT_INIT = 16'h6996;
    SB_CARRY add_564_5 (.CI(n36488), .I0(byte_transmit_counter_c[3]), .I1(n3840), 
            .CO(n36489));
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n24034));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n24033));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_12 (.CI(n36464), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n36465));
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n24032));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n24031));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_564_4_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter_c[2]), 
            .I2(n3840), .I3(n36487), .O(n23892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_564_4_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_564_4 (.CI(n36487), .I0(byte_transmit_counter_c[2]), .I1(n3840), 
            .CO(n36488));
    SB_LUT4 add_41_3_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n36455), .O(n2_adj_3234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_982 (.I0(\data_in_frame[20] [1]), .I1(n43071), 
            .I2(\data_in_frame[17] [7]), .I3(GND_net), .O(n43891));
    defparam i2_3_lut_adj_982.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33878 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter_c[1]), .O(n49396));
    defparam byte_transmit_counter_0__bdd_4_lut_33878.LUT_INIT = 16'he4aa;
    SB_LUT4 i29085_4_lut (.I0(Kp_23__N_785), .I1(n43891), .I2(n10_adj_3236), 
            .I3(\data_in_frame[21] [2]), .O(n44596));
    defparam i29085_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 add_41_11_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n36463), .O(n2_adj_3222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_3 (.CI(n36455), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n36456));
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n24030));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10791_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[5]), .I3(\data_out_frame[14] [5]), .O(n24209));
    defparam i10791_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_564_3_lut (.I0(byte_transmit_counter_c[1]), .I1(byte_transmit_counter_c[1]), 
            .I2(n3840), .I3(n36486), .O(n23889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_564_3_lut.LUT_INIT = 16'hA3AC;
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n24029));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_564_3 (.CI(n36486), .I0(byte_transmit_counter_c[1]), .I1(n3840), 
            .CO(n36487));
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n24028));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n24027));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n24026));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_4_lut_adj_983 (.I0(n39672), .I1(n43842), .I2(n10_adj_3200), 
            .I3(\data_in_frame[18] [2]), .O(n10_adj_3237));
    defparam i2_4_lut_adj_983.LUT_INIT = 16'hedde;
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n24025));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10792_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[4]), .I3(\data_out_frame[14] [4]), .O(n24210));
    defparam i10792_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10793_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[3]), .I3(\data_out_frame[14] [3]), .O(n24211));
    defparam i10793_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_984 (.I0(\data_in_frame[16] [5]), .I1(n43618), 
            .I2(n10_adj_3202), .I3(\data_in_frame[20] [7]), .O(n11));
    defparam i3_4_lut_adj_984.LUT_INIT = 16'hdeed;
    SB_LUT4 add_564_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_2639), .I3(GND_net), .O(n2241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_564_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10794_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[2]), .I3(\data_out_frame[14] [2]), .O(n24212));
    defparam i10794_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_4_lut_adj_985 (.I0(\data_in_frame[20] [3]), .I1(n44463), 
            .I2(n8_adj_3199), .I3(n43017), .O(n9));
    defparam i1_4_lut_adj_985.LUT_INIT = 16'hdeed;
    SB_LUT4 i1_rep_20_2_lut (.I0(\data_in_frame[19] [0]), .I1(n23470), .I2(GND_net), 
            .I3(GND_net), .O(n49513));   // verilog/coms.v(72[16:43])
    defparam i1_rep_20_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10795_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[1]), .I3(\data_out_frame[14] [1]), .O(n24213));
    defparam i10795_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i5_4_lut_adj_986 (.I0(n43139), .I1(n49513), .I2(\data_in_frame[21] [0]), 
            .I3(\data_in_frame[16] [7]), .O(n12_adj_3238));
    defparam i5_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_CARRY add_564_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_2639), 
            .CO(n36486));
    SB_LUT4 i10796_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[0]), .I3(\data_out_frame[14] [0]), .O(n24214));
    defparam i10796_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n24024));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n24023));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n24022));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n24021));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n24020));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n24019));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n24018));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n24017));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n24016));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n24015));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i5_4_lut_adj_987 (.I0(n23513), .I1(n23026), .I2(n43142), .I3(n39049), 
            .O(n12_adj_3239));
    defparam i5_4_lut_adj_987.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n24014));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n24013));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n24012));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n24011));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n24010));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49396_bdd_4_lut (.I0(n49396), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter_c[1]), 
            .O(n49399));
    defparam n49396_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_41_33_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n36485), .O(n2_adj_3189)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_988 (.I0(n23467), .I1(\data_in_frame[20] [2]), 
            .I2(n43017), .I3(n6_adj_3240), .O(n43615));
    defparam i4_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 i10797_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[15]), .I3(\data_out_frame[13] [7]), .O(n24215));
    defparam i10797_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_41_32_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n36484), .O(n2_adj_3203)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_989 (.I0(n22682), .I1(\data_in_frame[20] [5]), 
            .I2(\data_in_frame[18] [3]), .I3(\data_in_frame[18] [4]), .O(n8_adj_3241));
    defparam i3_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_990 (.I0(n9), .I1(n11), .I2(n10_adj_3237), .I3(n44596), 
            .O(n44547));
    defparam i7_4_lut_adj_990.LUT_INIT = 16'hfeff;
    SB_CARRY add_41_32 (.CI(n36484), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n36485));
    SB_LUT4 add_41_31_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n36483), .O(n2_adj_3204)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_991 (.I0(n39629), .I1(n12_adj_3238), .I2(n43313), 
            .I3(\data_in_frame[16] [3]), .O(n43841));
    defparam i6_4_lut_adj_991.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_992 (.I0(n42904), .I1(n42951), .I2(\data_in_frame[21] [6]), 
            .I3(GND_net), .O(n44167));
    defparam i2_3_lut_adj_992.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_993 (.I0(n42902), .I1(n39672), .I2(n8_adj_3241), 
            .I3(n39629), .O(n13_adj_3242));
    defparam i4_4_lut_adj_993.LUT_INIT = 16'h7dd7;
    SB_CARRY add_41_31 (.CI(n36483), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n36484));
    SB_LUT4 add_41_30_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n36482), .O(n2_adj_3205)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10798_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[14]), .I3(\data_out_frame[13] [6]), .O(n24216));
    defparam i10798_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n24009));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n24008));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n24007));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n24006));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n24005));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i6_4_lut_adj_994 (.I0(\data_in_frame[16] [3]), .I1(n12_adj_3239), 
            .I2(n23470), .I3(\data_in_frame[21] [1]), .O(n44377));
    defparam i6_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n24004));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n24003));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i3_4_lut_adj_995 (.I0(\data_in_frame[21] [4]), .I1(n43615), 
            .I2(n43196), .I3(n43241), .O(n12_adj_3243));
    defparam i3_4_lut_adj_995.LUT_INIT = 16'hedde;
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n24002));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n24001));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i7_4_lut_adj_996 (.I0(n13_adj_3242), .I1(n44167), .I2(n43841), 
            .I3(n44547), .O(n16_adj_3244));
    defparam i7_4_lut_adj_996.LUT_INIT = 16'hffbf;
    SB_LUT4 i10799_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[13]), .I3(\data_out_frame[13] [5]), .O(n24217));
    defparam i10799_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n24000));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n23999));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10848_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[12]), .I3(\data_out_frame[7] [4]), .O(n24266));
    defparam i10848_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_997 (.I0(\data_in_frame[20] [0]), .I1(n43238), 
            .I2(n43172), .I3(n43071), .O(n43617));
    defparam i3_4_lut_adj_997.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_998 (.I0(n43617), .I1(n16_adj_3244), .I2(n12_adj_3243), 
            .I3(n44377), .O(n31));
    defparam i8_4_lut_adj_998.LUT_INIT = 16'hfeff;
    SB_CARRY add_41_30 (.CI(n36482), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n36483));
    SB_LUT4 i10833_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[19]), .I3(\data_out_frame[9] [3]), .O(n24251));
    defparam i10833_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10831_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[21]), .I3(\data_out_frame[9] [5]), .O(n24249));
    defparam i10831_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10863_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(control_mode[5]), .I3(\data_out_frame[5] [5]), .O(n24281));
    defparam i10863_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10862_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(control_mode[6]), .I3(\data_out_frame[5] [6]), .O(n24280));
    defparam i10862_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10822_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[14]), .I3(\data_out_frame[10] [6]), .O(n24240));
    defparam i10822_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15097_2_lut (.I0(n31), .I1(n28473), .I2(GND_net), .I3(GND_net), 
            .O(n28496));
    defparam i15097_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10850_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[10]), .I3(\data_out_frame[7] [2]), .O(n24268));
    defparam i10850_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_41_29_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n36481), .O(n2_adj_3206)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_29_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n23998));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n23997));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n23996));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n23995));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n23994));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n23993));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n23992));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n23991));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_29 (.CI(n36481), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n36482));
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n23990));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n23989));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n23988));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n23987));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n23986));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n23985));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n23984));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n23983));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n23982));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n23981));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n23980));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n23979));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n23978));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n23977));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n23976));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i1 (.Q(\PWMLimit[1] ), .C(clk32MHz), .D(n23975));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i2 (.Q(\PWMLimit[2] ), .C(clk32MHz), .D(n23974));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i3 (.Q(\PWMLimit[3] ), .C(clk32MHz), .D(n23973));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i4 (.Q(\PWMLimit[4] ), .C(clk32MHz), .D(n23972));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i5 (.Q(\PWMLimit[5] ), .C(clk32MHz), .D(n23971));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i6 (.Q(\PWMLimit[6] ), .C(clk32MHz), .D(n23970));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i7 (.Q(\PWMLimit[7] ), .C(clk32MHz), .D(n28310));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i8 (.Q(\PWMLimit[8] ), .C(clk32MHz), .D(n23968));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i9 (.Q(\PWMLimit[9] ), .C(clk32MHz), .D(n23967));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10852_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[8]), .I3(\data_out_frame[7] [0]), .O(n24270));
    defparam i10852_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY add_41_11 (.CI(n36463), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n36464));
    SB_LUT4 i10853_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[23]), .I3(\data_out_frame[6] [7]), .O(n24271));
    defparam i10853_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state[2] ), .C(clk32MHz), 
           .D(n49493));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_28_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n36480), .O(n2_adj_3207)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_41_2_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2_adj_3245)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_41_10_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n36462), .O(n2_adj_3224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_28 (.CI(n36480), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n36481));
    SB_LUT4 add_41_27_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n36479), .O(n2_adj_3208)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_27 (.CI(n36479), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n36480));
    SB_CARRY add_41_10 (.CI(n36462), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n36463));
    SB_LUT4 i10774_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[14]), .I3(\data_out_frame[16] [6]), .O(n24192));
    defparam i10774_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_41_26_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n36478), .O(n2_adj_3209)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n36455));
    SB_CARRY add_41_26 (.CI(n36478), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n36479));
    SB_LUT4 add_41_9_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n36461), .O(n2_adj_3226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10821_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[15]), .I3(\data_out_frame[10] [7]), .O(n24239));
    defparam i10821_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY add_41_9 (.CI(n36461), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n36462));
    SB_LUT4 i10818_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder1_position[2]), .I3(\data_out_frame[11] [2]), .O(n24236));
    defparam i10818_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10809_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[19]), .I3(\data_out_frame[12] [3]), .O(n24227));
    defparam i10809_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10772_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[0]), .I3(\data_out_frame[17] [0]), .O(n24190));
    defparam i10772_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10768_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(pwm[4]), .I3(\data_out_frame[17] [4]), .O(n24186));
    defparam i10768_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10851_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(encoder0_position[9]), .I3(\data_out_frame[7] [1]), .O(n24269));
    defparam i10851_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_41_25_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n36477), .O(n2_adj_3210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_25 (.CI(n36477), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n36478));
    SB_LUT4 i10746_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[2]), .I3(\data_out_frame[20] [2]), .O(n24164));
    defparam i10746_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10800_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(setpoint[12]), .I3(\data_out_frame[13] [4]), .O(n24218));
    defparam i10800_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10755_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22498), 
            .I2(displacement[9]), .I3(\data_out_frame[19] [1]), .O(n24173));
    defparam i10755_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n24358));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n24357));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n24356));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n24355));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n24310));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33873 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n49384));
    defparam byte_transmit_counter_0__bdd_4_lut_33873.LUT_INIT = 16'he4aa;
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n24309));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n24354));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_4_lut_adj_999 (.I0(n5025), .I1(n28895), .I2(\FRAME_MATCHER.state_31__N_1924 [3]), 
            .I3(n5023), .O(n23616));
    defparam i1_4_lut_adj_999.LUT_INIT = 16'ha022;
    SB_LUT4 add_41_24_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n36476), .O(n2_adj_3211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_24_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n24308));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2054_2_lut (.I0(n3362), .I1(\FRAME_MATCHER.state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n5023));
    defparam i2054_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n24307));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n24353));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), .C(clk32MHz), 
           .D(n23897));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n49384_bdd_4_lut (.I0(n49384), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n49387));
    defparam n49384_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_41_24 (.CI(n36476), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n36477));
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), .C(clk32MHz), 
           .D(n23900));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), .C(clk32MHz), 
           .D(n23903));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), .C(clk32MHz), 
           .D(n23906));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), .C(clk32MHz), 
           .D(n23909));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSR tx_transmit_3220 (.Q(r_SM_Main_2__N_2747[0]), .C(clk32MHz), 
            .D(n46678), .R(n43341));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n24352));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_23_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n36475), .O(n2_adj_3212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_23 (.CI(n36475), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n36476));
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n24351));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kd_i1 (.Q(\Kd[1] ), .C(clk32MHz), .D(n24350));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kd_i2 (.Q(\Kd[2] ), .C(clk32MHz), .D(n24349));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n24382));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i6_4_lut_adj_1000 (.I0(\FRAME_MATCHER.state [10]), .I1(\FRAME_MATCHER.state [11]), 
            .I2(\FRAME_MATCHER.state [8]), .I3(\FRAME_MATCHER.state [15]), 
            .O(n14_adj_3246));
    defparam i6_4_lut_adj_1000.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33864 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter_c[1]), .O(n49378));
    defparam byte_transmit_counter_0__bdd_4_lut_33864.LUT_INIT = 16'he4aa;
    SB_LUT4 n49378_bdd_4_lut (.I0(n49378), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n49381));
    defparam n49378_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_41_22_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n36474), .O(n2_adj_3213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_4_lut_adj_1001 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(\FRAME_MATCHER.state [12]), .I3(\FRAME_MATCHER.state [9]), 
            .O(n13_adj_3247));
    defparam i5_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(n13_adj_3247), .I1(\FRAME_MATCHER.state [7]), 
            .I2(n14_adj_3246), .I3(GND_net), .O(n6_adj_3248));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1002 (.I0(\FRAME_MATCHER.state [5]), .I1(\FRAME_MATCHER.state [6]), 
            .I2(\FRAME_MATCHER.state [4]), .I3(n6_adj_3248), .O(n42743));
    defparam i4_4_lut_adj_1002.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1003 (.I0(\FRAME_MATCHER.state [18]), .I1(\FRAME_MATCHER.state [27]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [16]), 
            .O(n12_adj_3249));
    defparam i5_4_lut_adj_1003.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1004 (.I0(\FRAME_MATCHER.state [20]), .I1(n12_adj_3249), 
            .I2(\FRAME_MATCHER.state [23]), .I3(\FRAME_MATCHER.state [24]), 
            .O(n39501));
    defparam i6_4_lut_adj_1004.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1005 (.I0(\FRAME_MATCHER.state [25]), .I1(\FRAME_MATCHER.state [17]), 
            .I2(\FRAME_MATCHER.state [26]), .I3(GND_net), .O(n14_adj_3250));
    defparam i5_3_lut_adj_1005.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1006 (.I0(\FRAME_MATCHER.state [29]), .I1(\FRAME_MATCHER.state [21]), 
            .I2(\FRAME_MATCHER.state [28]), .I3(\FRAME_MATCHER.state [30]), 
            .O(n15_adj_3251));
    defparam i6_4_lut_adj_1006.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1007 (.I0(n15_adj_3251), .I1(\FRAME_MATCHER.state [22]), 
            .I2(n14_adj_3250), .I3(\FRAME_MATCHER.state [19]), .O(n42612));
    defparam i8_4_lut_adj_1007.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n22513));   // verilog/coms.v(248[5:27])
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1009 (.I0(n42612), .I1(n39501), .I2(n42743), 
            .I3(GND_net), .O(n29039));
    defparam i2_3_lut_adj_1009.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1010 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n22492));
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'h2222;
    SB_LUT4 i15_rep_4_2_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n49497));
    defparam i15_rep_4_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1011 (.I0(n49497), .I1(n29039), .I2(n4_adj_3252), 
            .I3(n22513), .O(n3362));
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'h3032;
    SB_DFF Kd_i3 (.Q(\Kd[3] ), .C(clk32MHz), .D(n24348));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kd_i4 (.Q(\Kd[4] ), .C(clk32MHz), .D(n24347));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kd_i5 (.Q(\Kd[5] ), .C(clk32MHz), .D(n24346));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kd_i6 (.Q(\Kd[6] ), .C(clk32MHz), .D(n24345));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_8_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n36460), .O(n2_adj_3228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_22 (.CI(n36474), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n36475));
    SB_DFF deadband_i0_i0 (.Q(\deadband[0] ), .C(clk32MHz), .D(n23829));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n23828));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n24272));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_3245), .S(n3_adj_3253));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_21_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n36473), .O(n2_adj_3214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_21 (.CI(n36473), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n36474));
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n24381));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n24380));   // verilog/coms.v(125[12] 284[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n42006));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_20_lut (.I0(n1508), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n36472), .O(n2_adj_3215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_20_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i0 (.Q(\PWMLimit[0] ), .C(clk32MHz), .D(n23811));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n23810));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n23809));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n23808));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n23807));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kd_i0 (.Q(\Kd[0] ), .C(clk32MHz), .D(n23806));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n23805));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n23804));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n23803));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 mux_956_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[16] [0]), .O(n3800));
    defparam mux_956_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[16] [1]), .O(n3801));
    defparam mux_956_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[16] [2]), .O(n3802));
    defparam mux_956_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[16] [3]), .O(n3803));
    defparam mux_956_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[16] [4]), .O(n3804));
    defparam mux_956_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[16] [5]), .O(n3805));
    defparam mux_956_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[16] [6]), .O(n3806));
    defparam mux_956_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[16] [7]), .O(n3807));
    defparam mux_956_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[15] [0]), .O(n3808));
    defparam mux_956_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[15] [1]), .O(n3809));
    defparam mux_956_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[15] [2]), .O(n3810));
    defparam mux_956_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[15] [3]), .O(n3811));
    defparam mux_956_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[15] [4]), .O(n3812));
    defparam mux_956_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[15] [5]), .O(n3813));
    defparam mux_956_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[15] [6]), .O(n3814));
    defparam mux_956_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[15] [7]), .O(n3815));
    defparam mux_956_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[14] [0]), .O(n3816));
    defparam mux_956_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44681), .I3(n44680), 
            .O(tx_data[7]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44678), .I3(n44677), 
            .O(tx_data[6]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44675), .I3(n44674), 
            .O(tx_data[5]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 mux_956_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[14] [1]), .O(n3817));
    defparam mux_956_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[14] [2]), .O(n3818));
    defparam mux_956_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44672), .I3(n44671), 
            .O(tx_data[3]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 mux_956_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[14] [3]), .O(n3819));
    defparam mux_956_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[14] [4]), .O(n3820));
    defparam mux_956_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(byte_transmit_counter_c[2]), 
            .I1(n44739), .I2(n48097), .I3(byte_transmit_counter_c[3]), 
            .O(n49372));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44663), .I3(n44662), 
            .O(tx_data[0]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44666), .I3(n44665), 
            .O(tx_data[1]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 mux_956_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[14] [5]), .O(n3821));
    defparam mux_956_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[14] [7]), .O(n3823));
    defparam mux_956_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_956_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n28475), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[14] [6]), .O(n3822));
    defparam mux_956_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n44669), .I3(n44668), 
            .O(tx_data[2]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 n49372_bdd_4_lut (.I0(n49372), .I1(n44689), .I2(n44688), .I3(byte_transmit_counter_c[3]), 
            .O(n49375));
    defparam n49372_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i29176_3_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter_c[1]), .I3(GND_net), .O(n44688));
    defparam i29176_3_lut.LUT_INIT = 16'hc2c2;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3254));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29177_4_lut (.I0(\data_out_frame[5] [4]), .I1(n5_adj_3254), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n44689));
    defparam i29177_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33859 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n49366));
    defparam byte_transmit_counter_0__bdd_4_lut_33859.LUT_INIT = 16'he4aa;
    SB_LUT4 n49366_bdd_4_lut (.I0(n49366), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n49369));
    defparam n49366_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15492_4_lut (.I0(n28473), .I1(n31), .I2(n31_adj_3255), .I3(\FRAME_MATCHER.state [1]), 
            .O(n28895));
    defparam i15492_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33850 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n49360));
    defparam byte_transmit_counter_0__bdd_4_lut_33850.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_3_lut_adj_1012 (.I0(n28895), .I1(n19960), .I2(n29039), 
            .I3(GND_net), .O(n44107));
    defparam i3_3_lut_adj_1012.LUT_INIT = 16'hfbfb;
    SB_LUT4 i12_4_lut (.I0(n16_adj_3179), .I1(n15_adj_3256), .I2(n22979), 
            .I3(n22770), .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i10_4_lut (.I0(n23229), .I1(n22853), .I2(n5_adj_3186), .I3(n23233), 
            .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n23032), .I1(n39331), .I2(n23449), .I3(n22977), 
            .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i9_4_lut_adj_1013 (.I0(n23347), .I1(n22858), .I2(n7), .I3(n10_adj_3157), 
            .O(n25));
    defparam i9_4_lut_adj_1013.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n31_adj_3255));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15078_2_lut (.I0(n31_adj_3255), .I1(n28473), .I2(GND_net), 
            .I3(GND_net), .O(n28475));
    defparam i15078_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1014 (.I0(n20014), .I1(n28496), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state[2] ), .O(n6_adj_3257));
    defparam i2_4_lut_adj_1014.LUT_INIT = 16'h5d55;
    SB_LUT4 i3_4_lut_adj_1015 (.I0(n29039), .I1(n6_adj_3257), .I2(n28475), 
            .I3(n22492), .O(n3840));
    defparam i3_4_lut_adj_1015.LUT_INIT = 16'hfeee;
    SB_LUT4 i15281_3_lut (.I0(n3840), .I1(\FRAME_MATCHER.state[0] ), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n28694));
    defparam i15281_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 mux_616_i1_4_lut (.I0(n28496), .I1(n29029), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n29035));   // verilog/coms.v(143[4] 283[11])
    defparam mux_616_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i31166_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n29035), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(n4_adj_3258), .O(n46678));   // verilog/coms.v(143[4] 283[11])
    defparam i31166_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3259));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31494_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n47008));   // verilog/coms.v(103[34:55])
    defparam i31494_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3260));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29147_4_lut (.I0(n19_adj_3259), .I1(\data_out_frame[22]_c [7]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n44659));
    defparam i29147_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29148_3_lut (.I0(n49363), .I1(n44659), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44660));
    defparam i29148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29167_4_lut (.I0(n5_adj_3260), .I1(n47008), .I2(n46420), 
            .I3(byte_transmit_counter[0]), .O(n44679));
    defparam i29167_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i29169_4_lut (.I0(n44679), .I1(n44660), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44681));
    defparam i29169_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29168_3_lut (.I0(n49429), .I1(n49423), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44680));
    defparam i29168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3261));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31487_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n47001));   // verilog/coms.v(103[34:55])
    defparam i31487_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3262));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29144_4_lut (.I0(n19_adj_3261), .I1(\data_out_frame[22]_c [6]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n44656));
    defparam i29144_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29145_3_lut (.I0(n49357), .I1(n44656), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44657));
    defparam i29145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29164_4_lut (.I0(n5_adj_3262), .I1(n47001), .I2(n46420), 
            .I3(byte_transmit_counter[0]), .O(n44676));
    defparam i29164_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i29166_4_lut (.I0(n44676), .I1(n44657), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44678));
    defparam i29166_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29165_3_lut (.I0(n49333), .I1(n49435), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44677));
    defparam i29165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3263));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter_c[1]), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n46994));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3264));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29141_4_lut (.I0(n19_adj_3263), .I1(\data_out_frame[22]_c [5]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n44653));
    defparam i29141_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29142_3_lut (.I0(n49351), .I1(n44653), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44654));
    defparam i29142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29161_4_lut (.I0(n5_adj_3264), .I1(byte_transmit_counter[0]), 
            .I2(n46420), .I3(n46994), .O(n44673));
    defparam i29161_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i29163_4_lut (.I0(n44673), .I1(n44654), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44675));
    defparam i29163_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29162_3_lut (.I0(n49369), .I1(n49339), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44674));
    defparam i29162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3265));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29138_4_lut (.I0(n19_adj_3265), .I1(\data_out_frame[22]_c [4]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n44650));
    defparam i29138_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29139_3_lut (.I0(n49345), .I1(n44650), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44651));
    defparam i29139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32748_4_lut (.I0(n49375), .I1(n44651), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(tx_data[4]));   // verilog/coms.v(103[34:55])
    defparam i32748_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31468_2_lut (.I0(\data_out_frame[0][3] ), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n46586));   // verilog/coms.v(103[34:55])
    defparam i31468_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(n46586), .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3266));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf0c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3267));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29158_3_lut (.I0(n5_adj_3267), .I1(n6_adj_3266), .I2(n46420), 
            .I3(GND_net), .O(n44670));
    defparam i29158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29160_4_lut (.I0(n44670), .I1(n49483), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44672));
    defparam i29160_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29159_3_lut (.I0(n49441), .I1(n49381), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44671));
    defparam i29159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31785_2_lut (.I0(\data_out_frame[0][2] ), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n46583));   // verilog/coms.v(103[34:55])
    defparam i31785_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3268));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5][2] ), 
            .I1(n46583), .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3269));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha00c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3270));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29183_4_lut (.I0(n19_adj_3268), .I1(\data_out_frame[22]_c [2]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n44695));
    defparam i29183_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29184_3_lut (.I0(n49405), .I1(n44695), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44696));
    defparam i29184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29155_3_lut (.I0(n5_adj_3270), .I1(n6_adj_3269), .I2(n46420), 
            .I3(GND_net), .O(n44667));
    defparam i29155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29157_4_lut (.I0(n44667), .I1(n44696), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44669));
    defparam i29157_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29156_3_lut (.I0(n49453), .I1(n49447), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44668));
    defparam i29156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3271));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31461_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n46974));   // verilog/coms.v(103[34:55])
    defparam i31461_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3272));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29180_4_lut (.I0(n19_adj_3271), .I1(\data_out_frame[22] [1]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n44692));
    defparam i29180_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29181_3_lut (.I0(n49399), .I1(n44692), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44693));
    defparam i29181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29130_4_lut (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[0] [2]), .O(n44642));
    defparam i29130_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29152_4_lut (.I0(n5_adj_3272), .I1(n46974), .I2(n46420), 
            .I3(byte_transmit_counter[0]), .O(n44664));
    defparam i29152_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i29154_4_lut (.I0(n44664), .I1(n44693), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n44666));
    defparam i29154_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29153_3_lut (.I0(n49465), .I1(n49459), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n44665));
    defparam i29153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [4]), .O(n38));
    defparam i14_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15_4_lut_adj_1016 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[2] [6]), .O(n39));
    defparam i15_4_lut_adj_1016.LUT_INIT = 16'h0002;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[1] [3]), .O(n37));
    defparam i13_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i29126_4_lut (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [1]), .O(n44638));
    defparam i29126_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1017 (.I0(n37), .I1(n39), .I2(n38), .I3(n44642), 
            .O(n46));
    defparam i22_4_lut_adj_1017.LUT_INIT = 16'h0080;
    SB_LUT4 i29128_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[2] [5]), .O(n44640));
    defparam i29128_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_3_lut (.I0(n44640), .I1(n46), .I2(n44638), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_1924 [3]));
    defparam i23_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2056_3_lut (.I0(n3362), .I1(\FRAME_MATCHER.state[2] ), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n5025));
    defparam i2056_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(n5025), .I1(\FRAME_MATCHER.state_31__N_1924 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n22498));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h8888;
    SB_LUT4 i15231_3_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n63_adj_3273), 
            .I2(n63_adj_3274), .I3(GND_net), .O(n122));   // verilog/coms.v(137[4] 139[7])
    defparam i15231_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_313_Select_2_i5_4_lut (.I0(n122), .I1(n22525), .I2(n2854), 
            .I3(n63), .O(n5));
    defparam select_313_Select_2_i5_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i15227_rep_520_2_lut (.I0(n122), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n50013));   // verilog/coms.v(140[4] 142[7])
    defparam i15227_rep_520_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n49360_bdd_4_lut (.I0(n49360), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n49363));
    defparam n49360_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15189_1_lut (.I0(n28588), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1508));
    defparam i15189_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_4_lut_adj_1019 (.I0(n42916), .I1(\data_out_frame[18] [4]), 
            .I2(\data_out_frame[18] [6]), .I3(n43175), .O(n10_adj_3277));
    defparam i4_4_lut_adj_1019.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1020 (.I0(\data_out_frame[16] [2]), .I1(n10_adj_3277), 
            .I2(n38965), .I3(GND_net), .O(n44444));
    defparam i5_3_lut_adj_1020.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_adj_1021 (.I0(n42813), .I1(n42863), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3278));
    defparam i2_2_lut_adj_1021.LUT_INIT = 16'h9999;
    SB_LUT4 i6_4_lut_adj_1022 (.I0(n43114), .I1(\data_out_frame[20] [7]), 
            .I2(n23356), .I3(n39622), .O(n14_adj_3279));
    defparam i6_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1023 (.I0(n44450), .I1(n14_adj_3279), .I2(n10_adj_3278), 
            .I3(n38900), .O(n44218));
    defparam i7_4_lut_adj_1023.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1024 (.I0(n38998), .I1(n39622), .I2(n43036), 
            .I3(n6_adj_3280), .O(n43632));
    defparam i4_4_lut_adj_1024.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(\data_out_frame[16] [6]), .I1(n39315), 
            .I2(GND_net), .I3(GND_net), .O(n39622));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1026 (.I0(\data_out_frame[19] [2]), .I1(n42863), 
            .I2(n43152), .I3(\data_out_frame[17] [1]), .O(n42936));
    defparam i1_4_lut_adj_1026.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1027 (.I0(n43304), .I1(n1692), .I2(\data_out_frame[16] [7]), 
            .I3(n43307), .O(n10_adj_3281));
    defparam i4_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1028 (.I0(n42883), .I1(n10_adj_3281), .I2(n23431), 
            .I3(n4_adj_3282), .O(n44450));
    defparam i5_4_lut_adj_1028.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1029 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[14] [7]), 
            .I2(n8_adj_3283), .I3(n1506), .O(n42813));   // verilog/coms.v(69[16:41])
    defparam i1_4_lut_adj_1029.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1030 (.I0(\data_out_frame[19] [4]), .I1(n43152), 
            .I2(n42813), .I3(\data_out_frame[17] [2]), .O(n43111));   // verilog/coms.v(69[16:41])
    defparam i3_4_lut_adj_1030.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1031 (.I0(n43111), .I1(n43127), .I2(\data_out_frame[19] [5]), 
            .I3(GND_net), .O(n44248));   // verilog/coms.v(69[16:41])
    defparam i2_3_lut_adj_1031.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1032 (.I0(n23371), .I1(n23546), .I2(n43205), 
            .I3(n42955), .O(n16_adj_3284));
    defparam i6_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1033 (.I0(\data_out_frame[8] [5]), .I1(n43187), 
            .I2(n43289), .I3(n42868), .O(n17_adj_3285));
    defparam i7_4_lut_adj_1033.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(\data_out_frame[17] [3]), .I1(n17_adj_3285), 
            .I2(n15_adj_3286), .I3(n16_adj_3284), .O(n38926));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1035 (.I0(n42791), .I1(n43096), .I2(n43062), 
            .I3(n38926), .O(n12_adj_3287));
    defparam i5_4_lut_adj_1035.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1036 (.I0(n22703), .I1(n12_adj_3287), .I2(n43268), 
            .I3(n39004), .O(n43849));
    defparam i6_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1037 (.I0(n39599), .I1(n43062), .I2(GND_net), 
            .I3(GND_net), .O(n23311));
    defparam i1_2_lut_adj_1037.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1038 (.I0(n23071), .I1(n23546), .I2(n23368), 
            .I3(n23522), .O(n44332));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33845 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n49354));
    defparam byte_transmit_counter_0__bdd_4_lut_33845.LUT_INIT = 16'he4aa;
    SB_LUT4 n49354_bdd_4_lut (.I0(n49354), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n49357));
    defparam n49354_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1039 (.I0(n43334), .I1(n42836), .I2(n44332), 
            .I3(GND_net), .O(n43127));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1039.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1040 (.I0(n43127), .I1(\data_out_frame[20] [0]), 
            .I2(n42791), .I3(GND_net), .O(n43062));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1040.LUT_INIT = 16'h9696;
    SB_LUT4 i10385_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[10] [0]), 
            .I3(IntegralLimit[0]), .O(n23803));
    defparam i10385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10386_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[0] ), .O(n23804));
    defparam i10386_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10387_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[3] [0]), 
            .I3(\Ki[0] ), .O(n23805));
    defparam i10387_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10388_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[4] [0]), 
            .I3(\Kd[0] ), .O(n23806));
    defparam i10388_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10389_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[19] [0]), 
            .I3(gearBoxRatio[0]), .O(n23807));
    defparam i10389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1041 (.I0(\FRAME_MATCHER.state_31__N_1860[1] ), .I1(\FRAME_MATCHER.state_31__N_1892 [1]), 
            .I2(n43447), .I3(n22512), .O(n6_adj_3289));
    defparam i2_4_lut_adj_1041.LUT_INIT = 16'h0ace;
    SB_LUT4 i3_4_lut_adj_1042 (.I0(n43773), .I1(n6_adj_3289), .I2(\FRAME_MATCHER.state_31__N_1988 [1]), 
            .I3(n22525), .O(n49489));
    defparam i3_4_lut_adj_1042.LUT_INIT = 16'hddfd;
    SB_LUT4 i10392_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[1] [0]), 
            .I3(control_mode[0]), .O(n23810));
    defparam i10392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1043 (.I0(\FRAME_MATCHER.state[3] ), .I1(n113), 
            .I2(n11_adj_3290), .I3(GND_net), .O(n13_adj_3291));
    defparam i1_3_lut_adj_1043.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut_adj_1044 (.I0(n22520), .I1(n13_adj_3291), .I2(n22492), 
            .I3(\FRAME_MATCHER.state_31__N_1924 [3]), .O(n42198));
    defparam i1_4_lut_adj_1044.LUT_INIT = 16'hdccc;
    SB_LUT4 i15514_2_lut (.I0(\FRAME_MATCHER.state [5]), .I1(n34109), .I2(GND_net), 
            .I3(GND_net), .O(n28918));
    defparam i15514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15515_2_lut (.I0(\FRAME_MATCHER.state [6]), .I1(n34109), .I2(GND_net), 
            .I3(GND_net), .O(n28920));
    defparam i15515_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10393_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[7] [0]), 
            .I3(\PWMLimit[0] ), .O(n23811));
    defparam i10393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(n34109), .I1(\FRAME_MATCHER.state [16]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3178));
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h8888;
    SB_LUT4 i33129_2_lut_3_lut (.I0(n5025), .I1(n3362), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(GND_net), .O(n23610));
    defparam i33129_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1046 (.I0(n34109), .I1(\FRAME_MATCHER.state [18]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3176));
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_1047 (.I0(\data_out_frame[18] [4]), .I1(n10_adj_3292), 
            .I2(\data_out_frame[16] [3]), .I3(\data_out_frame[16] [1]), 
            .O(n44037));
    defparam i5_3_lut_4_lut_adj_1047.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1048 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[9] [2]), .I3(GND_net), .O(n42865));
    defparam i1_2_lut_3_lut_adj_1048.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1049 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[11] [4]), .I3(GND_net), .O(n23485));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1049.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(n34109), .I1(\FRAME_MATCHER.state [20]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3175));
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1051 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[6] [2]), .O(n42752));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1052 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[13] [3]), .I3(GND_net), .O(n22664));   // verilog/coms.v(82[17:63])
    defparam i1_2_lut_3_lut_adj_1052.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1053 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[16] [0]), .I3(\data_out_frame[17] [7]), 
            .O(n42974));
    defparam i2_3_lut_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1054 (.I0(\data_out_frame[8] [6]), .I1(n42948), 
            .I2(n43156), .I3(\data_out_frame[5] [0]), .O(n22187));
    defparam i2_3_lut_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1055 (.I0(\data_out_frame[6] [5]), .I1(n43292), 
            .I2(n43199), .I3(\data_out_frame[9] [1]), .O(n1512));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1056 (.I0(\FRAME_MATCHER.state [23]), .I1(n34109), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3173));
    defparam i1_2_lut_adj_1056.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1057 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n43199));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1057.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(n34109), .I1(\FRAME_MATCHER.state [24]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3171));
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1059 (.I0(n22700), .I1(\data_out_frame[11] [5]), 
            .I2(n43280), .I3(GND_net), .O(n42789));   // verilog/coms.v(82[17:70])
    defparam i1_2_lut_3_lut_adj_1059.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(n34109), .I1(\FRAME_MATCHER.state [25]), 
            .I2(GND_net), .I3(GND_net), .O(n28932));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'h8888;
    SB_LUT4 i3_3_lut_4_lut_adj_1061 (.I0(\data_out_frame[12] [5]), .I1(n22292), 
            .I2(n1608), .I3(\data_out_frame[13] [0]), .O(n42871));
    defparam i3_3_lut_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(n34109), .I1(\FRAME_MATCHER.state [26]), 
            .I2(GND_net), .I3(GND_net), .O(n28539));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h8888;
    SB_LUT4 i15229_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n63_adj_3274), 
            .I2(n63_adj_3273), .I3(n63), .O(\FRAME_MATCHER.state_31__N_1860[1] ));
    defparam i15229_2_lut_3_lut_4_lut.LUT_INIT = 16'h80ff;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(\FRAME_MATCHER.state [27]), .I1(n34109), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3168));
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_1064 (.I0(\data_out_frame[8] [0]), .I1(n10_adj_3293), 
            .I2(\data_out_frame[7] [7]), .I3(\data_out_frame[5] [5]), .O(n23335));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[5][2] ), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[7] [3]), .O(n43280));   // verilog/coms.v(82[17:70])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10962_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[9] [0]), 
            .I3(IntegralLimit[8]), .O(n24380));
    defparam i10962_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1065 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n22712));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1065.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1066 (.I0(\data_out_frame[5][2] ), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n23128));
    defparam i1_2_lut_3_lut_adj_1066.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1067 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[10] [7]), .I3(GND_net), .O(n43159));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1067.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1068 (.I0(\FRAME_MATCHER.state [1]), .I1(n42694), 
            .I2(n20285), .I3(n22510), .O(n11_adj_3290));
    defparam i1_4_lut_adj_1068.LUT_INIT = 16'h4454;
    SB_LUT4 i1_2_lut_4_lut_adj_1069 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[13] [2]), .I3(n22664), .O(n43187));   // verilog/coms.v(82[17:63])
    defparam i1_2_lut_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1070 (.I0(\data_out_frame[6] [2]), .I1(n42836), 
            .I2(\data_out_frame[10] [4]), .I3(n43165), .O(n22292));
    defparam i1_2_lut_4_lut_adj_1070.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1071 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n22520), .I3(GND_net), .O(n44266));   // verilog/coms.v(156[5:29])
    defparam i2_3_lut_adj_1071.LUT_INIT = 16'hfbfb;
    SB_LUT4 i4_4_lut_adj_1072 (.I0(n22518), .I1(n28588), .I2(n43773), 
            .I3(n44266), .O(n10_adj_3294));
    defparam i4_4_lut_adj_1072.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_1073 (.I0(\FRAME_MATCHER.state[0] ), .I1(n10_adj_3294), 
            .I2(n63_adj_3288), .I3(n22517), .O(n2119));
    defparam i5_4_lut_adj_1073.LUT_INIT = 16'hc080;
    SB_LUT4 i10963_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[10] [7]), 
            .I3(IntegralLimit[7]), .O(n24381));
    defparam i10963_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_2_lut_3_lut (.I0(\data_out_frame[18] [5]), .I1(n22967), .I2(n43152), 
            .I3(GND_net), .O(n16_adj_3295));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1074 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[8] [4]), 
            .I2(n42786), .I3(\data_out_frame[10] [5]), .O(n43020));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i29662_2_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n46420));
    defparam i29662_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(\FRAME_MATCHER.state [1]), .I1(n22524), 
            .I2(GND_net), .I3(GND_net), .O(n22517));   // verilog/coms.v(201[5:16])
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_3_lut_adj_1076 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[14] [7]), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n6_adj_3296));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1076.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1077 (.I0(byte_transmit_counter_c[7]), .I1(byte_transmit_counter_c[6]), 
            .I2(byte_transmit_counter_c[5]), .I3(GND_net), .O(n4_adj_3297));   // verilog/coms.v(202[6] 209[9])
    defparam i2_3_lut_adj_1077.LUT_INIT = 16'hfefe;
    SB_LUT4 i15619_4_lut (.I0(n46420), .I1(n4_adj_3297), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n29027));
    defparam i15619_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_3_lut_adj_1078 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [3]), 
            .I2(n39653), .I3(GND_net), .O(n43175));
    defparam i1_2_lut_3_lut_adj_1078.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1079 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[14] [4]), 
            .I2(n43325), .I3(GND_net), .O(n39653));
    defparam i1_2_lut_3_lut_adj_1079.LUT_INIT = 16'h9696;
    SB_LUT4 i15214_4_lut (.I0(n10_adj_3298), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n22570), .O(n3758));   // verilog/coms.v(244[9:58])
    defparam i15214_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i12_3_lut_4_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[18] [7]), .I3(n42746), .O(n35));
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [28]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3299));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1080 (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i [22]), 
            .I2(\FRAME_MATCHER.i [27]), .I3(\FRAME_MATCHER.i [15]), .O(n36));
    defparam i14_4_lut_adj_1080.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1081 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [19]), 
            .I2(\FRAME_MATCHER.i [16]), .I3(\FRAME_MATCHER.i [9]), .O(n44306));
    defparam i3_4_lut_adj_1081.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1082 (.I0(\FRAME_MATCHER.i [18]), .I1(n44306), 
            .I2(\FRAME_MATCHER.i [8]), .I3(\FRAME_MATCHER.i [25]), .O(n34));
    defparam i12_4_lut_adj_1082.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n36), .I2(n26_adj_3299), 
            .I3(\FRAME_MATCHER.i [10]), .O(n40));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [29]), .I3(\FRAME_MATCHER.i [24]), .O(n38_adj_3300));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n34), .I2(\FRAME_MATCHER.i [23]), 
            .I3(GND_net), .O(n39_adj_3301));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1083 (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [13]), 
            .I2(\FRAME_MATCHER.i [14]), .I3(\FRAME_MATCHER.i [30]), .O(n37_adj_3302));
    defparam i15_4_lut_adj_1083.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1084 (.I0(n37_adj_3302), .I1(n39_adj_3301), .I2(n38_adj_3300), 
            .I3(n40), .O(n22570));
    defparam i21_4_lut_adj_1084.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1085 (.I0(n22636), .I1(\data_in[1] [4]), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [6]), .O(n10_adj_3303));
    defparam i3_4_lut_adj_1085.LUT_INIT = 16'hffef;
    SB_LUT4 i29122_3_lut (.I0(\data_in[3] [0]), .I1(\data_in[2] [2]), .I2(\data_in[1] [5]), 
            .I3(GND_net), .O(n44634));
    defparam i29122_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6_4_lut_adj_1086 (.I0(n44634), .I1(\data_in[2] [4]), .I2(n10_adj_3303), 
            .I3(\data_in[0] [3]), .O(n22422));
    defparam i6_4_lut_adj_1086.LUT_INIT = 16'hfdff;
    SB_LUT4 i6_4_lut_adj_1087 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_3304));
    defparam i6_4_lut_adj_1087.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1088 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_3305));
    defparam i7_4_lut_adj_1088.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1089 (.I0(n17_adj_3305), .I1(\data_in[1] [6]), 
            .I2(n16_adj_3304), .I3(\data_in[3] [7]), .O(n22501));
    defparam i9_4_lut_adj_1089.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1090 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_3306));
    defparam i4_4_lut_adj_1090.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1091 (.I0(\data_in[3] [4]), .I1(n10_adj_3306), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n22636));
    defparam i5_3_lut_adj_1091.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_2_lut_adj_1092 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3307));
    defparam i2_2_lut_adj_1092.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1093 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_3308));
    defparam i6_4_lut_adj_1093.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1094 (.I0(\data_in[3] [6]), .I1(n14_adj_3308), 
            .I2(n10_adj_3307), .I3(\data_in[2] [1]), .O(n22544));
    defparam i7_4_lut_adj_1094.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_1095 (.I0(\data_in[2] [4]), .I1(n22544), .I2(\data_in[1] [5]), 
            .I3(n22636), .O(n18_adj_3309));
    defparam i7_4_lut_adj_1095.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1096 (.I0(\data_in[0] [6]), .I1(n18_adj_3309), 
            .I2(\data_in[3] [0]), .I3(n22501), .O(n20_adj_3310));
    defparam i9_4_lut_adj_1096.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut_adj_1097 (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3311));
    defparam i4_2_lut_adj_1097.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1098 (.I0(n15_adj_3311), .I1(n20_adj_3310), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_adj_3273));
    defparam i10_4_lut_adj_1098.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1099 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n22422), .O(n16_adj_3312));
    defparam i6_4_lut_adj_1099.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1100 (.I0(n22501), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_3313));
    defparam i7_4_lut_adj_1100.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1101 (.I0(n17_adj_3313), .I1(\data_in[3] [5]), 
            .I2(n16_adj_3312), .I3(\data_in[3] [3]), .O(n63_adj_3274));
    defparam i9_4_lut_adj_1101.LUT_INIT = 16'hfbff;
    SB_LUT4 i5883_2_lut (.I0(n63_adj_3274), .I1(n63_adj_3273), .I2(GND_net), 
            .I3(GND_net), .O(n19202));   // verilog/coms.v(137[4] 139[7])
    defparam i5883_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8_4_lut_adj_1102 (.I0(n22544), .I1(\data_in[1] [3]), .I2(n22422), 
            .I3(\data_in[2] [0]), .O(n20_adj_3314));
    defparam i8_4_lut_adj_1102.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1103 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19_adj_3315));
    defparam i7_4_lut_adj_1103.LUT_INIT = 16'hfeff;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33840 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n49348));
    defparam byte_transmit_counter_0__bdd_4_lut_33840.LUT_INIT = 16'he4aa;
    SB_LUT4 i29124_4_lut (.I0(\data_in[1] [2]), .I1(\data_in[3] [2]), .I2(\data_in[2] [5]), 
            .I3(\data_in[0] [5]), .O(n44636));
    defparam i29124_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n44636), .I1(n19_adj_3315), .I2(n20_adj_3314), 
            .I3(GND_net), .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1104 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n43124));
    defparam i1_2_lut_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1105 (.I0(n22416), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3316));
    defparam i1_2_lut_adj_1105.LUT_INIT = 16'heeee;
    SB_LUT4 i15209_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_3316), .I3(\FRAME_MATCHER.i [1]), .O(n737));   // verilog/coms.v(152[9:60])
    defparam i15209_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\FRAME_MATCHER.state[0] ), .I1(n22520), 
            .I2(GND_net), .I3(GND_net), .O(n22510));   // verilog/coms.v(239[5:25])
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(n20156), .I1(n737), .I2(GND_net), .I3(GND_net), 
            .O(n20285));
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h2222;
    SB_LUT4 i10411_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[13] [0]), 
            .I3(\deadband[0] ), .O(n23829));
    defparam i10411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1108 (.I0(n22525), .I1(n44), .I2(n20211), .I3(n40_adj_3317), 
            .O(n34109));
    defparam i2_4_lut_adj_1108.LUT_INIT = 16'hffdc;
    SB_LUT4 i1_2_lut_adj_1109 (.I0(\FRAME_MATCHER.state [31]), .I1(n34109), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3164));
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1110 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[13] [1]), .I3(GND_net), .O(n23194));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_3_lut_adj_1110.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1111 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[7] [0]), .I3(n43265), .O(n6_adj_3318));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1112 (.I0(\data_out_frame[6] [1]), .I1(n10_adj_3319), 
            .I2(\data_out_frame[12] [7]), .I3(n1506), .O(n23431));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i10927_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[4] [6]), 
            .I3(\Kd[6] ), .O(n24345));
    defparam i10927_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1113 (.I0(n43165), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[12] [3]), .I3(n23335), .O(n38682));
    defparam i1_2_lut_3_lut_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i10928_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[4] [5]), 
            .I3(\Kd[5] ), .O(n24346));
    defparam i10928_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10929_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[4] [4]), 
            .I3(\Kd[4] ), .O(n24347));
    defparam i10929_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_2_lut_3_lut_4_lut (.I0(\data_out_frame[14] [7]), .I1(n22700), 
            .I2(\data_out_frame[11] [5]), .I3(n43280), .O(n15_adj_3286));
    defparam i5_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1114 (.I0(\FRAME_MATCHER.state[0] ), 
            .I1(\FRAME_MATCHER.state [1]), .I2(n22524), .I3(n745), .O(n3));
    defparam i1_2_lut_3_lut_4_lut_adj_1114.LUT_INIT = 16'h0800;
    SB_LUT4 i27940_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n22520), .I3(n3758), .O(n43447));
    defparam i27940_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1115 (.I0(n2854), .I1(n63), .I2(n63_adj_3274), 
            .I3(n63_adj_3273), .O(n20211));   // verilog/coms.v(216[6] 218[9])
    defparam i1_2_lut_3_lut_4_lut_adj_1115.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1116 (.I0(n63), .I1(n63_adj_3274), 
            .I2(n63_adj_3273), .I3(n2119), .O(n44));   // verilog/coms.v(152[6] 154[9])
    defparam i1_2_lut_3_lut_4_lut_adj_1116.LUT_INIT = 16'h8000;
    SB_LUT4 i10930_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[4] [3]), 
            .I3(\Kd[3] ), .O(n24348));
    defparam i10930_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1117 (.I0(n20156), .I1(n737), .I2(n22512), 
            .I3(GND_net), .O(n40_adj_3317));   // verilog/coms.v(147[5:27])
    defparam i1_2_lut_3_lut_adj_1117.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_adj_1118 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n22520), .I3(GND_net), .O(n22512));   // verilog/coms.v(147[5:27])
    defparam i1_2_lut_3_lut_adj_1118.LUT_INIT = 16'hfbfb;
    SB_LUT4 i2_2_lut_3_lut_adj_1119 (.I0(n63), .I1(n63_adj_3274), .I2(n63_adj_3273), 
            .I3(GND_net), .O(n20156));   // verilog/coms.v(152[6] 154[9])
    defparam i2_2_lut_3_lut_adj_1119.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut (.I0(n22518), .I1(n63), .I2(n19202), .I3(n745), 
            .O(n113));   // verilog/coms.v(201[5:16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i171_3_lut_4_lut (.I0(n22511), .I1(n63), .I2(n19202), .I3(n3758), 
            .O(n48));   // verilog/coms.v(112[11:12])
    defparam i171_3_lut_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_3_lut_adj_1120 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n22520), .I3(GND_net), .O(n22511));   // verilog/coms.v(239[5:25])
    defparam i1_2_lut_3_lut_adj_1120.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1121 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n22524), .I3(GND_net), .O(n22518));   // verilog/coms.v(201[5:16])
    defparam i1_2_lut_3_lut_adj_1121.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_3_lut_4_lut_adj_1122 (.I0(\FRAME_MATCHER.state[0] ), .I1(n2854), 
            .I2(n20156), .I3(n22524), .O(n42694));
    defparam i1_3_lut_4_lut_adj_1122.LUT_INIT = 16'h0020;
    SB_LUT4 i10964_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[10] [6]), 
            .I3(IntegralLimit[6]), .O(n24382));
    defparam i10964_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1123 (.I0(\FRAME_MATCHER.state[3] ), .I1(n20156), 
            .I2(n2119), .I3(n48), .O(n41956));
    defparam i1_3_lut_4_lut_adj_1123.LUT_INIT = 16'haa80;
    SB_LUT4 i10931_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[4] [2]), 
            .I3(\Kd[2] ), .O(n24349));
    defparam i10931_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10932_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[4] [1]), 
            .I3(\Kd[1] ), .O(n24350));
    defparam i10932_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10933_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[3] [7]), 
            .I3(\Ki[7] ), .O(n24351));
    defparam i10933_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10934_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[3] [6]), 
            .I3(\Ki[6] ), .O(n24352));
    defparam i10934_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10935_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[3] [5]), 
            .I3(\Ki[5] ), .O(n24353));
    defparam i10935_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10936_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[3] [4]), 
            .I3(\Ki[4] ), .O(n24354));
    defparam i10936_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10937_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[3] [3]), 
            .I3(\Ki[3] ), .O(n24355));
    defparam i10937_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1124 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(n42874), .I3(GND_net), .O(n42791));
    defparam i1_2_lut_3_lut_adj_1124.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1125 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[12] [7]), .I3(GND_net), .O(n23546));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1125.LUT_INIT = 16'h9696;
    SB_LUT4 i10938_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[3] [2]), 
            .I3(\Ki[2] ), .O(n24356));
    defparam i10938_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1126 (.I0(\data_out_frame[19] [1]), .I1(n42936), 
            .I2(\data_out_frame[16] [6]), .I3(n39315), .O(n43950));
    defparam i2_3_lut_4_lut_adj_1126.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31802_2_lut (.I0(\data_out_frame[22]_c [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46624));
    defparam i31802_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3149));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10939_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[3] [1]), 
            .I3(\Ki[1] ), .O(n24357));
    defparam i10939_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1127 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[19] [1]), .I3(GND_net), .O(n6_adj_3280));
    defparam i1_2_lut_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_LUT4 i10940_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[7] ), .O(n24358));
    defparam i10940_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10549_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[6] [1]), 
            .I3(\PWMLimit[9] ), .O(n23967));
    defparam i10549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10550_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[6] [0]), 
            .I3(\PWMLimit[8] ), .O(n23968));
    defparam i10550_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14911_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[7] [7]), 
            .I3(\PWMLimit[7] ), .O(n28310));
    defparam i14911_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10552_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[7] [6]), 
            .I3(\PWMLimit[6] ), .O(n23970));
    defparam i10552_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14829_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[7] [5]), 
            .I3(\PWMLimit[5] ), .O(n23971));
    defparam i14829_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14778_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[7] [4]), 
            .I3(\PWMLimit[4] ), .O(n23972));
    defparam i14778_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10555_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[7] [3]), 
            .I3(\PWMLimit[3] ), .O(n23973));
    defparam i10555_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10556_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[7] [2]), 
            .I3(\PWMLimit[2] ), .O(n23974));
    defparam i10556_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10557_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[7] [1]), 
            .I3(\PWMLimit[1] ), .O(n23975));
    defparam i10557_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10558_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[1] [7]), 
            .I3(control_mode[7]), .O(n23976));
    defparam i10558_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10559_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[1] [6]), 
            .I3(control_mode[6]), .O(n23977));
    defparam i10559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n49348_bdd_4_lut (.I0(n49348), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n49351));
    defparam n49348_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33835 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n49342));
    defparam byte_transmit_counter_0__bdd_4_lut_33835.LUT_INIT = 16'he4aa;
    SB_LUT4 n49342_bdd_4_lut (.I0(n49342), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n49345));
    defparam n49342_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33830 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n49336));
    defparam byte_transmit_counter_0__bdd_4_lut_33830.LUT_INIT = 16'he4aa;
    SB_LUT4 n49336_bdd_4_lut (.I0(n49336), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n49339));
    defparam n49336_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10560_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[1] [5]), 
            .I3(control_mode[5]), .O(n23978));
    defparam i10560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10561_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[1] [4]), 
            .I3(control_mode[4]), .O(n23979));
    defparam i10561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10562_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[1] [3]), 
            .I3(control_mode[3]), .O(n23980));
    defparam i10562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10563_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[1] [2]), 
            .I3(control_mode[2]), .O(n23981));
    defparam i10563_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10564_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[1] [1]), 
            .I3(control_mode[1]), .O(n23982));
    defparam i10564_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10965_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[10] [5]), 
            .I3(IntegralLimit[5]), .O(n24383));
    defparam i10965_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10941_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[6] ), .O(n24359));
    defparam i10941_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10966_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[10] [4]), 
            .I3(IntegralLimit[4]), .O(n24384));
    defparam i10966_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10967_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[10] [3]), 
            .I3(IntegralLimit[3]), .O(n24385));
    defparam i10967_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1128 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n29039), .I3(GND_net), .O(n4_adj_3258));
    defparam i1_2_lut_3_lut_adj_1128.LUT_INIT = 16'hfefe;
    SB_LUT4 i10968_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[10] [2]), 
            .I3(IntegralLimit[2]), .O(n24386));
    defparam i10968_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_567_i1_3_lut_4_lut (.I0(n31_adj_3255), .I1(n28473), .I2(tx_transmit_N_2639), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n29029));   // verilog/coms.v(143[4] 283[11])
    defparam mux_567_i1_3_lut_4_lut.LUT_INIT = 16'h0fee;
    SB_LUT4 i27839_4_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n29039), .I3(n2_adj_3321), .O(n43341));
    defparam i27839_4_lut_4_lut.LUT_INIT = 16'hfbf8;
    SB_LUT4 i1_2_lut_3_lut_adj_1129 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n2_adj_3321));
    defparam i1_2_lut_3_lut_adj_1129.LUT_INIT = 16'ha8a8;
    SB_LUT4 i10969_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[10] [1]), 
            .I3(IntegralLimit[1]), .O(n24387));
    defparam i10969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n20014));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h4046;
    SB_LUT4 i10942_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[5] ), .O(n24360));
    defparam i10942_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_1045_i15_2_lut_3_lut (.I0(n5_adj_3190), .I1(n23446), .I2(\data_in_frame[4] [6]), 
            .I3(GND_net), .O(n15_adj_3256));   // verilog/coms.v(225[9:81])
    defparam equal_1045_i15_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i10943_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[4] ), .O(n24361));
    defparam i10943_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10954_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[8] [0]), 
            .I3(IntegralLimit[16]), .O(n24372));
    defparam i10954_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10953_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[8] [1]), 
            .I3(IntegralLimit[17]), .O(n24371));
    defparam i10953_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10952_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[8] [2]), 
            .I3(IntegralLimit[18]), .O(n24370));
    defparam i10952_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10951_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[8] [3]), 
            .I3(IntegralLimit[19]), .O(n24369));
    defparam i10951_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10950_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[8] [4]), 
            .I3(IntegralLimit[20]), .O(n24368));
    defparam i10950_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10961_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[9] [1]), 
            .I3(IntegralLimit[9]), .O(n24379));
    defparam i10961_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33825 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n49330));
    defparam byte_transmit_counter_0__bdd_4_lut_33825.LUT_INIT = 16'he4aa;
    SB_LUT4 n49330_bdd_4_lut (.I0(n49330), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n49333));
    defparam n49330_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10926_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[4] [7]), 
            .I3(\Kd[7] ), .O(n24344));
    defparam i10926_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10925_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[19] [1]), 
            .I3(gearBoxRatio[1]), .O(n24343));
    defparam i10925_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10924_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[19] [2]), 
            .I3(gearBoxRatio[2]), .O(n24342));
    defparam i10924_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10923_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[19] [3]), 
            .I3(gearBoxRatio[3]), .O(n24341));
    defparam i10923_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10912_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[18] [6]), 
            .I3(gearBoxRatio[14]), .O(n24330));
    defparam i10912_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10913_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[18] [5]), 
            .I3(gearBoxRatio[13]), .O(n24331));
    defparam i10913_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10914_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[18] [4]), 
            .I3(gearBoxRatio[12]), .O(n24332));
    defparam i10914_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10915_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[18] [3]), 
            .I3(gearBoxRatio[11]), .O(n24333));
    defparam i10915_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10916_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[18] [2]), 
            .I3(gearBoxRatio[10]), .O(n24334));
    defparam i10916_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10959_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[9] [3]), 
            .I3(IntegralLimit[11]), .O(n24377));
    defparam i10959_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10917_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[18] [1]), 
            .I3(gearBoxRatio[9]), .O(n24335));
    defparam i10917_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10918_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[18] [0]), 
            .I3(gearBoxRatio[8]), .O(n24336));
    defparam i10918_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10919_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[19] [7]), 
            .I3(gearBoxRatio[7]), .O(n24337));
    defparam i10919_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10920_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[19] [6]), 
            .I3(gearBoxRatio[6]), .O(n24338));
    defparam i10920_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10921_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[19] [5]), 
            .I3(gearBoxRatio[5]), .O(n24339));
    defparam i10921_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut_adj_1130 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(\FRAME_MATCHER.state [1]), 
            .O(n4_adj_3252));
    defparam i1_4_lut_4_lut_adj_1130.LUT_INIT = 16'h0504;
    SB_LUT4 i6617_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n19960));
    defparam i6617_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i10922_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[19] [4]), 
            .I3(gearBoxRatio[4]), .O(n24340));
    defparam i10922_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11071_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[12] [0]), 
            .I3(\deadband[8] ), .O(n24489));
    defparam i11071_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11072_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[12] [1]), 
            .I3(\deadband[9] ), .O(n24490));
    defparam i11072_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10903_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[17] [7]), 
            .I3(gearBoxRatio[23]), .O(n24321));
    defparam i10903_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10904_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[17] [6]), 
            .I3(gearBoxRatio[22]), .O(n24322));
    defparam i10904_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10905_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[17] [5]), 
            .I3(gearBoxRatio[21]), .O(n24323));
    defparam i10905_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1131 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n22524), .I3(GND_net), .O(n63_adj_3288));   // verilog/coms.v(248[5:27])
    defparam i1_2_lut_3_lut_adj_1131.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1132 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[9] [4]), .I3(\data_out_frame[7] [1]), .O(n22700));   // verilog/coms.v(82[17:70])
    defparam i2_3_lut_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[17] [6]), .I3(GND_net), .O(n16_adj_3322));   // verilog/coms.v(82[17:70])
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1133 (.I0(\data_in_frame[21] [7]), .I1(n42904), 
            .I2(n43172), .I3(n23467), .O(n42902));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1134 (.I0(\data_out_frame[13] [1]), .I1(n43187), 
            .I2(n42871), .I3(n42789), .O(n38984));   // verilog/coms.v(82[17:63])
    defparam i2_3_lut_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1135 (.I0(n39672), .I1(\data_in_frame[17] [6]), 
            .I2(n42782), .I3(n39055), .O(n6_adj_3240));
    defparam i1_2_lut_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1136 (.I0(\data_out_frame[13] [1]), .I1(n43187), 
            .I2(n43211), .I3(n42987), .O(n43307));   // verilog/coms.v(82[17:63])
    defparam i2_3_lut_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1137 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(n42999), .I3(GND_net), .O(n6_adj_3194));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1137.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1138 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[6] [3]), .I3(\data_out_frame[6] [1]), .O(n42786));   // verilog/coms.v(70[16:34])
    defparam i3_3_lut_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1139 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[11] [0]), .O(n42868));   // verilog/coms.v(70[16:34])
    defparam i2_3_lut_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i10906_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[17] [4]), 
            .I3(gearBoxRatio[20]), .O(n24324));
    defparam i10906_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10907_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[17] [3]), 
            .I3(gearBoxRatio[19]), .O(n24325));
    defparam i10907_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut_adj_1140 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[8] [2]), .I3(n5_adj_3323), .O(n42836));   // verilog/coms.v(70[16:34])
    defparam i3_3_lut_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1141 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[9] [2]), .I3(GND_net), .O(n42826));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1141.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1142 (.I0(n43050), .I1(n43256), .I2(n23032), 
            .I3(n43077), .O(n23113));
    defparam i1_2_lut_4_lut_adj_1142.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1143 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n43169));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1143.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1144 (.I0(n5_adj_3190), .I1(n23446), .I2(\data_in_frame[7] [0]), 
            .I3(GND_net), .O(n23164));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_3_lut_adj_1144.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1145 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[1] [1]), .O(n43117));   // verilog/coms.v(70[16:34])
    defparam i2_3_lut_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1146 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n42762));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1146.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1147 (.I0(n5_adj_3190), .I1(n23446), .I2(\data_in_frame[7] [2]), 
            .I3(GND_net), .O(n43053));
    defparam i1_2_lut_3_lut_adj_1147.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1148 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[1] [0]), .O(n23528));   // verilog/coms.v(68[16:69])
    defparam i2_3_lut_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1149 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[9] [0]), .I3(\data_out_frame[11] [1]), .O(n23368));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i10908_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[17] [2]), 
            .I3(gearBoxRatio[18]), .O(n24326));
    defparam i10908_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1150 (.I0(n43165), .I1(\data_out_frame[12] [4]), 
            .I2(n42883), .I3(GND_net), .O(n23000));
    defparam i2_2_lut_3_lut_adj_1150.LUT_INIT = 16'h9696;
    SB_LUT4 i10909_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[17] [1]), 
            .I3(gearBoxRatio[17]), .O(n24327));
    defparam i10909_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1151 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[7] [4]), 
            .I2(\data_in_frame[7] [5]), .I3(GND_net), .O(n43081));
    defparam i1_2_lut_3_lut_adj_1151.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1152 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(\data_in_frame[9] [4]), .I3(n43259), .O(n8_adj_3184));
    defparam i3_3_lut_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i10910_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[17] [0]), 
            .I3(gearBoxRatio[16]), .O(n24328));
    defparam i10910_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1153 (.I0(n38682), .I1(n42929), .I2(\data_out_frame[14] [5]), 
            .I3(\data_out_frame[17] [0]), .O(n42863));
    defparam i1_2_lut_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1154 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[7] [3]), 
            .I2(\data_in_frame[9] [5]), .I3(GND_net), .O(n43050));
    defparam i1_2_lut_3_lut_adj_1154.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1155 (.I0(n38682), .I1(n42929), .I2(\data_out_frame[14] [5]), 
            .I3(n1713), .O(n38998));
    defparam i1_2_lut_4_lut_adj_1155.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_4_lut_adj_1156 (.I0(n38984), .I1(n1608), .I2(n43307), 
            .I3(n1592), .O(n8_adj_3283));
    defparam i3_3_lut_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1157 (.I0(n38984), .I1(n1608), .I2(\data_out_frame[15] [1]), 
            .I3(GND_net), .O(n43205));
    defparam i1_2_lut_3_lut_adj_1157.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1158 (.I0(\data_in_frame[4] [7]), .I1(n39661), 
            .I2(n43053), .I3(GND_net), .O(n43074));
    defparam i1_2_lut_3_lut_adj_1158.LUT_INIT = 16'h6969;
    SB_LUT4 i10911_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[18] [7]), 
            .I3(gearBoxRatio[15]), .O(n24329));
    defparam i10911_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10391_3_lut_4_lut (.I0(n8), .I1(n42714), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n23809));
    defparam i10391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10733_3_lut_4_lut (.I0(n8), .I1(n42714), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n24151));
    defparam i10733_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1159 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[9] [1]), 
            .I2(Kp_23__N_325), .I3(\data_in_frame[7] [0]), .O(n23519));   // verilog/coms.v(71[16:43])
    defparam i2_3_lut_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i10734_3_lut_4_lut (.I0(n8), .I1(n42714), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n24152));
    defparam i10734_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1160 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[15] [7]), 
            .I2(\data_in_frame[14] [0]), .I3(n43310), .O(n6_adj_3182));
    defparam i1_2_lut_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i10735_3_lut_4_lut (.I0(n8), .I1(n42714), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n24153));
    defparam i10735_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10736_3_lut_4_lut (.I0(n8), .I1(n42714), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n24154));
    defparam i10736_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10737_3_lut_4_lut (.I0(n8), .I1(n42714), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n24155));
    defparam i10737_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14777_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[13] [4]), 
            .I3(\deadband[4] ), .O(n24485));
    defparam i14777_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1161 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[14] [0]), 
            .I2(n43310), .I3(GND_net), .O(n42907));
    defparam i1_2_lut_3_lut_adj_1161.LUT_INIT = 16'h9696;
    SB_LUT4 i10738_3_lut_4_lut (.I0(n8), .I1(n42714), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n24156));
    defparam i10738_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10739_3_lut_4_lut (.I0(n8), .I1(n42714), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n24157));
    defparam i10739_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1162 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[16] [2]), 
            .I2(n39257), .I3(GND_net), .O(n43064));
    defparam i1_2_lut_3_lut_adj_1162.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1163 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n28467), .O(n42723));   // verilog/coms.v(149[7:23])
    defparam i2_3_lut_4_lut_adj_1163.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_4_lut_adj_1164 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n28467), .O(n42714));   // verilog/coms.v(149[7:23])
    defparam i2_3_lut_4_lut_adj_1164.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_2_lut_3_lut_adj_1165 (.I0(\data_in_frame[8] [0]), .I1(Kp_23__N_458), 
            .I2(\data_in_frame[5] [6]), .I3(GND_net), .O(n22826));   // verilog/coms.v(82[17:28])
    defparam i2_2_lut_3_lut_adj_1165.LUT_INIT = 16'h9696;
    SB_LUT4 equal_61_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(149[7:23])
    defparam equal_61_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_60_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3126));   // verilog/coms.v(149[7:23])
    defparam equal_60_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i10725_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42714), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n24143));
    defparam i10725_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11068_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[13] [5]), 
            .I3(\deadband[5] ), .O(n24486));
    defparam i11068_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1166 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[12] [2]), 
            .I2(n22977), .I3(\data_in_frame[10] [0]), .O(n43262));
    defparam i2_3_lut_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i10726_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42714), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n24144));
    defparam i10726_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10727_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42714), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n24145));
    defparam i10727_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1167 (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[3] [4]), 
            .I2(n42821), .I3(\data_in_frame[1] [1]), .O(n43274));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1168 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(\data_in_frame[6] [0]), .I3(\data_in_frame[10] [2]), .O(n42925));
    defparam i1_2_lut_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i10728_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42714), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n24146));
    defparam i10728_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10729_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42714), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n24147));
    defparam i10729_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10730_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42714), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n24148));
    defparam i10730_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11069_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[13] [6]), 
            .I3(\deadband[6] ), .O(n24487));
    defparam i11069_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1169 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(n42840), .I3(\data_in_frame[14] [7]), .O(n43228));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i10731_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42714), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n24149));
    defparam i10731_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1170 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [7]), .I3(GND_net), .O(n43253));   // verilog/coms.v(225[9:81])
    defparam i1_2_lut_3_lut_adj_1170.LUT_INIT = 16'h9696;
    SB_LUT4 i10732_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42714), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n24150));
    defparam i10732_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10717_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42714), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n24135));
    defparam i10717_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10718_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42714), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n24136));
    defparam i10718_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1171 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[1] [5]), .O(n43008));   // verilog/coms.v(225[9:81])
    defparam i2_3_lut_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i10719_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42714), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n24137));
    defparam i10719_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10720_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42714), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n24138));
    defparam i10720_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10721_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42714), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n24139));
    defparam i10721_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10722_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42714), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n24140));
    defparam i10722_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10723_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42714), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n24141));
    defparam i10723_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14912_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[13] [7]), 
            .I3(\deadband[7] ), .O(n24488));
    defparam i14912_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1172 (.I0(Kp_23__N_515), .I1(n43059), .I2(n10_adj_3155), 
            .I3(n5_adj_3186), .O(n23018));
    defparam i5_3_lut_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i10724_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42714), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n24142));
    defparam i10724_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1173 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [1]), 
            .I2(\data_in_frame[16] [4]), .I3(\data_in_frame[16] [2]), .O(n43105));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(148[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1174 (.I0(n23519), .I1(\data_in_frame[8] [7]), 
            .I2(n22858), .I3(GND_net), .O(n42913));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_3_lut_adj_1174.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1175 (.I0(n23519), .I1(n43283), .I2(n10_adj_3151), 
            .I3(\data_in_frame[10] [7]), .O(n23266));   // verilog/coms.v(71[16:43])
    defparam i5_3_lut_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 equal_66_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3132));   // verilog/coms.v(149[7:23])
    defparam equal_66_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_3_lut_adj_1176 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[8] [3]), 
            .I2(\data_in_frame[10] [4]), .I3(GND_net), .O(n43322));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1176.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1177 (.I0(n44318), .I1(n44327), .I2(\data_in_frame[18] [7]), 
            .I3(\data_in_frame[16] [6]), .O(n42919));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1178 (.I0(\data_in_frame[8] [0]), .I1(n7), 
            .I2(\data_in_frame[14] [4]), .I3(\data_in_frame[12] [3]), .O(n14_adj_3148));
    defparam i5_3_lut_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 equal_67_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3131));   // verilog/coms.v(149[7:23])
    defparam equal_67_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i10709_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42714), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n24127));
    defparam i10709_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10710_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42714), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n24128));
    defparam i10710_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10711_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42714), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n24129));
    defparam i10711_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1179 (.I0(n42969), .I1(\data_in_frame[14] [5]), 
            .I2(n23018), .I3(n44327), .O(Kp_23__N_945));
    defparam i1_2_lut_4_lut_adj_1179.LUT_INIT = 16'h9669;
    SB_LUT4 i10712_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42714), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n24130));
    defparam i10712_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10713_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42714), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n24131));
    defparam i10713_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10714_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42714), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n24132));
    defparam i10714_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10715_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42714), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n24133));
    defparam i10715_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10716_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42714), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n24134));
    defparam i10716_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10701_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42714), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n24119));
    defparam i10701_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10702_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42714), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n24120));
    defparam i10702_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10703_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42714), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n24121));
    defparam i10703_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10704_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42714), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n24122));
    defparam i10704_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10705_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42714), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n24123));
    defparam i10705_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10706_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42714), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n24124));
    defparam i10706_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10707_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42714), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n24125));
    defparam i10707_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10708_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42714), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n24126));
    defparam i10708_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_64_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3135));   // verilog/coms.v(149[7:23])
    defparam equal_64_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_65_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3133));   // verilog/coms.v(149[7:23])
    defparam equal_65_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i10693_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42714), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n24111));
    defparam i10693_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10694_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42714), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n24112));
    defparam i10694_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10949_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[8] [5]), 
            .I3(IntegralLimit[21]), .O(n24367));
    defparam i10949_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10695_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42714), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n24113));
    defparam i10695_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10696_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42714), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n24114));
    defparam i10696_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10697_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42714), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n24115));
    defparam i10697_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10698_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42714), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n24116));
    defparam i10698_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10699_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42714), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n24117));
    defparam i10699_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1180 (.I0(n42868), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[6] [5]), .I3(n43159), .O(n10_adj_3319));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1181 (.I0(\data_out_frame[6] [1]), .I1(n10_adj_3319), 
            .I2(\data_out_frame[12] [7]), .I3(GND_net), .O(n1592));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1182 (.I0(n42746), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[15] [5]), .I3(GND_net), .O(n42874));
    defparam i2_3_lut_adj_1182.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1183 (.I0(n22967), .I1(n38965), .I2(GND_net), 
            .I3(GND_net), .O(n38679));
    defparam i1_2_lut_adj_1183.LUT_INIT = 16'h6666;
    SB_LUT4 i10700_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42714), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n24118));
    defparam i10700_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10685_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42714), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n24103));
    defparam i10685_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1184 (.I0(n22766), .I1(n42886), .I2(n1713), .I3(n38679), 
            .O(n38980));   // verilog/coms.v(71[16:43])
    defparam i3_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i10686_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42714), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n24104));
    defparam i10686_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1185 (.I0(\data_out_frame[15] [3]), .I1(n23194), 
            .I2(\data_out_frame[19] [7]), .I3(n23326), .O(n12_adj_3325));   // verilog/coms.v(71[16:43])
    defparam i5_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1186 (.I0(\data_out_frame[17] [5]), .I1(n12_adj_3325), 
            .I2(n42874), .I3(n23431), .O(n39334));   // verilog/coms.v(71[16:43])
    defparam i6_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i10687_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42714), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n24105));
    defparam i10687_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1187 (.I0(\data_out_frame[16] [2]), .I1(n42749), 
            .I2(n38679), .I3(n44449), .O(n39432));
    defparam i3_4_lut_adj_1187.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1188 (.I0(n38994), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[13] [2]), .I3(n1661), .O(n44381));
    defparam i3_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i10688_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42714), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n24106));
    defparam i10688_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1189 (.I0(n43169), .I1(n43156), .I2(n44381), 
            .I3(GND_net), .O(n14_adj_3326));
    defparam i5_3_lut_adj_1189.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1190 (.I0(n43292), .I1(\data_out_frame[15] [6]), 
            .I2(n43331), .I3(n42857), .O(n15_adj_3327));
    defparam i6_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i10689_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42714), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n24107));
    defparam i10689_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10690_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42714), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n24108));
    defparam i10690_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1191 (.I0(n15_adj_3327), .I1(\data_out_frame[8] [6]), 
            .I2(n14_adj_3326), .I3(n42871), .O(n44449));
    defparam i8_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i10691_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42714), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n24109));
    defparam i10691_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10948_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[8] [6]), 
            .I3(IntegralLimit[22]), .O(n24366));
    defparam i10948_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42916));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1193 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(n39342), .I3(GND_net), .O(n39601));
    defparam i2_3_lut_adj_1193.LUT_INIT = 16'h9696;
    SB_LUT4 i10692_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42714), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n24110));
    defparam i10692_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1194 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n23356));
    defparam i1_2_lut_adj_1194.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42776));
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_LUT4 i15212_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n22416), .I3(\FRAME_MATCHER.i [31]), .O(n2854));
    defparam i15212_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 i1842_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [4]), .O(n10_adj_3298));
    defparam i1842_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i15140_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n28540));
    defparam i15140_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 equal_63_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3324));
    defparam equal_63_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i10677_3_lut_4_lut (.I0(n28540), .I1(n42714), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n24095));
    defparam i10677_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n22675));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1197 (.I0(n23488), .I1(n42863), .I2(GND_net), 
            .I3(GND_net), .O(n42889));
    defparam i1_2_lut_adj_1197.LUT_INIT = 16'h9999;
    SB_LUT4 i10678_3_lut_4_lut (.I0(n28540), .I1(n42714), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n24096));
    defparam i10678_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10679_3_lut_4_lut (.I0(n28540), .I1(n42714), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n24097));
    defparam i10679_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1198 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42749));
    defparam i1_2_lut_adj_1198.LUT_INIT = 16'h6666;
    SB_LUT4 i14786_3_lut_4_lut (.I0(n28540), .I1(n42714), .I2(\data_in_frame[7] [4]), 
            .I3(rx_data[4]), .O(n24098));
    defparam i14786_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n23243));
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i10947_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[8] [7]), 
            .I3(IntegralLimit[23]), .O(n24365));
    defparam i10947_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10681_3_lut_4_lut (.I0(n28540), .I1(n42714), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n24099));
    defparam i10681_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1200 (.I0(n22187), .I1(n23368), .I2(n42752), 
            .I3(n22639), .O(n43211));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i10684_3_lut_4_lut (.I0(n28540), .I1(n42714), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n24102));
    defparam i10684_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1201 (.I0(\data_out_frame[13] [2]), .I1(n43211), 
            .I2(\data_out_frame[13] [4]), .I3(\data_out_frame[15] [4]), 
            .O(n42746));
    defparam i3_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n22766));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43250));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h6666;
    SB_LUT4 i10683_3_lut_4_lut (.I0(n28540), .I1(n42714), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n24101));
    defparam i10683_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10682_3_lut_4_lut (.I0(n28540), .I1(n42714), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n24100));
    defparam i10682_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1204 (.I0(\data_out_frame[6] [7]), .I1(n23371), 
            .I2(n43087), .I3(n6_adj_3318), .O(n1506));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i10669_3_lut_4_lut (.I0(n8), .I1(n42723), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n24087));
    defparam i10669_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42886));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i10670_3_lut_4_lut (.I0(n8), .I1(n42723), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n24088));
    defparam i10670_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10671_3_lut_4_lut (.I0(n8), .I1(n42723), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n24089));
    defparam i10671_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10672_3_lut_4_lut (.I0(n8), .I1(n42723), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n24090));
    defparam i10672_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10946_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[1] ), .O(n24364));
    defparam i10946_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10673_3_lut_4_lut (.I0(n8), .I1(n42723), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n24091));
    defparam i10673_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10674_3_lut_4_lut (.I0(n8), .I1(n42723), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n24092));
    defparam i10674_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10945_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[2] ), .O(n24363));
    defparam i10945_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10675_3_lut_4_lut (.I0(n8), .I1(n42723), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n24093));
    defparam i10675_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10676_3_lut_4_lut (.I0(n8), .I1(n42723), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n24094));
    defparam i10676_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1206 (.I0(n1506), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43215));
    defparam i1_2_lut_adj_1206.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_out_frame[19] [5]), .I1(n23488), 
            .I2(GND_net), .I3(GND_net), .O(n43096));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i10661_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42723), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n24079));
    defparam i10661_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10662_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42723), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n24080));
    defparam i10662_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10663_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42723), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n24081));
    defparam i10663_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10960_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[9] [2]), 
            .I3(IntegralLimit[10]), .O(n24378));
    defparam i10960_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10664_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42723), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n24082));
    defparam i10664_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(n38984), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n38994));
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_LUT4 i10665_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42723), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n24083));
    defparam i10665_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10666_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42723), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n24084));
    defparam i10666_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42857));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43023));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1211 (.I0(n23485), .I1(n43124), .I2(n23128), 
            .I3(n22720), .O(n12_adj_3328));
    defparam i5_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i10667_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42723), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n24085));
    defparam i10667_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10668_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42723), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n24086));
    defparam i10668_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1212 (.I0(\data_out_frame[11] [6]), .I1(n12_adj_3328), 
            .I2(\data_out_frame[14] [0]), .I3(n42826), .O(n38965));
    defparam i6_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1213 (.I0(\data_out_frame[14] [3]), .I1(n42880), 
            .I2(n22720), .I3(\data_out_frame[12] [2]), .O(n23488));   // verilog/coms.v(82[17:70])
    defparam i3_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1214 (.I0(n43190), .I1(n43193), .I2(\data_out_frame[14] [2]), 
            .I3(n42945), .O(n12_adj_3329));
    defparam i5_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1215 (.I0(\data_out_frame[10] [0]), .I1(n12_adj_3329), 
            .I2(n43301), .I3(\data_out_frame[12] [1]), .O(n23317));
    defparam i6_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(n23317), .I1(n23488), .I2(GND_net), 
            .I3(GND_net), .O(n1713));
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1217 (.I0(\data_out_frame[13] [5]), .I1(n42987), 
            .I2(n38965), .I3(GND_net), .O(n39342));
    defparam i2_3_lut_adj_1217.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42955));
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1219 (.I0(n23356), .I1(n42977), .I2(n43205), 
            .I3(\data_out_frame[14] [5]), .O(n43304));
    defparam i1_4_lut_adj_1219.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1220 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(n42955), .I3(\data_out_frame[13] [2]), .O(n43334));
    defparam i3_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i10653_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42723), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n24071));
    defparam i10653_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1221 (.I0(n39342), .I1(n22967), .I2(n38998), 
            .I3(n1692), .O(n12_adj_3330));
    defparam i5_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1222 (.I0(n42977), .I1(n12_adj_3330), .I2(n23000), 
            .I3(n38994), .O(n44360));
    defparam i6_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i6_2_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3331));
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1223 (.I0(n43334), .I1(n43304), .I2(n38986), 
            .I3(\data_out_frame[11] [5]), .O(n23));
    defparam i9_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1224 (.I0(\data_out_frame[9] [1]), .I1(n42974), 
            .I2(n43023), .I3(n43124), .O(n44199));
    defparam i3_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1225 (.I0(n23194), .I1(n23096), .I2(n44199), 
            .I3(n43277), .O(n22));
    defparam i8_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1226 (.I0(n23), .I1(\data_out_frame[15] [6]), 
            .I2(n20_adj_3331), .I3(n44360), .O(n26_adj_3332));
    defparam i12_4_lut_adj_1226.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1227 (.I0(\data_out_frame[17] [3]), .I1(n26_adj_3332), 
            .I2(n22), .I3(\data_out_frame[13] [4]), .O(n44382));
    defparam i13_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1228 (.I0(n42939), .I1(n23243), .I2(n42749), 
            .I3(n1512), .O(n38_adj_3333));
    defparam i15_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1229 (.I0(n43096), .I1(n43215), .I2(\data_out_frame[19] [2]), 
            .I3(n42886), .O(n36_adj_3334));
    defparam i13_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1230 (.I0(n39653), .I1(n43250), .I2(\data_out_frame[19] [4]), 
            .I3(n43202), .O(n37_adj_3335));
    defparam i14_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i10944_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[3] ), .O(n24362));
    defparam i10944_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17_4_lut (.I0(n44382), .I1(n42889), .I2(\data_out_frame[16] [7]), 
            .I3(n22675), .O(n40_adj_3336));
    defparam i17_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i10654_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42723), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n24072));
    defparam i10654_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21_4_lut_adj_1231 (.I0(n35), .I1(n37_adj_3335), .I2(n36_adj_3334), 
            .I3(n38_adj_3333), .O(n44_adj_3337));
    defparam i21_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i10655_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42723), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n24073));
    defparam i10655_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10656_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42723), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n24074));
    defparam i10656_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10657_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42723), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n24075));
    defparam i10657_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10658_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42723), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n24076));
    defparam i10658_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10659_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42723), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n24077));
    defparam i10659_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10660_3_lut_4_lut (.I0(n8_adj_3131), .I1(n42723), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n24078));
    defparam i10660_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10645_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42723), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n24063));
    defparam i10645_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10646_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42723), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n24064));
    defparam i10646_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10647_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42723), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n24065));
    defparam i10647_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10648_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42723), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n24066));
    defparam i10648_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10649_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42723), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n24067));
    defparam i10649_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10650_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42723), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n24068));
    defparam i10650_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10651_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42723), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n24069));
    defparam i10651_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10652_3_lut_4_lut (.I0(n8_adj_3132), .I1(n42723), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n24070));
    defparam i10652_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10637_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42723), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n24055));
    defparam i10637_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10638_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42723), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n24056));
    defparam i10638_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10639_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42723), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n24057));
    defparam i10639_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10640_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42723), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n24058));
    defparam i10640_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut_adj_1232 (.I0(n43023), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[19] [3]), .I3(n23326), .O(n39_adj_3338));
    defparam i16_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1233 (.I0(\data_out_frame[17] [5]), .I1(n39_adj_3338), 
            .I2(n44_adj_3337), .I3(n40_adj_3336), .O(n43114));
    defparam i1_4_lut_adj_1233.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1234 (.I0(n23000), .I1(n42776), .I2(\data_out_frame[18] [7]), 
            .I3(\data_out_frame[16] [5]), .O(n12_adj_3339));
    defparam i5_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1235 (.I0(\data_out_frame[14] [6]), .I1(n12_adj_3339), 
            .I2(n42889), .I3(n22292), .O(n39315));
    defparam i6_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_out_frame[14] [4]), .I1(n43325), 
            .I2(GND_net), .I3(GND_net), .O(n42929));
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i10641_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42723), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n24059));
    defparam i10641_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1237 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n22703));
    defparam i1_2_lut_adj_1237.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1238 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n42945));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1238.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1239 (.I0(\data_out_frame[7] [4]), .I1(n42945), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n22720));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1239.LUT_INIT = 16'h9696;
    SB_LUT4 i10642_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42723), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n24060));
    defparam i10642_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1240 (.I0(n42789), .I1(\data_out_frame[12] [0]), 
            .I2(\data_out_frame[14] [1]), .I3(n43093), .O(n10_adj_3340));   // verilog/coms.v(82[17:70])
    defparam i4_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1241 (.I0(n22720), .I1(n10_adj_3340), .I2(\data_out_frame[13] [7]), 
            .I3(GND_net), .O(n22967));   // verilog/coms.v(82[17:70])
    defparam i5_3_lut_adj_1241.LUT_INIT = 16'h9696;
    SB_LUT4 i10643_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42723), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n24061));
    defparam i10643_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10958_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[9] [4]), 
            .I3(IntegralLimit[12]), .O(n24376));
    defparam i10958_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1242 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3341));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1243 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[5] [5]), 
            .I2(n43108), .I3(n6_adj_3341), .O(n42883));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i10644_3_lut_4_lut (.I0(n8_adj_3133), .I1(n42723), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n24062));
    defparam i10644_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10629_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42723), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n24047));
    defparam i10629_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10630_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42723), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n24048));
    defparam i10630_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10631_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42723), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n24049));
    defparam i10631_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14790_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42723), .I2(\data_in_frame[13] [4]), 
            .I3(rx_data[4]), .O(n24050));
    defparam i14790_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i10633_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42723), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n24051));
    defparam i10633_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i936_2_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1692));   // verilog/coms.v(68[16:27])
    defparam i936_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10636_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42723), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n24054));
    defparam i10636_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1244 (.I0(n23000), .I1(n23329), .I2(n43020), 
            .I3(n6_adj_3296), .O(n43152));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_out_frame[18] [5]), .I1(n22967), 
            .I2(GND_net), .I3(GND_net), .O(n43268));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\data_out_frame[12] [3]), .I1(n23335), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3282));
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 i10635_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42723), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n24053));
    defparam i10635_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\data_out_frame[15] [0]), .I1(n38682), 
            .I2(GND_net), .I3(GND_net), .O(n38986));
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43036));
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 i10634_3_lut_4_lut (.I0(n8_adj_3135), .I1(n42723), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n24052));
    defparam i10634_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1249 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n28467), .O(n42698));   // verilog/coms.v(149[7:23])
    defparam i2_3_lut_4_lut_adj_1249.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_4_lut_adj_1250 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n22570), .I3(\FRAME_MATCHER.i [4]), .O(n22416));   // verilog/coms.v(149[7:23])
    defparam i2_3_lut_4_lut_adj_1250.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1251 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n42098));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1251.LUT_INIT = 16'he0e0;
    SB_LUT4 i15095_2_lut_3_lut (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n28493));   // verilog/coms.v(112[11:12])
    defparam i15095_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i9_4_lut_adj_1252 (.I0(n43036), .I1(n38986), .I2(n43020), 
            .I3(\data_out_frame[14] [5]), .O(n22_adj_3342));
    defparam i9_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(\data_out_frame[14] [7]), .I1(n39315), .I2(n43114), 
            .I3(GND_net), .O(n20_adj_3343));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1253 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n42044));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1253.LUT_INIT = 16'he0e0;
    SB_LUT4 i11_4_lut_adj_1254 (.I0(n43175), .I1(n22_adj_3342), .I2(n16_adj_3295), 
            .I3(\data_out_frame[17] [0]), .O(n24));
    defparam i11_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1255 (.I0(n43165), .I1(n24), .I2(n20_adj_3343), 
            .I3(n42776), .O(n38900));
    defparam i12_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43331));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1257 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n42100));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1257.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3344));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1259 (.I0(n23151), .I1(\data_out_frame[8] [2]), 
            .I2(n42809), .I3(n6_adj_3344), .O(n43165));   // verilog/coms.v(70[16:34])
    defparam i4_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1260 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n42102));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1260.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1261 (.I0(\data_out_frame[6] [2]), .I1(n42836), 
            .I2(\data_out_frame[10] [4]), .I3(GND_net), .O(n23329));   // verilog/coms.v(70[16:34])
    defparam i2_3_lut_adj_1261.LUT_INIT = 16'h9696;
    SB_LUT4 i11061_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[13] [1]), 
            .I3(\deadband[1] ), .O(n24479));
    defparam i11061_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1262 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n42104));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1262.LUT_INIT = 16'he0e0;
    SB_LUT4 i11065_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[13] [2]), 
            .I3(\deadband[2] ), .O(n24483));
    defparam i11065_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1263 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n42106));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1263.LUT_INIT = 16'he0e0;
    SB_LUT4 i905_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1661));   // verilog/coms.v(82[17:28])
    defparam i905_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1264 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n42108));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1264.LUT_INIT = 16'he0e0;
    SB_LUT4 i11066_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[13] [3]), 
            .I3(\deadband[3] ), .O(n24484));
    defparam i11066_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n23071));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42779));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43265));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1268 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n42110));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1268.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1269 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n42112));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1269.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1270 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n22639));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1270.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42898));
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1272 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n42809));
    defparam i2_3_lut_adj_1272.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1273 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n42114));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1273.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1274 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n42116));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1274.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1275 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n7_adj_3177));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1275.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1276 (.I0(\data_out_frame[6] [0]), .I1(n42809), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n43108));
    defparam i2_3_lut_adj_1276.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1277 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n42118));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1277.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_adj_1278 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3345));
    defparam i2_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1279 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n28495));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1279.LUT_INIT = 16'he0e0;
    SB_LUT4 i6_4_lut_adj_1280 (.I0(n22712), .I1(\data_out_frame[5][2] ), 
            .I2(n43108), .I3(\data_out_frame[10] [2]), .O(n14_adj_3346));
    defparam i6_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1281 (.I0(\data_out_frame[7] [4]), .I1(n14_adj_3346), 
            .I2(n10_adj_3345), .I3(\data_out_frame[12] [3]), .O(n43325));
    defparam i7_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1282 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n42120));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1282.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1283 (.I0(\data_out_frame[8] [4]), .I1(n42786), 
            .I2(\data_out_frame[10] [5]), .I3(GND_net), .O(n22738));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1283.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1284 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n7_adj_3174));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1284.LUT_INIT = 16'he0e0;
    SB_LUT4 i10957_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[9] [5]), 
            .I3(IntegralLimit[13]), .O(n24375));
    defparam i10957_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1285 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n42122));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1285.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1286 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n42124));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1286.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1287 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n7_adj_3172));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1287.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1288 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n7_adj_3170));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1288.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1289 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n42136));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1289.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1290 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n7_adj_3169));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1290.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1291 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n7_adj_3167));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1291.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1292 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n42200));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1292.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1293 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n42084));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1293.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1294 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n42088));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1294.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1295 (.I0(n113), .I1(n48), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n7_adj_3163));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_3_lut_adj_1295.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1296 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n41958));
    defparam i1_2_lut_3_lut_adj_1296.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1297 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n42030));
    defparam i1_2_lut_3_lut_adj_1297.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1298 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n42028));
    defparam i1_2_lut_3_lut_adj_1298.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1299 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n42026));
    defparam i1_2_lut_3_lut_adj_1299.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1300 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n42024));
    defparam i1_2_lut_3_lut_adj_1300.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1301 (.I0(n42799), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[5] [4]), .O(n43301));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i15070_2_lut_2_lut_3_lut (.I0(n28588), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n28467));
    defparam i15070_2_lut_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i10955_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[9] [7]), 
            .I3(IntegralLimit[15]), .O(n24373));
    defparam i10955_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1302 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n42022));
    defparam i1_2_lut_3_lut_adj_1302.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1303 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n42020));
    defparam i1_2_lut_3_lut_adj_1303.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1304 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3323));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1305 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n42018));
    defparam i1_2_lut_3_lut_adj_1305.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1306 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n42016));
    defparam i1_2_lut_3_lut_adj_1306.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1307 (.I0(n5_adj_3323), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[8] [2]), .I3(\data_out_frame[6] [2]), .O(n43289));   // verilog/coms.v(70[16:34])
    defparam i4_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1308 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n42014));
    defparam i1_2_lut_3_lut_adj_1308.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1309 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43218));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1309.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43002));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n23151));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1312 (.I0(\data_out_frame[5][2] ), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n42860));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1312.LUT_INIT = 16'h9696;
    SB_LUT4 i10956_3_lut_4_lut (.I0(n28496), .I1(n63_adj_3288), .I2(\data_in_frame[9] [6]), 
            .I3(IntegralLimit[14]), .O(n24374));
    defparam i10956_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1313 (.I0(\data_in_frame[2] [3]), .I1(n42772), 
            .I2(n5_adj_3190), .I3(\data_in_frame[4] [5]), .O(n22858));   // verilog/coms.v(161[9:87])
    defparam i2_3_lut_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1314 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[9] [6]), 
            .I2(n42860), .I3(\data_out_frame[7] [5]), .O(n43093));   // verilog/coms.v(82[17:70])
    defparam i3_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1315 (.I0(n43002), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[10] [1]), .I3(n43218), .O(n10_adj_3293));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1316 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n42012));
    defparam i1_2_lut_3_lut_adj_1316.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1317 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n42010));
    defparam i1_2_lut_3_lut_adj_1317.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43087));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1319 (.I0(n23335), .I1(n43093), .I2(\data_out_frame[12] [1]), 
            .I3(GND_net), .O(n42880));   // verilog/coms.v(82[17:70])
    defparam i2_3_lut_adj_1319.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1320 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n42008));
    defparam i1_2_lut_3_lut_adj_1320.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1321 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43190));
    defparam i1_2_lut_adj_1321.LUT_INIT = 16'h6666;
    SB_LUT4 i18_4_lut_adj_1322 (.I0(\data_out_frame[11] [0]), .I1(n43190), 
            .I2(n42880), .I3(n43087), .O(n52));   // verilog/coms.v(70[16:27])
    defparam i18_4_lut_adj_1322.LUT_INIT = 16'h6996;
    SB_LUT4 i26_3_lut (.I0(\data_out_frame[7] [7]), .I1(n52), .I2(\data_out_frame[8] [0]), 
            .I3(GND_net), .O(n60_adj_3347));   // verilog/coms.v(70[16:27])
    defparam i26_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i24_4_lut_adj_1323 (.I0(\data_out_frame[7] [1]), .I1(n42786), 
            .I2(n43289), .I3(\data_out_frame[8] [1]), .O(n58_adj_3348));   // verilog/coms.v(70[16:27])
    defparam i24_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1324 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n41966));
    defparam i1_2_lut_3_lut_adj_1324.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1325 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n41892));
    defparam i1_2_lut_3_lut_adj_1325.LUT_INIT = 16'he0e0;
    SB_LUT4 i25_4_lut_adj_1326 (.I0(n43301), .I1(n42860), .I2(n43169), 
            .I3(n42762), .O(n59_adj_3349));   // verilog/coms.v(70[16:27])
    defparam i25_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1327 (.I0(n42948), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[9] [0]), .I3(n22639), .O(n57_adj_3350));   // verilog/coms.v(70[16:27])
    defparam i23_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1328 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n41998));
    defparam i1_2_lut_3_lut_adj_1328.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1329 (.I0(\data_in_frame[2] [3]), .I1(n42772), 
            .I2(\data_in_frame[0] [0]), .I3(n42769), .O(Kp_23__N_319));   // verilog/coms.v(161[9:87])
    defparam i2_3_lut_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1330 (.I0(n22738), .I1(n43280), .I2(n43325), 
            .I3(\data_out_frame[12] [4]), .O(n38_adj_3351));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(n44), .I1(n11_adj_3290), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n42004));
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'he0e0;
    SB_LUT4 i20_4_lut_adj_1332 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[11] [3]), .I3(n22700), .O(n54));   // verilog/coms.v(70[16:27])
    defparam i20_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1333 (.I0(n43265), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[6] [3]), .I3(n43218), .O(n56_adj_3352));   // verilog/coms.v(70[16:27])
    defparam i22_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1334 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [2]), .I3(GND_net), .O(n6_adj_3185));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1334.LUT_INIT = 16'h9696;
    SB_LUT4 i21_4_lut_adj_1335 (.I0(n42779), .I1(n42898), .I2(n23071), 
            .I3(n43193), .O(n55_adj_3353));   // verilog/coms.v(70[16:27])
    defparam i21_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i32_4_lut (.I0(n57_adj_3350), .I1(n59_adj_3349), .I2(n58_adj_3348), 
            .I3(n60_adj_3347), .O(n66));   // verilog/coms.v(70[16:27])
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut_adj_1336 (.I0(n43159), .I1(n54), .I2(n38_adj_3351), 
            .I3(n42977), .O(n61_adj_3354));   // verilog/coms.v(70[16:27])
    defparam i27_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut_adj_1337 (.I0(n61_adj_3354), .I1(n66), .I2(n55_adj_3353), 
            .I3(n56_adj_3352), .O(n1608));   // verilog/coms.v(70[16:27])
    defparam i33_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1338 (.I0(\FRAME_MATCHER.state [1]), .I1(n19202), 
            .I2(n2854), .I3(n63), .O(\FRAME_MATCHER.state_31__N_1988 [1]));
    defparam i2_3_lut_4_lut_adj_1338.LUT_INIT = 16'hf8ff;
    SB_LUT4 i1_2_lut_adj_1339 (.I0(\data_out_frame[12] [5]), .I1(n22292), 
            .I2(GND_net), .I3(GND_net), .O(n42977));
    defparam i1_2_lut_adj_1339.LUT_INIT = 16'h6666;
    SB_LUT4 i15151_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n19202), 
            .I2(n737), .I3(n63), .O(\FRAME_MATCHER.state_31__N_1892 [1]));
    defparam i15151_2_lut_3_lut_4_lut.LUT_INIT = 16'hf8ff;
    SB_LUT4 i1_4_lut_4_lut_adj_1340 (.I0(n63), .I1(n737), .I2(n3), .I3(n22512), 
            .O(n5_adj_3));   // verilog/coms.v(152[6] 154[9])
    defparam i1_4_lut_4_lut_adj_1340.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_2_lut_adj_1341 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42799));
    defparam i1_2_lut_adj_1341.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1342 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23096));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1342.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(n22700), .I1(\data_out_frame[11] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43121));
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h6666;
    SB_LUT4 i10621_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42723), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n24039));
    defparam i10621_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10622_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42723), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n24040));
    defparam i10622_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10623_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42723), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n24041));
    defparam i10623_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10624_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42723), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n24042));
    defparam i10624_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10625_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42723), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n24043));
    defparam i10625_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10626_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42723), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n24044));
    defparam i10626_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1344 (.I0(n23313), .I1(\data_out_frame[5][2] ), 
            .I2(n42799), .I3(\data_out_frame[7] [3]), .O(n43277));
    defparam i3_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i10627_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42723), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n24045));
    defparam i10627_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10628_3_lut_4_lut (.I0(n8_adj_3324), .I1(n42723), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n24046));
    defparam i10628_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10613_3_lut_4_lut (.I0(n28540), .I1(n42723), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n24031));
    defparam i10613_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10614_3_lut_4_lut (.I0(n28540), .I1(n42723), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n24032));
    defparam i10614_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10615_3_lut_4_lut (.I0(n28540), .I1(n42723), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n24033));
    defparam i10615_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10616_3_lut_4_lut (.I0(n28540), .I1(n42723), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n24034));
    defparam i10616_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10617_3_lut_4_lut (.I0(n28540), .I1(n42723), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n24035));
    defparam i10617_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10618_3_lut_4_lut (.I0(n28540), .I1(n42723), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n24036));
    defparam i10618_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10619_3_lut_4_lut (.I0(n28540), .I1(n42723), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n24037));
    defparam i10619_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1345 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[11] [2]), .I3(n43199), .O(n43156));
    defparam i3_4_lut_adj_1345.LUT_INIT = 16'h6996;
    SB_LUT4 i10620_3_lut_4_lut (.I0(n28540), .I1(n42723), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n24038));
    defparam i10620_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1346 (.I0(\data_out_frame[20] [5]), .I1(n44037), 
            .I2(n39432), .I3(\data_out_frame[20] [4]), .O(n42924));
    defparam i1_2_lut_3_lut_4_lut_adj_1346.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1347 (.I0(\data_out_frame[20] [5]), .I1(n44037), 
            .I2(\data_out_frame[20] [6]), .I3(n38980), .O(n44064));
    defparam i2_3_lut_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1348 (.I0(\data_out_frame[20] [4]), .I1(n39432), 
            .I2(n39012), .I3(\data_out_frame[20] [3]), .O(n23309));
    defparam i1_2_lut_3_lut_4_lut_adj_1348.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1349 (.I0(\data_out_frame[20] [3]), .I1(n39012), 
            .I2(n38931), .I3(\data_out_frame[20] [2]), .O(n22958));
    defparam i1_2_lut_3_lut_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1350 (.I0(\data_out_frame[20] [2]), .I1(n38931), 
            .I2(n39334), .I3(\data_out_frame[20] [1]), .O(n42897));
    defparam i1_2_lut_3_lut_4_lut_adj_1350.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(\data_out_frame[20] [1]), .I1(n39334), 
            .I2(n43062), .I3(GND_net), .O(n43063));
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1352 (.I0(\data_out_frame[19] [3]), .I1(n44450), 
            .I2(n42936), .I3(\data_out_frame[16] [6]), .O(n44323));
    defparam i2_3_lut_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1353 (.I0(\data_out_frame[19] [3]), .I1(n44450), 
            .I2(n43111), .I3(n38926), .O(n44212));
    defparam i2_3_lut_4_lut_adj_1353.LUT_INIT = 16'h9669;
    SB_LUT4 select_278_Select_0_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [0]), .O(n3_adj_3253));
    defparam select_278_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_1_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_3235));
    defparam select_278_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_2_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_3233));
    defparam select_278_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_3_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_3232));
    defparam select_278_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_adj_1354 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n21084));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1354.LUT_INIT = 16'h9696;
    SB_LUT4 select_278_Select_4_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_3231));
    defparam select_278_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_5_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_3230));
    defparam select_278_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_6_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_3229));
    defparam select_278_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i3_4_lut_adj_1355 (.I0(n1512), .I1(n42826), .I2(n43277), .I3(n43121), 
            .O(n42987));
    defparam i3_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 select_278_Select_7_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_3227));
    defparam select_278_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1356 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42939));   // verilog/coms.v(82[17:63])
    defparam i1_2_lut_adj_1356.LUT_INIT = 16'h6666;
    SB_LUT4 select_278_Select_8_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_3225));
    defparam select_278_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_4_lut_adj_1357 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[3] [5]), .O(Kp_23__N_458));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1358 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n23522));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1358.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1359 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43202));
    defparam i1_2_lut_adj_1359.LUT_INIT = 16'h6666;
    SB_LUT4 select_278_Select_9_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_3223));
    defparam select_278_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_278_Select_10_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_3221));
    defparam select_278_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1360 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23371));
    defparam i1_2_lut_adj_1360.LUT_INIT = 16'h6666;
    SB_LUT4 select_278_Select_11_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_3220));
    defparam select_278_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1361 (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(n43008), .I3(\data_in_frame[6] [3]), .O(n42958));   // verilog/coms.v(69[16:41])
    defparam i1_2_lut_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1362 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n23313));
    defparam i1_2_lut_adj_1362.LUT_INIT = 16'h6666;
    SB_LUT4 select_278_Select_12_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_3219));
    defparam select_278_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_adj_1363 (.I0(\data_out_frame[7] [2]), .I1(n23485), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n43292));
    defparam i2_3_lut_adj_1363.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1364 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42948));
    defparam i1_2_lut_adj_1364.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1365 (.I0(\data_out_frame[6] [5]), .I1(n43292), 
            .I2(GND_net), .I3(GND_net), .O(n42964));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1365.LUT_INIT = 16'h6666;
    SB_LUT4 select_278_Select_13_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_3218));
    defparam select_278_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1366 (.I0(\data_out_frame[13] [2]), .I1(n22664), 
            .I2(GND_net), .I3(GND_net), .O(n42932));   // verilog/coms.v(82[17:63])
    defparam i1_2_lut_adj_1366.LUT_INIT = 16'h6666;
    SB_LUT4 select_278_Select_14_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_3217));
    defparam select_278_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i7_4_lut_adj_1367 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[8] [4]), 
            .I2(n42932), .I3(\data_out_frame[18] [0]), .O(n18_adj_3356));
    defparam i7_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n6_adj_3187));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1369 (.I0(n23528), .I1(n38906), .I2(n21084), 
            .I3(n4_c), .O(n39675));
    defparam i1_2_lut_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 select_278_Select_15_i3_2_lut_4_lut (.I0(n28588), .I1(n22513), 
            .I2(n22520), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_3216));
    defparam select_278_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_4_lut_adj_1370 (.I0(n23528), .I1(n38906), .I2(n21084), 
            .I3(n23446), .O(n39661));
    defparam i1_2_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1371 (.I0(n23371), .I1(n18_adj_3356), .I2(n42752), 
            .I3(n43202), .O(n20_adj_3357));
    defparam i9_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1372 (.I0(n42964), .I1(n20_adj_3357), .I2(n16_adj_3322), 
            .I3(n42865), .O(n23326));
    defparam i10_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1373 (.I0(n42974), .I1(n42987), .I2(n38984), 
            .I3(n22187), .O(n12_adj_3358));
    defparam i5_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1374 (.I0(n38994), .I1(n12_adj_3358), .I2(n43215), 
            .I3(n22664), .O(n38920));
    defparam i6_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1375 (.I0(n38920), .I1(n23326), .I2(GND_net), 
            .I3(GND_net), .O(n38931));
    defparam i1_2_lut_adj_1375.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1376 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[20] [4]), 
            .I2(n38900), .I3(\data_out_frame[20] [3]), .O(n12_adj_3359));   // verilog/coms.v(68[16:27])
    defparam i5_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1377 (.I0(\data_out_frame[20] [5]), .I1(n12_adj_3359), 
            .I2(n42916), .I3(\data_out_frame[20] [1]), .O(n39004));   // verilog/coms.v(68[16:27])
    defparam i6_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1378 (.I0(\data_out_frame[18] [3]), .I1(n39601), 
            .I2(n22967), .I3(n23317), .O(n10_adj_3292));
    defparam i4_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1379 (.I0(n38920), .I1(\data_out_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3360));
    defparam i2_2_lut_adj_1379.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1380 (.I0(n7_adj_3360), .I1(n44449), .I2(\data_out_frame[16] [1]), 
            .I3(n39601), .O(n39012));
    defparam i4_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1381 (.I0(\data_in_frame[8] [5]), .I1(n10_adj_3157), 
            .I2(\data_in_frame[11] [1]), .I3(n10_adj_3142), .O(n22891));   // verilog/coms.v(69[16:41])
    defparam i5_3_lut_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1382 (.I0(n39012), .I1(n44037), .I2(n39004), 
            .I3(n38931), .O(n12_adj_3361));
    defparam i5_4_lut_adj_1382.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1383 (.I0(n39432), .I1(n12_adj_3361), .I2(n39334), 
            .I3(n38980), .O(n39599));
    defparam i6_4_lut_adj_1383.LUT_INIT = 16'h6996;
    uart_tx tx (.n23847(n23847), .clk32MHz(clk32MHz), .n23850(n23850), 
            .n23853(n23853), .n23856(n23856), .n23859(n23859), .n23862(n23862), 
            .n23865(n23865), .n23868(n23868), .n23872(n23872), .r_Bit_Index({r_Bit_Index}), 
            .n23875(n23875), .n23845(n23845), .n23848(n23848), .tx_data({tx_data}), 
            .n23851(n23851), .n23915(n23915), .n23918(n23918), .n23854(n23854), 
            .n23857(n23857), .n23860(n23860), .n23863(n23863), .\r_SM_Main_2__N_2747[0] (r_SM_Main_2__N_2747[0]), 
            .GND_net(GND_net), .n23866(n23866), .n23913(n23913), .VCC_net(VCC_net), 
            .tx_o(tx_o), .n23655(n23655), .n23785(n23785), .n4038(n4038), 
            .n23914(n23914), .tx_enable(tx_enable), .n29027(n29027), .tx_transmit_N_2639(tx_transmit_N_2639), 
            .n745(n745)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(104[10:70])
    uart_rx rx (.clk32MHz(clk32MHz), .n23878(n23878), .r_Bit_Index({r_Bit_Index_adj_9}), 
            .n23881(n23881), .n24453(n24453), .rx_data({rx_data}), .VCC_net(VCC_net), 
            .rx_data_ready(rx_data_ready), .n29023(n29023), .r_SM_Main({\r_SM_Main[2] , 
            \r_SM_Main[1] , Open_14}), .r_Rx_Data(r_Rx_Data), .LED_c(LED_c), 
            .GND_net(GND_net), .n24391(n24391), .n23888(n23888), .n23887(n23887), 
            .n23886(n23886), .n23885(n23885), .n23884(n23884), .n23883(n23883), 
            .n23882(n23882), .n23817(n23817), .n46591(n46591), .n22534(n22534), 
            .n4(n4), .n28989(n28989), .n28517(n28517), .n4_adj_1(n4_adj_7), 
            .n4_adj_2(n4_adj_8), .n23649(n23649), .n23783(n23783), .n4016(n4016), 
            .n22539(n22539), .n1(n1), .n46590(n46590)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(90[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n23847, clk32MHz, n23850, n23853, n23856, n23859, 
            n23862, n23865, n23868, n23872, r_Bit_Index, n23875, 
            n23845, n23848, tx_data, n23851, n23915, n23918, n23854, 
            n23857, n23860, n23863, \r_SM_Main_2__N_2747[0] , GND_net, 
            n23866, n23913, VCC_net, tx_o, n23655, n23785, n4038, 
            n23914, tx_enable, n29027, tx_transmit_N_2639, n745) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n23847;
    input clk32MHz;
    input n23850;
    input n23853;
    input n23856;
    input n23859;
    input n23862;
    input n23865;
    input n23868;
    input n23872;
    output [2:0]r_Bit_Index;
    input n23875;
    output n23845;
    output n23848;
    input [7:0]tx_data;
    output n23851;
    input n23915;
    input n23918;
    output n23854;
    output n23857;
    output n23860;
    output n23863;
    input \r_SM_Main_2__N_2747[0] ;
    input GND_net;
    output n23866;
    output n23913;
    input VCC_net;
    output tx_o;
    output n23655;
    output n23785;
    output n4038;
    output n23914;
    output tx_enable;
    input n29027;
    output tx_transmit_N_2639;
    output n745;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n42504;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    
    wire n36507, n36506, n20351;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n36505, n36504, n36503, n36502, n36501, n5, n36500, n44742, 
        n44743, n49390, n44686, n44685, o_Tx_Serial_N_2775, n43619, 
        n23824, n25739, tx_active, n10;
    wire [2:0]r_SM_Main_2__N_2744;
    
    wire n29007, n12, n23583, n28903, n19663, n38461, n10_adj_3109, 
        n44628, n9, n44626;
    
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .D(n23847));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n23850));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n23853));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n23856));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n23859));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n23862));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n23865));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n23868));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n23872));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n23875));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n42504));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[8]), 
            .I2(r_SM_Main[2]), .I3(n36507), .O(n23845)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_59_9_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[7]), 
            .I2(r_SM_Main[2]), .I3(n36506), .O(n23848)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hA3AC;
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n20351), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_9 (.CI(n36506), .I0(r_Clock_Count[7]), .I1(r_SM_Main[2]), 
            .CO(n36507));
    SB_LUT4 add_59_8_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[6]), 
            .I2(r_SM_Main[2]), .I3(n36505), .O(n23851)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hA3AC;
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n23915));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n23918));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_8 (.CI(n36505), .I0(r_Clock_Count[6]), .I1(r_SM_Main[2]), 
            .CO(n36506));
    SB_LUT4 add_59_7_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[5]), 
            .I2(r_SM_Main[2]), .I3(n36504), .O(n23854)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_7 (.CI(n36504), .I0(r_Clock_Count[5]), .I1(r_SM_Main[2]), 
            .CO(n36505));
    SB_LUT4 add_59_6_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[4]), 
            .I2(r_SM_Main[2]), .I3(n36503), .O(n23857)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_6 (.CI(n36503), .I0(r_Clock_Count[4]), .I1(r_SM_Main[2]), 
            .CO(n36504));
    SB_LUT4 add_59_5_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[3]), 
            .I2(r_SM_Main[2]), .I3(n36502), .O(n23860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_5 (.CI(n36502), .I0(r_Clock_Count[3]), .I1(r_SM_Main[2]), 
            .CO(n36503));
    SB_LUT4 add_59_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[2]), 
            .I2(r_SM_Main[2]), .I3(n36501), .O(n23863)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_4 (.CI(n36501), .I0(r_Clock_Count[2]), .I1(r_SM_Main[2]), 
            .CO(n36502));
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_2747[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 add_59_3_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[1]), 
            .I2(r_SM_Main[2]), .I3(n36500), .O(n23866)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_3 (.CI(n36500), .I0(r_Clock_Count[1]), .I1(r_SM_Main[2]), 
            .CO(n36501));
    SB_LUT4 add_59_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[0]), 
            .I2(r_SM_Main[2]), .I3(VCC_net), .O(n23913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(r_SM_Main[2]), 
            .CO(n36500));
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n44742), 
            .I2(n44743), .I3(r_Bit_Index[2]), .O(n49390));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49390_bdd_4_lut (.I0(n49390), .I1(n44686), .I2(n44685), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_2775));
    defparam n49390_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n20351), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n20351), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n20351), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n20351), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n20351), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n20351), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n20351), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n43619));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n23824));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n25739));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n10));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i15599_2_lut (.I0(r_SM_Main_2__N_2744[1]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29007));
    defparam i15599_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_2775), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n12));
    defparam i26_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i25_3_lut (.I0(n12), .I1(tx_o), .I2(r_SM_Main[2]), .I3(GND_net), 
            .O(n10));
    defparam i25_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i2_4_lut (.I0(n5), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), .I3(n29007), 
            .O(n23583));
    defparam i2_4_lut.LUT_INIT = 16'h3202;
    SB_LUT4 i12324_3_lut (.I0(n23583), .I1(r_SM_Main[1]), .I2(tx_active), 
            .I3(GND_net), .O(n25739));   // verilog/uart_tx.v(31[16:25])
    defparam i12324_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i6357_4_lut (.I0(\r_SM_Main_2__N_2747[0] ), .I1(n28903), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_2744[1]), .O(n19663));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i6357_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n19663), .I2(r_SM_Main_2__N_2744[1]), 
            .I3(r_SM_Main[0]), .O(n23824));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n28903));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), .I2(n38461), 
            .I3(r_Clock_Count[8]), .O(n10_adj_3109));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10_adj_3109), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(r_SM_Main_2__N_2744[1]));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_826 (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_2744[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n23655));
    defparam i2_4_lut_adj_826.LUT_INIT = 16'h0405;
    SB_LUT4 i10367_3_lut (.I0(n23655), .I1(n28903), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n23785));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10367_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1123_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4038));   // verilog/uart_tx.v(98[36:51])
    defparam i1123_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), .I2(r_Clock_Count[3]), 
            .I3(r_Clock_Count[2]), .O(n38461));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i29116_2_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[4]), 
            .I2(GND_net), .I3(GND_net), .O(n44628));
    defparam i29116_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_827 (.I0(r_Clock_Count[6]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n9));
    defparam i2_3_lut_adj_827.LUT_INIT = 16'h5454;
    SB_LUT4 i29114_3_lut (.I0(r_Clock_Count[7]), .I1(n38461), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n44626));
    defparam i29114_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_828 (.I0(r_SM_Main[2]), .I1(n44626), .I2(n9), 
            .I3(n44628), .O(n23914));   // verilog/uart_tx.v(31[16:25])
    defparam i1_4_lut_adj_828.LUT_INIT = 16'haaba;
    SB_LUT4 i29173_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n44685));
    defparam i29173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29174_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n44686));
    defparam i29174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29231_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n44743));
    defparam i29231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29230_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n44742));
    defparam i29230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main_2__N_2744[1]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n43619));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_2744[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n42504));   // verilog/uart_tx.v(31[16:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1540;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_2747[0] ), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n20351));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i33795_2_lut_3_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_2747[0] ), 
            .I2(n29027), .I3(GND_net), .O(tx_transmit_N_2639));
    defparam i33795_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i233_2_lut_3_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_2747[0] ), 
            .I2(n29027), .I3(GND_net), .O(n745));
    defparam i233_2_lut_3_lut.LUT_INIT = 16'hefef;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (clk32MHz, n23878, r_Bit_Index, n23881, n24453, rx_data, 
            VCC_net, rx_data_ready, n29023, r_SM_Main, r_Rx_Data, 
            LED_c, GND_net, n24391, n23888, n23887, n23886, n23885, 
            n23884, n23883, n23882, n23817, n46591, n22534, n4, 
            n28989, n28517, n4_adj_1, n4_adj_2, n23649, n23783, 
            n4016, n22539, n1, n46590) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input n23878;
    output [2:0]r_Bit_Index;
    input n23881;
    input n24453;
    output [7:0]rx_data;
    input VCC_net;
    output rx_data_ready;
    input n29023;
    output [2:0]r_SM_Main;
    output r_Rx_Data;
    input LED_c;
    input GND_net;
    input n24391;
    input n23888;
    input n23887;
    input n23886;
    input n23885;
    input n23884;
    input n23883;
    input n23882;
    input n23817;
    output n46591;
    output n22534;
    output n4;
    output n28989;
    output n28517;
    output n4_adj_1;
    output n4_adj_2;
    output n23649;
    output n23783;
    output n4016;
    output n22539;
    output n1;
    output n46590;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n23820;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n23827, n42138, n23835, n23838, n23841, n23844, n42096, 
        r_Rx_Data_R, n23912, n46472, n43339, n30103, n4_c;
    wire [2:0]r_SM_Main_2__N_2673;
    
    wire n42675, n46475, n36499, n108, n46474, n36498, n46618, 
        n36497, n46471, n36496, n46473, n36495, n46476, n36494, 
        n46470, n36493;
    wire [2:0]r_SM_Main_c;   // verilog/uart_rx.v(36[17:26])
    
    wire n22386, n28897, n44585, n42732, n11, n46627, n46625, 
        n38;
    wire [2:0]r_SM_Main_2__N_2679;
    
    wire n43887, n23570;
    
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n23820));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n23827));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n42138));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n23835));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n23838));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n23841));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n23844));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n23878));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n23881));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n24453));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n42096));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n29023));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(LED_c));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n23912));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i16771_3_lut (.I0(r_Clock_Count[0]), .I1(n46472), .I2(n43339), 
            .I3(GND_net), .O(n23912));
    defparam i16771_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n24391));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i15498_3_lut_4_lut (.I0(r_Clock_Count[0]), .I1(n30103), .I2(n4_c), 
            .I3(r_Clock_Count[3]), .O(r_SM_Main_2__N_2673[2]));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15498_3_lut_4_lut.LUT_INIT = 16'hf8f0;
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_2673[2]), 
            .R(n42675));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_9_lut (.I0(n108), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n36499), .O(n46475)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(n108), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n36498), .O(n46474)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_8 (.CI(n36498), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n36499));
    SB_LUT4 add_62_7_lut (.I0(n108), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n36497), .O(n46618)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_7 (.CI(n36497), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n36498));
    SB_LUT4 add_62_6_lut (.I0(n108), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n36496), .O(n46471)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n36496), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n36497));
    SB_LUT4 add_62_5_lut (.I0(n108), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n36495), .O(n46473)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_5 (.CI(n36495), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n36496));
    SB_LUT4 add_62_4_lut (.I0(n108), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n36494), .O(n46476)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_4 (.CI(n36494), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n36495));
    SB_LUT4 add_62_3_lut (.I0(n108), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n36493), .O(n46470)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_3 (.CI(n36493), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n36494));
    SB_LUT4 add_62_2_lut (.I0(n108), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n46472)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n36493));
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n23888));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n23887));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n23886));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n23885));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n23884));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n23883));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n23882));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n23817));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i31789_2_lut (.I0(r_SM_Main_2__N_2673[2]), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46591));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i31789_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main_2__N_2673[2]), .O(n22386));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut (.I0(r_Bit_Index[0]), .I1(n22386), .I2(GND_net), 
            .I3(GND_net), .O(n22534));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_77_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_77_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n28897), .I1(r_SM_Main_2__N_2673[2]), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n28989));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 i15118_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n28517));
    defparam i15118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_73_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_73_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_75_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_75_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n28897));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_2673[2]), .I2(r_SM_Main_c[0]), 
            .I3(r_SM_Main[1]), .O(n23649));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i10365_3_lut (.I0(n23649), .I1(n28897), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n23783));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10365_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1101_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4016));   // verilog/uart_rx.v(102[36:51])
    defparam i1101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16759_3_lut (.I0(r_Clock_Count[1]), .I1(n46470), .I2(n43339), 
            .I3(GND_net), .O(n23844));
    defparam i16759_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16789_3_lut (.I0(r_Clock_Count[2]), .I1(n46476), .I2(n43339), 
            .I3(GND_net), .O(n23841));
    defparam i16789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_821 (.I0(n22386), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n22539));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_821.LUT_INIT = 16'hbbbb;
    SB_LUT4 i16775_3_lut (.I0(r_Clock_Count[3]), .I1(n46473), .I2(n43339), 
            .I3(GND_net), .O(n23838));
    defparam i16775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16765_3_lut (.I0(r_Clock_Count[4]), .I1(n46471), .I2(n43339), 
            .I3(GND_net), .O(n23835));
    defparam i16765_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_3_lut (.I0(r_Clock_Count[5]), .I1(n46618), .I2(n43339), 
            .I3(GND_net), .O(n42138));
    defparam i11_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16779_3_lut (.I0(r_Clock_Count[6]), .I1(n46474), .I2(n43339), 
            .I3(GND_net), .O(n23827));
    defparam i16779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29075_2_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[3]), 
            .I2(GND_net), .I3(GND_net), .O(n44585));
    defparam i29075_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(r_Rx_Data), .I1(r_Clock_Count[4]), .I2(n42732), 
            .I3(GND_net), .O(n11));
    defparam i3_3_lut.LUT_INIT = 16'h3131;
    SB_LUT4 i31790_4_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[5]), 
            .I2(n30103), .I3(r_Clock_Count[0]), .O(n46627));
    defparam i31790_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i31472_4_lut (.I0(n46627), .I1(r_SM_Main_c[0]), .I2(n11), 
            .I3(n44585), .O(n46625));
    defparam i31472_4_lut.LUT_INIT = 16'h33b3;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n46625), .I2(r_SM_Main_2__N_2673[2]), 
            .I3(r_SM_Main[1]), .O(n38));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1_2_lut_adj_822 (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[1]), 
            .I2(GND_net), .I3(GND_net), .O(n30103));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_822.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_823 (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(r_Clock_Count[4]), .O(n4_c));
    defparam i1_4_lut_adj_823.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_824 (.I0(r_Clock_Count[3]), .I1(n42732), .I2(GND_net), 
            .I3(GND_net), .O(r_SM_Main_2__N_2679[0]));   // verilog/uart_rx.v(68[17:52])
    defparam i1_2_lut_adj_824.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_825 (.I0(r_SM_Main[1]), .I1(r_SM_Main_2__N_2679[0]), 
            .I2(r_Rx_Data), .I3(r_SM_Main_c[0]), .O(n43887));
    defparam i3_4_lut_adj_825.LUT_INIT = 16'h1000;
    SB_LUT4 i27837_3_lut (.I0(r_SM_Main[2]), .I1(n38), .I2(n43887), .I3(GND_net), 
            .O(n43339));
    defparam i27837_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i16783_3_lut (.I0(r_Clock_Count[7]), .I1(n46475), .I2(n43339), 
            .I3(GND_net), .O(n23820));
    defparam i16783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33803_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_c[0]), 
            .I3(GND_net), .O(n42675));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i33803_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_2673[2]), 
            .I3(r_SM_Main_c[0]), .O(n23570));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n23570), 
            .I3(rx_data_ready), .O(n42096));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i39_1_lut_4_lut (.I0(r_SM_Main[2]), .I1(n46625), .I2(r_SM_Main_2__N_2673[2]), 
            .I3(r_SM_Main[1]), .O(n108));
    defparam i39_1_lut_4_lut.LUT_INIT = 16'hafbb;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_4_lut (.I0(r_Rx_Data), .I1(r_Clock_Count[3]), 
            .I2(n42732), .I3(r_SM_Main_c[0]), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_4_lut.LUT_INIT = 16'hfc55;
    SB_LUT4 i31492_3_lut_4_lut (.I0(r_SM_Main_c[0]), .I1(r_Clock_Count[3]), 
            .I2(n42732), .I3(r_Rx_Data), .O(n46590));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i31492_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), 
            .I2(r_Clock_Count[1]), .I3(n4_c), .O(n42732));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n24406, encoder1_position, clk32MHz, 
            n24405, n24404, n24422, n24421, n24420, n24419, n24418, 
            n24417, n24416, n24415, n24414, n24413, n24412, n24411, 
            n24410, n24409, n24408, n24407, n24403, data_o, n24402, 
            n24401, n24388, count_enable, n2242, GND_net, n23815, 
            n24452, PIN_23_c_0, reg_B, PIN_24_c_1, n23821, n44154) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n24406;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n24405;
    input n24404;
    input n24422;
    input n24421;
    input n24420;
    input n24419;
    input n24418;
    input n24417;
    input n24416;
    input n24415;
    input n24414;
    input n24413;
    input n24412;
    input n24411;
    input n24410;
    input n24409;
    input n24408;
    input n24407;
    input n24403;
    output [1:0]data_o;
    input n24402;
    input n24401;
    input n24388;
    output count_enable;
    output [23:0]n2242;
    input GND_net;
    input n23815;
    input n24452;
    input PIN_23_c_0;
    output [1:0]reg_B;
    input PIN_24_c_1;
    input n23821;
    output n44154;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire B_delayed, A_delayed, n2234, n36598, n36597, n36596, n36595, 
        n36594, n36593, n36592, n36591, n36590, n36589, n36588, 
        n36587, n36586, n36585, n36584, n36583, n36582, n36581, 
        n36580, n36579, n36578, n36577, n36576, count_direction, 
        n36575;
    
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n24406));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n24405));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n24404));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n24422));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n24421));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n24420));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n24419));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n24418));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n24417));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n24416));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n24415));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n24414));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n24413));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n24412));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n24411));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n24410));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n24409));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n24408));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n24407));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n24403));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n24402));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n24401));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n24388));   // quad.v(35[10] 41[6])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_524_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2234), 
            .I3(n36598), .O(n2242[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_524_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2234), 
            .I3(n36597), .O(n2242[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_24 (.CI(n36597), .I0(encoder1_position[22]), .I1(n2234), 
            .CO(n36598));
    SB_LUT4 add_524_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2234), 
            .I3(n36596), .O(n2242[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_23 (.CI(n36596), .I0(encoder1_position[21]), .I1(n2234), 
            .CO(n36597));
    SB_LUT4 add_524_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2234), 
            .I3(n36595), .O(n2242[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_22 (.CI(n36595), .I0(encoder1_position[20]), .I1(n2234), 
            .CO(n36596));
    SB_LUT4 add_524_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2234), 
            .I3(n36594), .O(n2242[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_21 (.CI(n36594), .I0(encoder1_position[19]), .I1(n2234), 
            .CO(n36595));
    SB_LUT4 add_524_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2234), 
            .I3(n36593), .O(n2242[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_20 (.CI(n36593), .I0(encoder1_position[18]), .I1(n2234), 
            .CO(n36594));
    SB_LUT4 add_524_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2234), 
            .I3(n36592), .O(n2242[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_19 (.CI(n36592), .I0(encoder1_position[17]), .I1(n2234), 
            .CO(n36593));
    SB_LUT4 add_524_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2234), 
            .I3(n36591), .O(n2242[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_18 (.CI(n36591), .I0(encoder1_position[16]), .I1(n2234), 
            .CO(n36592));
    SB_LUT4 add_524_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2234), 
            .I3(n36590), .O(n2242[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_17 (.CI(n36590), .I0(encoder1_position[15]), .I1(n2234), 
            .CO(n36591));
    SB_LUT4 add_524_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2234), 
            .I3(n36589), .O(n2242[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_16 (.CI(n36589), .I0(encoder1_position[14]), .I1(n2234), 
            .CO(n36590));
    SB_LUT4 add_524_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2234), 
            .I3(n36588), .O(n2242[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_15 (.CI(n36588), .I0(encoder1_position[13]), .I1(n2234), 
            .CO(n36589));
    SB_LUT4 add_524_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2234), 
            .I3(n36587), .O(n2242[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_14 (.CI(n36587), .I0(encoder1_position[12]), .I1(n2234), 
            .CO(n36588));
    SB_LUT4 add_524_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2234), 
            .I3(n36586), .O(n2242[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_13 (.CI(n36586), .I0(encoder1_position[11]), .I1(n2234), 
            .CO(n36587));
    SB_LUT4 add_524_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2234), 
            .I3(n36585), .O(n2242[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_12 (.CI(n36585), .I0(encoder1_position[10]), .I1(n2234), 
            .CO(n36586));
    SB_LUT4 add_524_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2234), 
            .I3(n36584), .O(n2242[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_11 (.CI(n36584), .I0(encoder1_position[9]), .I1(n2234), 
            .CO(n36585));
    SB_LUT4 add_524_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2234), 
            .I3(n36583), .O(n2242[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_10 (.CI(n36583), .I0(encoder1_position[8]), .I1(n2234), 
            .CO(n36584));
    SB_LUT4 add_524_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2234), 
            .I3(n36582), .O(n2242[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_9 (.CI(n36582), .I0(encoder1_position[7]), .I1(n2234), 
            .CO(n36583));
    SB_LUT4 add_524_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2234), 
            .I3(n36581), .O(n2242[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_8 (.CI(n36581), .I0(encoder1_position[6]), .I1(n2234), 
            .CO(n36582));
    SB_LUT4 add_524_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2234), 
            .I3(n36580), .O(n2242[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_7 (.CI(n36580), .I0(encoder1_position[5]), .I1(n2234), 
            .CO(n36581));
    SB_LUT4 add_524_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2234), 
            .I3(n36579), .O(n2242[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_6 (.CI(n36579), .I0(encoder1_position[4]), .I1(n2234), 
            .CO(n36580));
    SB_LUT4 add_524_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2234), 
            .I3(n36578), .O(n2242[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_5 (.CI(n36578), .I0(encoder1_position[3]), .I1(n2234), 
            .CO(n36579));
    SB_LUT4 add_524_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2234), 
            .I3(n36577), .O(n2242[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_4 (.CI(n36577), .I0(encoder1_position[2]), .I1(n2234), 
            .CO(n36578));
    SB_LUT4 add_524_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2234), 
            .I3(n36576), .O(n2242[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_3 (.CI(n36576), .I0(encoder1_position[1]), .I1(n2234), 
            .CO(n36577));
    SB_LUT4 add_524_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n36575), .O(n2242[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_524_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_524_2 (.CI(n36575), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n36576));
    SB_CARRY add_524_1 (.CI(GND_net), .I0(n2234), .I1(n2234), .CO(n36575));
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n23815));   // quad.v(35[10] 41[6])
    SB_LUT4 i786_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2234));   // quad.v(37[5] 40[8])
    defparam i786_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    \grp_debouncer(2,5)  debounce (.n24452(n24452), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .PIN_23_c_0(PIN_23_c_0), .reg_B({reg_B}), .PIN_24_c_1(PIN_24_c_1), 
            .n23821(n23821), .n44154(n44154), .GND_net(GND_net)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n24452, data_o, clk32MHz, PIN_23_c_0, reg_B, 
            PIN_24_c_1, n23821, n44154, GND_net) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n24452;
    output [1:0]data_o;
    input clk32MHz;
    input PIN_23_c_0;
    output [1:0]reg_B;
    input PIN_24_c_1;
    input n23821;
    output n44154;
    input GND_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3104, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n24452));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_23_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_24_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1051__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1051__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n23821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1051__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n44154));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i22884_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22884_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22877_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22877_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n44154), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22875_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22875_1_lut.LUT_INIT = 16'h5555;
    
endmodule
