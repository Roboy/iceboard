// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Feb 24 2020 16:03:38

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    TX,
    SDA,
    SCL,
    RX,
    NEOPXL,
    LED,
    INLC,
    INLB,
    INLA,
    INHC,
    INHB,
    INHA,
    HALL3,
    HALL2,
    HALL1,
    FAULT_N,
    ENCODER1_B,
    ENCODER1_A,
    ENCODER0_B,
    ENCODER0_A,
    DE,
    CS_MISO,
    CS_CLK,
    CS,
    CLK);

    inout USBPU;
    inout TX;
    inout SDA;
    inout SCL;
    inout RX;
    output NEOPXL;
    output LED;
    inout INLC;
    inout INLB;
    inout INLA;
    inout INHC;
    inout INHB;
    inout INHA;
    inout HALL3;
    inout HALL2;
    inout HALL1;
    inout FAULT_N;
    inout ENCODER1_B;
    inout ENCODER1_A;
    inout ENCODER0_B;
    inout ENCODER0_A;
    inout DE;
    inout CS_MISO;
    inout CS_CLK;
    inout CS;
    input CLK;

    wire N__47950;
    wire N__47949;
    wire N__47948;
    wire N__47941;
    wire N__47940;
    wire N__47939;
    wire N__47932;
    wire N__47931;
    wire N__47930;
    wire N__47923;
    wire N__47922;
    wire N__47921;
    wire N__47914;
    wire N__47913;
    wire N__47912;
    wire N__47905;
    wire N__47904;
    wire N__47903;
    wire N__47896;
    wire N__47895;
    wire N__47894;
    wire N__47887;
    wire N__47886;
    wire N__47885;
    wire N__47878;
    wire N__47877;
    wire N__47876;
    wire N__47869;
    wire N__47868;
    wire N__47867;
    wire N__47860;
    wire N__47859;
    wire N__47858;
    wire N__47851;
    wire N__47850;
    wire N__47849;
    wire N__47842;
    wire N__47841;
    wire N__47840;
    wire N__47833;
    wire N__47832;
    wire N__47831;
    wire N__47824;
    wire N__47823;
    wire N__47822;
    wire N__47815;
    wire N__47814;
    wire N__47813;
    wire N__47806;
    wire N__47805;
    wire N__47804;
    wire N__47797;
    wire N__47796;
    wire N__47795;
    wire N__47788;
    wire N__47787;
    wire N__47786;
    wire N__47779;
    wire N__47778;
    wire N__47777;
    wire N__47770;
    wire N__47769;
    wire N__47768;
    wire N__47761;
    wire N__47760;
    wire N__47759;
    wire N__47752;
    wire N__47751;
    wire N__47750;
    wire N__47743;
    wire N__47742;
    wire N__47741;
    wire N__47734;
    wire N__47733;
    wire N__47732;
    wire N__47725;
    wire N__47724;
    wire N__47723;
    wire N__47706;
    wire N__47703;
    wire N__47700;
    wire N__47697;
    wire N__47696;
    wire N__47695;
    wire N__47694;
    wire N__47693;
    wire N__47690;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47677;
    wire N__47676;
    wire N__47675;
    wire N__47674;
    wire N__47673;
    wire N__47672;
    wire N__47669;
    wire N__47668;
    wire N__47667;
    wire N__47666;
    wire N__47665;
    wire N__47664;
    wire N__47663;
    wire N__47660;
    wire N__47659;
    wire N__47658;
    wire N__47657;
    wire N__47654;
    wire N__47651;
    wire N__47648;
    wire N__47647;
    wire N__47646;
    wire N__47643;
    wire N__47642;
    wire N__47641;
    wire N__47638;
    wire N__47637;
    wire N__47636;
    wire N__47635;
    wire N__47632;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47624;
    wire N__47621;
    wire N__47618;
    wire N__47611;
    wire N__47610;
    wire N__47607;
    wire N__47604;
    wire N__47601;
    wire N__47600;
    wire N__47599;
    wire N__47598;
    wire N__47595;
    wire N__47594;
    wire N__47591;
    wire N__47590;
    wire N__47587;
    wire N__47586;
    wire N__47585;
    wire N__47584;
    wire N__47583;
    wire N__47582;
    wire N__47581;
    wire N__47578;
    wire N__47577;
    wire N__47570;
    wire N__47563;
    wire N__47560;
    wire N__47555;
    wire N__47550;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47539;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47523;
    wire N__47520;
    wire N__47519;
    wire N__47518;
    wire N__47517;
    wire N__47516;
    wire N__47515;
    wire N__47514;
    wire N__47509;
    wire N__47506;
    wire N__47503;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47489;
    wire N__47488;
    wire N__47485;
    wire N__47484;
    wire N__47483;
    wire N__47482;
    wire N__47481;
    wire N__47480;
    wire N__47479;
    wire N__47478;
    wire N__47475;
    wire N__47470;
    wire N__47461;
    wire N__47460;
    wire N__47459;
    wire N__47456;
    wire N__47453;
    wire N__47450;
    wire N__47447;
    wire N__47444;
    wire N__47437;
    wire N__47432;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47415;
    wire N__47412;
    wire N__47407;
    wire N__47402;
    wire N__47397;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47380;
    wire N__47377;
    wire N__47372;
    wire N__47369;
    wire N__47368;
    wire N__47367;
    wire N__47364;
    wire N__47363;
    wire N__47360;
    wire N__47355;
    wire N__47350;
    wire N__47347;
    wire N__47344;
    wire N__47341;
    wire N__47336;
    wire N__47333;
    wire N__47330;
    wire N__47329;
    wire N__47326;
    wire N__47325;
    wire N__47324;
    wire N__47323;
    wire N__47318;
    wire N__47315;
    wire N__47308;
    wire N__47305;
    wire N__47302;
    wire N__47301;
    wire N__47300;
    wire N__47299;
    wire N__47296;
    wire N__47277;
    wire N__47272;
    wire N__47269;
    wire N__47264;
    wire N__47259;
    wire N__47256;
    wire N__47251;
    wire N__47234;
    wire N__47229;
    wire N__47226;
    wire N__47221;
    wire N__47218;
    wire N__47215;
    wire N__47208;
    wire N__47199;
    wire N__47194;
    wire N__47183;
    wire N__47176;
    wire N__47157;
    wire N__47156;
    wire N__47155;
    wire N__47154;
    wire N__47153;
    wire N__47150;
    wire N__47149;
    wire N__47148;
    wire N__47147;
    wire N__47146;
    wire N__47143;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47130;
    wire N__47127;
    wire N__47126;
    wire N__47125;
    wire N__47124;
    wire N__47123;
    wire N__47122;
    wire N__47121;
    wire N__47120;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47110;
    wire N__47107;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47085;
    wire N__47082;
    wire N__47079;
    wire N__47076;
    wire N__47073;
    wire N__47072;
    wire N__47069;
    wire N__47066;
    wire N__47061;
    wire N__47058;
    wire N__47053;
    wire N__47048;
    wire N__47043;
    wire N__47040;
    wire N__47039;
    wire N__47038;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47028;
    wire N__47025;
    wire N__47022;
    wire N__47019;
    wire N__47014;
    wire N__47005;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46990;
    wire N__46985;
    wire N__46982;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46950;
    wire N__46947;
    wire N__46944;
    wire N__46941;
    wire N__46938;
    wire N__46935;
    wire N__46934;
    wire N__46931;
    wire N__46928;
    wire N__46923;
    wire N__46922;
    wire N__46921;
    wire N__46920;
    wire N__46919;
    wire N__46918;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46913;
    wire N__46912;
    wire N__46911;
    wire N__46910;
    wire N__46909;
    wire N__46908;
    wire N__46907;
    wire N__46906;
    wire N__46905;
    wire N__46904;
    wire N__46903;
    wire N__46902;
    wire N__46901;
    wire N__46900;
    wire N__46899;
    wire N__46898;
    wire N__46897;
    wire N__46896;
    wire N__46895;
    wire N__46894;
    wire N__46893;
    wire N__46892;
    wire N__46891;
    wire N__46890;
    wire N__46889;
    wire N__46888;
    wire N__46887;
    wire N__46886;
    wire N__46885;
    wire N__46884;
    wire N__46883;
    wire N__46882;
    wire N__46881;
    wire N__46880;
    wire N__46879;
    wire N__46878;
    wire N__46877;
    wire N__46876;
    wire N__46875;
    wire N__46874;
    wire N__46873;
    wire N__46872;
    wire N__46871;
    wire N__46870;
    wire N__46869;
    wire N__46868;
    wire N__46867;
    wire N__46866;
    wire N__46865;
    wire N__46864;
    wire N__46863;
    wire N__46862;
    wire N__46861;
    wire N__46860;
    wire N__46859;
    wire N__46858;
    wire N__46857;
    wire N__46856;
    wire N__46855;
    wire N__46854;
    wire N__46853;
    wire N__46852;
    wire N__46851;
    wire N__46850;
    wire N__46849;
    wire N__46848;
    wire N__46847;
    wire N__46846;
    wire N__46845;
    wire N__46844;
    wire N__46843;
    wire N__46842;
    wire N__46841;
    wire N__46840;
    wire N__46839;
    wire N__46668;
    wire N__46665;
    wire N__46662;
    wire N__46659;
    wire N__46656;
    wire N__46653;
    wire N__46650;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46629;
    wire N__46626;
    wire N__46623;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46602;
    wire N__46599;
    wire N__46596;
    wire N__46593;
    wire N__46590;
    wire N__46587;
    wire N__46584;
    wire N__46581;
    wire N__46578;
    wire N__46575;
    wire N__46572;
    wire N__46571;
    wire N__46568;
    wire N__46567;
    wire N__46566;
    wire N__46565;
    wire N__46564;
    wire N__46563;
    wire N__46560;
    wire N__46559;
    wire N__46556;
    wire N__46555;
    wire N__46552;
    wire N__46549;
    wire N__46546;
    wire N__46545;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46533;
    wire N__46530;
    wire N__46527;
    wire N__46524;
    wire N__46523;
    wire N__46522;
    wire N__46517;
    wire N__46514;
    wire N__46513;
    wire N__46512;
    wire N__46511;
    wire N__46510;
    wire N__46509;
    wire N__46508;
    wire N__46505;
    wire N__46498;
    wire N__46491;
    wire N__46486;
    wire N__46481;
    wire N__46478;
    wire N__46473;
    wire N__46470;
    wire N__46467;
    wire N__46464;
    wire N__46459;
    wire N__46454;
    wire N__46451;
    wire N__46448;
    wire N__46445;
    wire N__46428;
    wire N__46425;
    wire N__46422;
    wire N__46419;
    wire N__46416;
    wire N__46413;
    wire N__46412;
    wire N__46411;
    wire N__46410;
    wire N__46409;
    wire N__46408;
    wire N__46407;
    wire N__46406;
    wire N__46405;
    wire N__46402;
    wire N__46397;
    wire N__46396;
    wire N__46393;
    wire N__46392;
    wire N__46387;
    wire N__46386;
    wire N__46385;
    wire N__46384;
    wire N__46383;
    wire N__46378;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46357;
    wire N__46352;
    wire N__46349;
    wire N__46346;
    wire N__46345;
    wire N__46344;
    wire N__46343;
    wire N__46338;
    wire N__46337;
    wire N__46336;
    wire N__46335;
    wire N__46332;
    wire N__46329;
    wire N__46324;
    wire N__46323;
    wire N__46322;
    wire N__46321;
    wire N__46320;
    wire N__46315;
    wire N__46308;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46289;
    wire N__46284;
    wire N__46281;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46269;
    wire N__46264;
    wire N__46257;
    wire N__46248;
    wire N__46233;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46203;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46166;
    wire N__46165;
    wire N__46162;
    wire N__46157;
    wire N__46152;
    wire N__46151;
    wire N__46148;
    wire N__46147;
    wire N__46146;
    wire N__46145;
    wire N__46144;
    wire N__46143;
    wire N__46142;
    wire N__46141;
    wire N__46140;
    wire N__46139;
    wire N__46138;
    wire N__46137;
    wire N__46136;
    wire N__46133;
    wire N__46132;
    wire N__46129;
    wire N__46126;
    wire N__46121;
    wire N__46118;
    wire N__46115;
    wire N__46112;
    wire N__46111;
    wire N__46110;
    wire N__46107;
    wire N__46104;
    wire N__46099;
    wire N__46098;
    wire N__46097;
    wire N__46096;
    wire N__46095;
    wire N__46094;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46067;
    wire N__46064;
    wire N__46061;
    wire N__46054;
    wire N__46049;
    wire N__46046;
    wire N__46041;
    wire N__46026;
    wire N__46019;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45995;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45987;
    wire N__45982;
    wire N__45981;
    wire N__45980;
    wire N__45979;
    wire N__45978;
    wire N__45975;
    wire N__45974;
    wire N__45973;
    wire N__45972;
    wire N__45971;
    wire N__45970;
    wire N__45965;
    wire N__45962;
    wire N__45961;
    wire N__45960;
    wire N__45959;
    wire N__45958;
    wire N__45957;
    wire N__45956;
    wire N__45953;
    wire N__45952;
    wire N__45949;
    wire N__45944;
    wire N__45941;
    wire N__45936;
    wire N__45931;
    wire N__45926;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45902;
    wire N__45901;
    wire N__45900;
    wire N__45899;
    wire N__45898;
    wire N__45893;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45856;
    wire N__45853;
    wire N__45848;
    wire N__45845;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45812;
    wire N__45811;
    wire N__45808;
    wire N__45803;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45789;
    wire N__45788;
    wire N__45787;
    wire N__45784;
    wire N__45781;
    wire N__45778;
    wire N__45773;
    wire N__45768;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45752;
    wire N__45751;
    wire N__45748;
    wire N__45745;
    wire N__45742;
    wire N__45735;
    wire N__45732;
    wire N__45729;
    wire N__45726;
    wire N__45723;
    wire N__45720;
    wire N__45717;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45707;
    wire N__45704;
    wire N__45701;
    wire N__45696;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45682;
    wire N__45681;
    wire N__45678;
    wire N__45675;
    wire N__45672;
    wire N__45671;
    wire N__45670;
    wire N__45669;
    wire N__45668;
    wire N__45665;
    wire N__45664;
    wire N__45661;
    wire N__45658;
    wire N__45655;
    wire N__45654;
    wire N__45653;
    wire N__45652;
    wire N__45651;
    wire N__45650;
    wire N__45649;
    wire N__45646;
    wire N__45645;
    wire N__45644;
    wire N__45643;
    wire N__45642;
    wire N__45641;
    wire N__45638;
    wire N__45635;
    wire N__45634;
    wire N__45631;
    wire N__45628;
    wire N__45627;
    wire N__45624;
    wire N__45619;
    wire N__45616;
    wire N__45615;
    wire N__45612;
    wire N__45611;
    wire N__45608;
    wire N__45605;
    wire N__45602;
    wire N__45599;
    wire N__45598;
    wire N__45597;
    wire N__45596;
    wire N__45593;
    wire N__45592;
    wire N__45589;
    wire N__45588;
    wire N__45587;
    wire N__45584;
    wire N__45581;
    wire N__45578;
    wire N__45575;
    wire N__45574;
    wire N__45571;
    wire N__45570;
    wire N__45569;
    wire N__45568;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45560;
    wire N__45557;
    wire N__45556;
    wire N__45553;
    wire N__45550;
    wire N__45547;
    wire N__45544;
    wire N__45539;
    wire N__45538;
    wire N__45535;
    wire N__45534;
    wire N__45531;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45515;
    wire N__45512;
    wire N__45509;
    wire N__45508;
    wire N__45507;
    wire N__45502;
    wire N__45499;
    wire N__45498;
    wire N__45497;
    wire N__45494;
    wire N__45493;
    wire N__45492;
    wire N__45489;
    wire N__45488;
    wire N__45487;
    wire N__45482;
    wire N__45481;
    wire N__45478;
    wire N__45475;
    wire N__45472;
    wire N__45467;
    wire N__45466;
    wire N__45463;
    wire N__45462;
    wire N__45461;
    wire N__45458;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45452;
    wire N__45449;
    wire N__45446;
    wire N__45443;
    wire N__45438;
    wire N__45431;
    wire N__45426;
    wire N__45419;
    wire N__45408;
    wire N__45403;
    wire N__45398;
    wire N__45393;
    wire N__45388;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45361;
    wire N__45356;
    wire N__45351;
    wire N__45348;
    wire N__45345;
    wire N__45338;
    wire N__45333;
    wire N__45316;
    wire N__45305;
    wire N__45302;
    wire N__45295;
    wire N__45270;
    wire N__45269;
    wire N__45268;
    wire N__45267;
    wire N__45264;
    wire N__45263;
    wire N__45262;
    wire N__45261;
    wire N__45258;
    wire N__45255;
    wire N__45254;
    wire N__45253;
    wire N__45252;
    wire N__45251;
    wire N__45250;
    wire N__45247;
    wire N__45240;
    wire N__45237;
    wire N__45234;
    wire N__45231;
    wire N__45226;
    wire N__45219;
    wire N__45210;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45192;
    wire N__45189;
    wire N__45186;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45107;
    wire N__45106;
    wire N__45105;
    wire N__45102;
    wire N__45101;
    wire N__45100;
    wire N__45099;
    wire N__45098;
    wire N__45095;
    wire N__45092;
    wire N__45091;
    wire N__45090;
    wire N__45089;
    wire N__45086;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45062;
    wire N__45059;
    wire N__45056;
    wire N__45053;
    wire N__45046;
    wire N__45037;
    wire N__45034;
    wire N__45021;
    wire N__45020;
    wire N__45019;
    wire N__45014;
    wire N__45011;
    wire N__45010;
    wire N__45007;
    wire N__45006;
    wire N__45003;
    wire N__45000;
    wire N__44997;
    wire N__44996;
    wire N__44995;
    wire N__44992;
    wire N__44991;
    wire N__44990;
    wire N__44985;
    wire N__44982;
    wire N__44981;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44969;
    wire N__44968;
    wire N__44965;
    wire N__44964;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44946;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44929;
    wire N__44926;
    wire N__44913;
    wire N__44912;
    wire N__44911;
    wire N__44910;
    wire N__44909;
    wire N__44908;
    wire N__44907;
    wire N__44904;
    wire N__44903;
    wire N__44902;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44892;
    wire N__44891;
    wire N__44890;
    wire N__44887;
    wire N__44886;
    wire N__44883;
    wire N__44880;
    wire N__44879;
    wire N__44878;
    wire N__44875;
    wire N__44874;
    wire N__44873;
    wire N__44872;
    wire N__44871;
    wire N__44868;
    wire N__44863;
    wire N__44860;
    wire N__44855;
    wire N__44854;
    wire N__44853;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44837;
    wire N__44832;
    wire N__44831;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44819;
    wire N__44816;
    wire N__44807;
    wire N__44802;
    wire N__44799;
    wire N__44790;
    wire N__44787;
    wire N__44784;
    wire N__44777;
    wire N__44770;
    wire N__44765;
    wire N__44754;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44739;
    wire N__44738;
    wire N__44737;
    wire N__44734;
    wire N__44729;
    wire N__44724;
    wire N__44721;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44708;
    wire N__44705;
    wire N__44702;
    wire N__44699;
    wire N__44698;
    wire N__44695;
    wire N__44692;
    wire N__44689;
    wire N__44686;
    wire N__44679;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44643;
    wire N__44642;
    wire N__44639;
    wire N__44636;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44619;
    wire N__44616;
    wire N__44615;
    wire N__44612;
    wire N__44609;
    wire N__44608;
    wire N__44605;
    wire N__44600;
    wire N__44595;
    wire N__44592;
    wire N__44589;
    wire N__44586;
    wire N__44585;
    wire N__44582;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44569;
    wire N__44562;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44544;
    wire N__44541;
    wire N__44540;
    wire N__44539;
    wire N__44538;
    wire N__44537;
    wire N__44536;
    wire N__44535;
    wire N__44534;
    wire N__44533;
    wire N__44532;
    wire N__44531;
    wire N__44530;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44509;
    wire N__44504;
    wire N__44503;
    wire N__44500;
    wire N__44497;
    wire N__44494;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44474;
    wire N__44471;
    wire N__44468;
    wire N__44463;
    wire N__44460;
    wire N__44453;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44435;
    wire N__44432;
    wire N__44431;
    wire N__44430;
    wire N__44427;
    wire N__44426;
    wire N__44423;
    wire N__44422;
    wire N__44421;
    wire N__44418;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44405;
    wire N__44402;
    wire N__44399;
    wire N__44396;
    wire N__44393;
    wire N__44390;
    wire N__44389;
    wire N__44388;
    wire N__44387;
    wire N__44384;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44355;
    wire N__44350;
    wire N__44339;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44310;
    wire N__44309;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44282;
    wire N__44279;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44269;
    wire N__44266;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44231;
    wire N__44228;
    wire N__44225;
    wire N__44220;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44204;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44184;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44168;
    wire N__44165;
    wire N__44162;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44114;
    wire N__44113;
    wire N__44112;
    wire N__44111;
    wire N__44108;
    wire N__44107;
    wire N__44106;
    wire N__44105;
    wire N__44102;
    wire N__44099;
    wire N__44096;
    wire N__44095;
    wire N__44092;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44076;
    wire N__44073;
    wire N__44070;
    wire N__44067;
    wire N__44064;
    wire N__44063;
    wire N__44060;
    wire N__44055;
    wire N__44052;
    wire N__44047;
    wire N__44044;
    wire N__44041;
    wire N__44036;
    wire N__44033;
    wire N__44028;
    wire N__44021;
    wire N__44016;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43989;
    wire N__43988;
    wire N__43985;
    wire N__43982;
    wire N__43977;
    wire N__43976;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43955;
    wire N__43952;
    wire N__43951;
    wire N__43948;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43940;
    wire N__43939;
    wire N__43936;
    wire N__43933;
    wire N__43932;
    wire N__43929;
    wire N__43926;
    wire N__43925;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43913;
    wire N__43912;
    wire N__43911;
    wire N__43910;
    wire N__43907;
    wire N__43902;
    wire N__43899;
    wire N__43898;
    wire N__43897;
    wire N__43896;
    wire N__43895;
    wire N__43894;
    wire N__43893;
    wire N__43892;
    wire N__43891;
    wire N__43890;
    wire N__43887;
    wire N__43884;
    wire N__43879;
    wire N__43876;
    wire N__43875;
    wire N__43874;
    wire N__43869;
    wire N__43866;
    wire N__43861;
    wire N__43858;
    wire N__43853;
    wire N__43846;
    wire N__43843;
    wire N__43840;
    wire N__43837;
    wire N__43836;
    wire N__43833;
    wire N__43828;
    wire N__43825;
    wire N__43824;
    wire N__43823;
    wire N__43822;
    wire N__43819;
    wire N__43818;
    wire N__43817;
    wire N__43814;
    wire N__43811;
    wire N__43806;
    wire N__43797;
    wire N__43794;
    wire N__43791;
    wire N__43788;
    wire N__43783;
    wire N__43780;
    wire N__43777;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43765;
    wire N__43762;
    wire N__43755;
    wire N__43752;
    wire N__43745;
    wire N__43740;
    wire N__43737;
    wire N__43716;
    wire N__43715;
    wire N__43712;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43701;
    wire N__43698;
    wire N__43693;
    wire N__43692;
    wire N__43691;
    wire N__43688;
    wire N__43685;
    wire N__43682;
    wire N__43681;
    wire N__43680;
    wire N__43677;
    wire N__43676;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43668;
    wire N__43663;
    wire N__43660;
    wire N__43653;
    wire N__43652;
    wire N__43651;
    wire N__43648;
    wire N__43645;
    wire N__43642;
    wire N__43641;
    wire N__43640;
    wire N__43637;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43614;
    wire N__43611;
    wire N__43606;
    wire N__43601;
    wire N__43600;
    wire N__43597;
    wire N__43596;
    wire N__43593;
    wire N__43592;
    wire N__43589;
    wire N__43588;
    wire N__43585;
    wire N__43584;
    wire N__43581;
    wire N__43576;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43541;
    wire N__43536;
    wire N__43533;
    wire N__43528;
    wire N__43521;
    wire N__43506;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43492;
    wire N__43491;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43473;
    wire N__43470;
    wire N__43467;
    wire N__43464;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43449;
    wire N__43446;
    wire N__43443;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43431;
    wire N__43430;
    wire N__43429;
    wire N__43428;
    wire N__43425;
    wire N__43424;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43399;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43381;
    wire N__43378;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43340;
    wire N__43337;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43308;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43272;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43245;
    wire N__43244;
    wire N__43243;
    wire N__43242;
    wire N__43241;
    wire N__43240;
    wire N__43239;
    wire N__43238;
    wire N__43237;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43225;
    wire N__43218;
    wire N__43211;
    wire N__43200;
    wire N__43197;
    wire N__43194;
    wire N__43191;
    wire N__43190;
    wire N__43187;
    wire N__43186;
    wire N__43185;
    wire N__43184;
    wire N__43183;
    wire N__43180;
    wire N__43175;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43148;
    wire N__43143;
    wire N__43140;
    wire N__43137;
    wire N__43128;
    wire N__43125;
    wire N__43122;
    wire N__43119;
    wire N__43116;
    wire N__43115;
    wire N__43112;
    wire N__43109;
    wire N__43104;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43092;
    wire N__43091;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43074;
    wire N__43073;
    wire N__43070;
    wire N__43067;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43043;
    wire N__43042;
    wire N__43039;
    wire N__43034;
    wire N__43029;
    wire N__43026;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43010;
    wire N__43009;
    wire N__43006;
    wire N__43001;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42977;
    wire N__42974;
    wire N__42971;
    wire N__42966;
    wire N__42963;
    wire N__42960;
    wire N__42957;
    wire N__42954;
    wire N__42951;
    wire N__42950;
    wire N__42947;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42908;
    wire N__42907;
    wire N__42904;
    wire N__42899;
    wire N__42894;
    wire N__42891;
    wire N__42888;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42880;
    wire N__42879;
    wire N__42878;
    wire N__42877;
    wire N__42876;
    wire N__42875;
    wire N__42874;
    wire N__42869;
    wire N__42862;
    wire N__42853;
    wire N__42850;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42831;
    wire N__42828;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42807;
    wire N__42804;
    wire N__42801;
    wire N__42798;
    wire N__42797;
    wire N__42794;
    wire N__42791;
    wire N__42786;
    wire N__42785;
    wire N__42782;
    wire N__42779;
    wire N__42776;
    wire N__42771;
    wire N__42768;
    wire N__42767;
    wire N__42764;
    wire N__42761;
    wire N__42756;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42744;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42732;
    wire N__42729;
    wire N__42728;
    wire N__42725;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42715;
    wire N__42712;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42698;
    wire N__42695;
    wire N__42694;
    wire N__42691;
    wire N__42688;
    wire N__42685;
    wire N__42682;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42639;
    wire N__42636;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42628;
    wire N__42627;
    wire N__42622;
    wire N__42619;
    wire N__42616;
    wire N__42615;
    wire N__42614;
    wire N__42613;
    wire N__42610;
    wire N__42605;
    wire N__42604;
    wire N__42603;
    wire N__42600;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42588;
    wire N__42587;
    wire N__42584;
    wire N__42583;
    wire N__42582;
    wire N__42579;
    wire N__42578;
    wire N__42575;
    wire N__42572;
    wire N__42569;
    wire N__42566;
    wire N__42561;
    wire N__42558;
    wire N__42553;
    wire N__42550;
    wire N__42547;
    wire N__42542;
    wire N__42539;
    wire N__42536;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42509;
    wire N__42506;
    wire N__42503;
    wire N__42498;
    wire N__42495;
    wire N__42494;
    wire N__42491;
    wire N__42488;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42476;
    wire N__42473;
    wire N__42470;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42435;
    wire N__42434;
    wire N__42433;
    wire N__42432;
    wire N__42431;
    wire N__42428;
    wire N__42427;
    wire N__42424;
    wire N__42423;
    wire N__42420;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42398;
    wire N__42395;
    wire N__42392;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42362;
    wire N__42359;
    wire N__42356;
    wire N__42353;
    wire N__42350;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42332;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42312;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42300;
    wire N__42299;
    wire N__42298;
    wire N__42297;
    wire N__42296;
    wire N__42295;
    wire N__42294;
    wire N__42293;
    wire N__42290;
    wire N__42289;
    wire N__42288;
    wire N__42287;
    wire N__42284;
    wire N__42283;
    wire N__42282;
    wire N__42281;
    wire N__42280;
    wire N__42279;
    wire N__42276;
    wire N__42275;
    wire N__42274;
    wire N__42271;
    wire N__42270;
    wire N__42269;
    wire N__42268;
    wire N__42267;
    wire N__42264;
    wire N__42263;
    wire N__42262;
    wire N__42259;
    wire N__42258;
    wire N__42257;
    wire N__42256;
    wire N__42255;
    wire N__42254;
    wire N__42253;
    wire N__42252;
    wire N__42251;
    wire N__42244;
    wire N__42239;
    wire N__42230;
    wire N__42229;
    wire N__42226;
    wire N__42225;
    wire N__42224;
    wire N__42223;
    wire N__42222;
    wire N__42221;
    wire N__42220;
    wire N__42219;
    wire N__42218;
    wire N__42217;
    wire N__42216;
    wire N__42215;
    wire N__42214;
    wire N__42213;
    wire N__42212;
    wire N__42211;
    wire N__42210;
    wire N__42209;
    wire N__42208;
    wire N__42207;
    wire N__42206;
    wire N__42205;
    wire N__42204;
    wire N__42203;
    wire N__42202;
    wire N__42201;
    wire N__42200;
    wire N__42199;
    wire N__42198;
    wire N__42197;
    wire N__42196;
    wire N__42195;
    wire N__42194;
    wire N__42193;
    wire N__42188;
    wire N__42187;
    wire N__42176;
    wire N__42175;
    wire N__42174;
    wire N__42173;
    wire N__42172;
    wire N__42171;
    wire N__42170;
    wire N__42169;
    wire N__42168;
    wire N__42163;
    wire N__42154;
    wire N__42145;
    wire N__42142;
    wire N__42141;
    wire N__42140;
    wire N__42139;
    wire N__42138;
    wire N__42129;
    wire N__42128;
    wire N__42127;
    wire N__42126;
    wire N__42125;
    wire N__42124;
    wire N__42123;
    wire N__42122;
    wire N__42121;
    wire N__42120;
    wire N__42113;
    wire N__42110;
    wire N__42105;
    wire N__42102;
    wire N__42099;
    wire N__42098;
    wire N__42097;
    wire N__42096;
    wire N__42095;
    wire N__42094;
    wire N__42093;
    wire N__42092;
    wire N__42091;
    wire N__42090;
    wire N__42089;
    wire N__42088;
    wire N__42087;
    wire N__42086;
    wire N__42077;
    wire N__42072;
    wire N__42071;
    wire N__42068;
    wire N__42067;
    wire N__42066;
    wire N__42065;
    wire N__42064;
    wire N__42063;
    wire N__42062;
    wire N__42061;
    wire N__42060;
    wire N__42059;
    wire N__42058;
    wire N__42057;
    wire N__42056;
    wire N__42055;
    wire N__42054;
    wire N__42053;
    wire N__42052;
    wire N__42051;
    wire N__42050;
    wire N__42049;
    wire N__42048;
    wire N__42047;
    wire N__42044;
    wire N__42043;
    wire N__42042;
    wire N__42041;
    wire N__42034;
    wire N__42033;
    wire N__42032;
    wire N__42031;
    wire N__42030;
    wire N__42027;
    wire N__42026;
    wire N__42025;
    wire N__42024;
    wire N__42023;
    wire N__42022;
    wire N__42021;
    wire N__42020;
    wire N__42019;
    wire N__42016;
    wire N__42015;
    wire N__42014;
    wire N__42013;
    wire N__42012;
    wire N__42011;
    wire N__42010;
    wire N__42009;
    wire N__42006;
    wire N__42005;
    wire N__42004;
    wire N__42003;
    wire N__42002;
    wire N__42001;
    wire N__42000;
    wire N__41999;
    wire N__41998;
    wire N__41997;
    wire N__41988;
    wire N__41979;
    wire N__41978;
    wire N__41977;
    wire N__41976;
    wire N__41975;
    wire N__41974;
    wire N__41969;
    wire N__41968;
    wire N__41967;
    wire N__41966;
    wire N__41965;
    wire N__41964;
    wire N__41963;
    wire N__41960;
    wire N__41953;
    wire N__41948;
    wire N__41945;
    wire N__41944;
    wire N__41943;
    wire N__41940;
    wire N__41939;
    wire N__41938;
    wire N__41937;
    wire N__41936;
    wire N__41935;
    wire N__41932;
    wire N__41923;
    wire N__41914;
    wire N__41905;
    wire N__41896;
    wire N__41893;
    wire N__41886;
    wire N__41879;
    wire N__41876;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41868;
    wire N__41867;
    wire N__41866;
    wire N__41865;
    wire N__41864;
    wire N__41863;
    wire N__41862;
    wire N__41855;
    wire N__41850;
    wire N__41843;
    wire N__41836;
    wire N__41827;
    wire N__41820;
    wire N__41815;
    wire N__41814;
    wire N__41813;
    wire N__41812;
    wire N__41811;
    wire N__41810;
    wire N__41807;
    wire N__41806;
    wire N__41805;
    wire N__41802;
    wire N__41793;
    wire N__41786;
    wire N__41783;
    wire N__41772;
    wire N__41763;
    wire N__41754;
    wire N__41753;
    wire N__41752;
    wire N__41751;
    wire N__41750;
    wire N__41749;
    wire N__41748;
    wire N__41747;
    wire N__41746;
    wire N__41745;
    wire N__41744;
    wire N__41743;
    wire N__41742;
    wire N__41739;
    wire N__41732;
    wire N__41729;
    wire N__41724;
    wire N__41713;
    wire N__41704;
    wire N__41695;
    wire N__41688;
    wire N__41681;
    wire N__41680;
    wire N__41679;
    wire N__41672;
    wire N__41663;
    wire N__41658;
    wire N__41657;
    wire N__41656;
    wire N__41655;
    wire N__41654;
    wire N__41653;
    wire N__41652;
    wire N__41649;
    wire N__41648;
    wire N__41647;
    wire N__41646;
    wire N__41645;
    wire N__41644;
    wire N__41643;
    wire N__41642;
    wire N__41641;
    wire N__41640;
    wire N__41639;
    wire N__41638;
    wire N__41633;
    wire N__41632;
    wire N__41631;
    wire N__41630;
    wire N__41629;
    wire N__41628;
    wire N__41627;
    wire N__41620;
    wire N__41619;
    wire N__41618;
    wire N__41617;
    wire N__41616;
    wire N__41615;
    wire N__41614;
    wire N__41613;
    wire N__41612;
    wire N__41611;
    wire N__41610;
    wire N__41609;
    wire N__41608;
    wire N__41607;
    wire N__41606;
    wire N__41605;
    wire N__41604;
    wire N__41601;
    wire N__41600;
    wire N__41599;
    wire N__41598;
    wire N__41597;
    wire N__41596;
    wire N__41593;
    wire N__41592;
    wire N__41591;
    wire N__41590;
    wire N__41589;
    wire N__41586;
    wire N__41579;
    wire N__41578;
    wire N__41577;
    wire N__41574;
    wire N__41573;
    wire N__41572;
    wire N__41569;
    wire N__41568;
    wire N__41567;
    wire N__41566;
    wire N__41565;
    wire N__41562;
    wire N__41561;
    wire N__41560;
    wire N__41559;
    wire N__41552;
    wire N__41549;
    wire N__41540;
    wire N__41531;
    wire N__41524;
    wire N__41519;
    wire N__41512;
    wire N__41509;
    wire N__41502;
    wire N__41499;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41483;
    wire N__41480;
    wire N__41479;
    wire N__41478;
    wire N__41477;
    wire N__41476;
    wire N__41475;
    wire N__41474;
    wire N__41473;
    wire N__41472;
    wire N__41467;
    wire N__41462;
    wire N__41457;
    wire N__41454;
    wire N__41445;
    wire N__41436;
    wire N__41421;
    wire N__41414;
    wire N__41407;
    wire N__41400;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41372;
    wire N__41367;
    wire N__41360;
    wire N__41353;
    wire N__41342;
    wire N__41333;
    wire N__41324;
    wire N__41323;
    wire N__41322;
    wire N__41321;
    wire N__41318;
    wire N__41317;
    wire N__41316;
    wire N__41315;
    wire N__41314;
    wire N__41311;
    wire N__41310;
    wire N__41309;
    wire N__41308;
    wire N__41305;
    wire N__41298;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41278;
    wire N__41271;
    wire N__41264;
    wire N__41259;
    wire N__41252;
    wire N__41241;
    wire N__41232;
    wire N__41227;
    wire N__41224;
    wire N__41219;
    wire N__41210;
    wire N__41201;
    wire N__41192;
    wire N__41187;
    wire N__41184;
    wire N__41177;
    wire N__41174;
    wire N__41169;
    wire N__41164;
    wire N__41157;
    wire N__41146;
    wire N__41137;
    wire N__41128;
    wire N__41123;
    wire N__41116;
    wire N__41103;
    wire N__41094;
    wire N__41083;
    wire N__41078;
    wire N__41069;
    wire N__41064;
    wire N__41055;
    wire N__41042;
    wire N__41037;
    wire N__41014;
    wire N__41009;
    wire N__40994;
    wire N__40987;
    wire N__40974;
    wire N__40971;
    wire N__40966;
    wire N__40961;
    wire N__40956;
    wire N__40947;
    wire N__40946;
    wire N__40943;
    wire N__40940;
    wire N__40937;
    wire N__40934;
    wire N__40929;
    wire N__40928;
    wire N__40927;
    wire N__40926;
    wire N__40923;
    wire N__40922;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40914;
    wire N__40911;
    wire N__40908;
    wire N__40907;
    wire N__40904;
    wire N__40903;
    wire N__40902;
    wire N__40901;
    wire N__40900;
    wire N__40899;
    wire N__40898;
    wire N__40895;
    wire N__40894;
    wire N__40891;
    wire N__40886;
    wire N__40881;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40864;
    wire N__40863;
    wire N__40862;
    wire N__40861;
    wire N__40860;
    wire N__40859;
    wire N__40856;
    wire N__40849;
    wire N__40840;
    wire N__40835;
    wire N__40828;
    wire N__40819;
    wire N__40806;
    wire N__40803;
    wire N__40802;
    wire N__40799;
    wire N__40796;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40784;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40769;
    wire N__40766;
    wire N__40763;
    wire N__40758;
    wire N__40755;
    wire N__40752;
    wire N__40749;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40736;
    wire N__40733;
    wire N__40730;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40707;
    wire N__40704;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40692;
    wire N__40691;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40662;
    wire N__40659;
    wire N__40658;
    wire N__40655;
    wire N__40652;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40637;
    wire N__40634;
    wire N__40631;
    wire N__40628;
    wire N__40623;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40604;
    wire N__40601;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40584;
    wire N__40581;
    wire N__40578;
    wire N__40575;
    wire N__40572;
    wire N__40569;
    wire N__40566;
    wire N__40565;
    wire N__40562;
    wire N__40559;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40542;
    wire N__40539;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40523;
    wire N__40520;
    wire N__40517;
    wire N__40516;
    wire N__40513;
    wire N__40510;
    wire N__40507;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40475;
    wire N__40474;
    wire N__40471;
    wire N__40466;
    wire N__40463;
    wire N__40458;
    wire N__40455;
    wire N__40452;
    wire N__40449;
    wire N__40446;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40428;
    wire N__40425;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40408;
    wire N__40405;
    wire N__40402;
    wire N__40399;
    wire N__40396;
    wire N__40389;
    wire N__40386;
    wire N__40383;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40373;
    wire N__40372;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40360;
    wire N__40357;
    wire N__40354;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40322;
    wire N__40321;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40309;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40241;
    wire N__40238;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40228;
    wire N__40221;
    wire N__40218;
    wire N__40215;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40202;
    wire N__40201;
    wire N__40198;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40181;
    wire N__40176;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40163;
    wire N__40160;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40137;
    wire N__40134;
    wire N__40131;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40106;
    wire N__40105;
    wire N__40102;
    wire N__40101;
    wire N__40100;
    wire N__40099;
    wire N__40098;
    wire N__40097;
    wire N__40096;
    wire N__40095;
    wire N__40094;
    wire N__40093;
    wire N__40092;
    wire N__40091;
    wire N__40088;
    wire N__40085;
    wire N__40080;
    wire N__40079;
    wire N__40078;
    wire N__40077;
    wire N__40076;
    wire N__40065;
    wire N__40062;
    wire N__40059;
    wire N__40058;
    wire N__40055;
    wire N__40052;
    wire N__40051;
    wire N__40048;
    wire N__40047;
    wire N__40046;
    wire N__40039;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40023;
    wire N__40012;
    wire N__40005;
    wire N__40002;
    wire N__39987;
    wire N__39984;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39965;
    wire N__39962;
    wire N__39959;
    wire N__39956;
    wire N__39951;
    wire N__39950;
    wire N__39949;
    wire N__39944;
    wire N__39941;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39927;
    wire N__39924;
    wire N__39923;
    wire N__39922;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39899;
    wire N__39896;
    wire N__39893;
    wire N__39890;
    wire N__39887;
    wire N__39884;
    wire N__39881;
    wire N__39878;
    wire N__39873;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39855;
    wire N__39852;
    wire N__39849;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39839;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39824;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39806;
    wire N__39805;
    wire N__39802;
    wire N__39797;
    wire N__39794;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39770;
    wire N__39767;
    wire N__39764;
    wire N__39761;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39747;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39731;
    wire N__39728;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39710;
    wire N__39705;
    wire N__39702;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39669;
    wire N__39666;
    wire N__39663;
    wire N__39660;
    wire N__39657;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39644;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39603;
    wire N__39600;
    wire N__39599;
    wire N__39596;
    wire N__39593;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39545;
    wire N__39542;
    wire N__39539;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39522;
    wire N__39519;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39487;
    wire N__39484;
    wire N__39481;
    wire N__39478;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39453;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39391;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39359;
    wire N__39356;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39339;
    wire N__39338;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39306;
    wire N__39305;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39289;
    wire N__39284;
    wire N__39281;
    wire N__39278;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39173;
    wire N__39170;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39125;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39087;
    wire N__39086;
    wire N__39083;
    wire N__39080;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39062;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39020;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38978;
    wire N__38977;
    wire N__38974;
    wire N__38969;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38942;
    wire N__38939;
    wire N__38936;
    wire N__38931;
    wire N__38928;
    wire N__38927;
    wire N__38924;
    wire N__38921;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38913;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38890;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38861;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38825;
    wire N__38822;
    wire N__38821;
    wire N__38818;
    wire N__38815;
    wire N__38812;
    wire N__38809;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38773;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38724;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38711;
    wire N__38708;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38695;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38672;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38592;
    wire N__38591;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38574;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38531;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38519;
    wire N__38518;
    wire N__38513;
    wire N__38510;
    wire N__38505;
    wire N__38504;
    wire N__38503;
    wire N__38502;
    wire N__38501;
    wire N__38500;
    wire N__38499;
    wire N__38498;
    wire N__38497;
    wire N__38496;
    wire N__38493;
    wire N__38492;
    wire N__38489;
    wire N__38488;
    wire N__38487;
    wire N__38482;
    wire N__38479;
    wire N__38478;
    wire N__38475;
    wire N__38474;
    wire N__38471;
    wire N__38470;
    wire N__38469;
    wire N__38466;
    wire N__38465;
    wire N__38462;
    wire N__38461;
    wire N__38460;
    wire N__38457;
    wire N__38456;
    wire N__38445;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38431;
    wire N__38424;
    wire N__38419;
    wire N__38408;
    wire N__38391;
    wire N__38390;
    wire N__38387;
    wire N__38384;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38334;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38321;
    wire N__38318;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38298;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38290;
    wire N__38287;
    wire N__38284;
    wire N__38281;
    wire N__38278;
    wire N__38273;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38259;
    wire N__38258;
    wire N__38255;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38208;
    wire N__38205;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38187;
    wire N__38184;
    wire N__38181;
    wire N__38180;
    wire N__38177;
    wire N__38174;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38147;
    wire N__38144;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38105;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38022;
    wire N__38021;
    wire N__38018;
    wire N__38017;
    wire N__38016;
    wire N__38015;
    wire N__38014;
    wire N__38013;
    wire N__38012;
    wire N__38011;
    wire N__38010;
    wire N__38009;
    wire N__38008;
    wire N__38005;
    wire N__38004;
    wire N__38001;
    wire N__38000;
    wire N__37999;
    wire N__37996;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37988;
    wire N__37987;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37968;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37958;
    wire N__37949;
    wire N__37944;
    wire N__37939;
    wire N__37936;
    wire N__37925;
    wire N__37920;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37898;
    wire N__37897;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37879;
    wire N__37876;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37857;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37821;
    wire N__37818;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37805;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37766;
    wire N__37763;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37743;
    wire N__37740;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37718;
    wire N__37715;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37702;
    wire N__37695;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37674;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37662;
    wire N__37659;
    wire N__37658;
    wire N__37655;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37607;
    wire N__37606;
    wire N__37605;
    wire N__37604;
    wire N__37603;
    wire N__37602;
    wire N__37599;
    wire N__37598;
    wire N__37597;
    wire N__37596;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37588;
    wire N__37581;
    wire N__37580;
    wire N__37579;
    wire N__37576;
    wire N__37575;
    wire N__37570;
    wire N__37567;
    wire N__37566;
    wire N__37565;
    wire N__37564;
    wire N__37561;
    wire N__37560;
    wire N__37557;
    wire N__37556;
    wire N__37555;
    wire N__37552;
    wire N__37547;
    wire N__37544;
    wire N__37539;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37521;
    wire N__37518;
    wire N__37517;
    wire N__37514;
    wire N__37513;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37493;
    wire N__37486;
    wire N__37479;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37449;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37437;
    wire N__37436;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37422;
    wire N__37419;
    wire N__37418;
    wire N__37417;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37405;
    wire N__37402;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37383;
    wire N__37382;
    wire N__37381;
    wire N__37378;
    wire N__37375;
    wire N__37372;
    wire N__37367;
    wire N__37364;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37323;
    wire N__37322;
    wire N__37321;
    wire N__37320;
    wire N__37319;
    wire N__37318;
    wire N__37317;
    wire N__37314;
    wire N__37313;
    wire N__37312;
    wire N__37311;
    wire N__37308;
    wire N__37307;
    wire N__37306;
    wire N__37305;
    wire N__37304;
    wire N__37303;
    wire N__37300;
    wire N__37299;
    wire N__37298;
    wire N__37295;
    wire N__37294;
    wire N__37293;
    wire N__37288;
    wire N__37285;
    wire N__37280;
    wire N__37277;
    wire N__37276;
    wire N__37269;
    wire N__37264;
    wire N__37263;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37255;
    wire N__37252;
    wire N__37241;
    wire N__37232;
    wire N__37231;
    wire N__37228;
    wire N__37227;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37208;
    wire N__37201;
    wire N__37194;
    wire N__37189;
    wire N__37186;
    wire N__37173;
    wire N__37170;
    wire N__37167;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37159;
    wire N__37154;
    wire N__37151;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37104;
    wire N__37103;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37044;
    wire N__37041;
    wire N__37038;
    wire N__37035;
    wire N__37032;
    wire N__37029;
    wire N__37026;
    wire N__37023;
    wire N__37020;
    wire N__37017;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36948;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36936;
    wire N__36933;
    wire N__36930;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36912;
    wire N__36911;
    wire N__36908;
    wire N__36905;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36878;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36857;
    wire N__36854;
    wire N__36849;
    wire N__36846;
    wire N__36845;
    wire N__36842;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36822;
    wire N__36819;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36803;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36777;
    wire N__36774;
    wire N__36771;
    wire N__36768;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36690;
    wire N__36689;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36672;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36655;
    wire N__36648;
    wire N__36645;
    wire N__36642;
    wire N__36639;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36631;
    wire N__36628;
    wire N__36625;
    wire N__36622;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36600;
    wire N__36597;
    wire N__36594;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36564;
    wire N__36563;
    wire N__36562;
    wire N__36561;
    wire N__36560;
    wire N__36559;
    wire N__36558;
    wire N__36557;
    wire N__36554;
    wire N__36553;
    wire N__36552;
    wire N__36549;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36538;
    wire N__36535;
    wire N__36534;
    wire N__36533;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36525;
    wire N__36524;
    wire N__36519;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36501;
    wire N__36496;
    wire N__36491;
    wire N__36482;
    wire N__36475;
    wire N__36472;
    wire N__36459;
    wire N__36456;
    wire N__36455;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36442;
    wire N__36439;
    wire N__36436;
    wire N__36433;
    wire N__36430;
    wire N__36423;
    wire N__36422;
    wire N__36419;
    wire N__36416;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36401;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36387;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36333;
    wire N__36330;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36318;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36307;
    wire N__36302;
    wire N__36299;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36229;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36203;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36186;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36147;
    wire N__36144;
    wire N__36141;
    wire N__36138;
    wire N__36135;
    wire N__36132;
    wire N__36131;
    wire N__36128;
    wire N__36127;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36106;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36060;
    wire N__36059;
    wire N__36058;
    wire N__36057;
    wire N__36054;
    wire N__36049;
    wire N__36046;
    wire N__36045;
    wire N__36042;
    wire N__36039;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35995;
    wire N__35992;
    wire N__35989;
    wire N__35986;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35969;
    wire N__35968;
    wire N__35965;
    wire N__35962;
    wire N__35957;
    wire N__35954;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35850;
    wire N__35847;
    wire N__35844;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35836;
    wire N__35831;
    wire N__35828;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35805;
    wire N__35804;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35764;
    wire N__35761;
    wire N__35758;
    wire N__35755;
    wire N__35752;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35733;
    wire N__35730;
    wire N__35727;
    wire N__35724;
    wire N__35721;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35709;
    wire N__35706;
    wire N__35703;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35688;
    wire N__35685;
    wire N__35682;
    wire N__35679;
    wire N__35676;
    wire N__35673;
    wire N__35670;
    wire N__35667;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35622;
    wire N__35619;
    wire N__35616;
    wire N__35613;
    wire N__35612;
    wire N__35611;
    wire N__35608;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35596;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35577;
    wire N__35574;
    wire N__35571;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35560;
    wire N__35555;
    wire N__35552;
    wire N__35547;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35535;
    wire N__35532;
    wire N__35529;
    wire N__35528;
    wire N__35525;
    wire N__35522;
    wire N__35517;
    wire N__35516;
    wire N__35515;
    wire N__35512;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35486;
    wire N__35481;
    wire N__35478;
    wire N__35475;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35412;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35382;
    wire N__35379;
    wire N__35376;
    wire N__35373;
    wire N__35370;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35334;
    wire N__35331;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35316;
    wire N__35313;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35301;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35283;
    wire N__35282;
    wire N__35279;
    wire N__35276;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35258;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35234;
    wire N__35233;
    wire N__35232;
    wire N__35229;
    wire N__35226;
    wire N__35223;
    wire N__35220;
    wire N__35217;
    wire N__35214;
    wire N__35205;
    wire N__35202;
    wire N__35199;
    wire N__35196;
    wire N__35193;
    wire N__35190;
    wire N__35187;
    wire N__35186;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35150;
    wire N__35147;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35105;
    wire N__35100;
    wire N__35099;
    wire N__35096;
    wire N__35093;
    wire N__35090;
    wire N__35087;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35069;
    wire N__35066;
    wire N__35065;
    wire N__35062;
    wire N__35059;
    wire N__35056;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35040;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35027;
    wire N__35026;
    wire N__35021;
    wire N__35018;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34962;
    wire N__34959;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34947;
    wire N__34944;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34936;
    wire N__34931;
    wire N__34928;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34907;
    wire N__34904;
    wire N__34901;
    wire N__34896;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34884;
    wire N__34883;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34859;
    wire N__34856;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34805;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34790;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34717;
    wire N__34714;
    wire N__34711;
    wire N__34708;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34679;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34656;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34643;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34601;
    wire N__34600;
    wire N__34597;
    wire N__34592;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34571;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34499;
    wire N__34498;
    wire N__34495;
    wire N__34492;
    wire N__34489;
    wire N__34486;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34469;
    wire N__34466;
    wire N__34463;
    wire N__34460;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34443;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34344;
    wire N__34341;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34333;
    wire N__34330;
    wire N__34329;
    wire N__34328;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34313;
    wire N__34310;
    wire N__34303;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34266;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34254;
    wire N__34251;
    wire N__34250;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34176;
    wire N__34173;
    wire N__34172;
    wire N__34169;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34127;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34079;
    wire N__34078;
    wire N__34075;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34055;
    wire N__34052;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34028;
    wire N__34027;
    wire N__34026;
    wire N__34025;
    wire N__34024;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34007;
    wire N__34006;
    wire N__34005;
    wire N__34004;
    wire N__34003;
    wire N__34002;
    wire N__34001;
    wire N__33998;
    wire N__33995;
    wire N__33990;
    wire N__33989;
    wire N__33988;
    wire N__33987;
    wire N__33986;
    wire N__33985;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33977;
    wire N__33974;
    wire N__33973;
    wire N__33972;
    wire N__33969;
    wire N__33968;
    wire N__33967;
    wire N__33966;
    wire N__33963;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33955;
    wire N__33948;
    wire N__33943;
    wire N__33930;
    wire N__33915;
    wire N__33902;
    wire N__33891;
    wire N__33888;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33846;
    wire N__33845;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33779;
    wire N__33776;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33752;
    wire N__33749;
    wire N__33746;
    wire N__33745;
    wire N__33740;
    wire N__33737;
    wire N__33732;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33720;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33668;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33626;
    wire N__33623;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33581;
    wire N__33578;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33554;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33536;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33467;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33413;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33365;
    wire N__33362;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33352;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33329;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33311;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33248;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33209;
    wire N__33206;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33164;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33110;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33054;
    wire N__33051;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33043;
    wire N__33040;
    wire N__33035;
    wire N__33032;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33006;
    wire N__33005;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32948;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32924;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32875;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32861;
    wire N__32856;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32843;
    wire N__32840;
    wire N__32837;
    wire N__32834;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32798;
    wire N__32795;
    wire N__32794;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32768;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32740;
    wire N__32737;
    wire N__32732;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32708;
    wire N__32707;
    wire N__32704;
    wire N__32701;
    wire N__32698;
    wire N__32695;
    wire N__32692;
    wire N__32689;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32673;
    wire N__32670;
    wire N__32669;
    wire N__32666;
    wire N__32665;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32642;
    wire N__32639;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32580;
    wire N__32579;
    wire N__32578;
    wire N__32577;
    wire N__32576;
    wire N__32573;
    wire N__32572;
    wire N__32571;
    wire N__32570;
    wire N__32569;
    wire N__32566;
    wire N__32563;
    wire N__32562;
    wire N__32561;
    wire N__32560;
    wire N__32559;
    wire N__32558;
    wire N__32555;
    wire N__32554;
    wire N__32553;
    wire N__32552;
    wire N__32549;
    wire N__32542;
    wire N__32539;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32525;
    wire N__32518;
    wire N__32511;
    wire N__32506;
    wire N__32503;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32462;
    wire N__32459;
    wire N__32456;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32400;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32392;
    wire N__32391;
    wire N__32386;
    wire N__32383;
    wire N__32380;
    wire N__32377;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32354;
    wire N__32353;
    wire N__32350;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32332;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32304;
    wire N__32301;
    wire N__32298;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32281;
    wire N__32274;
    wire N__32271;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32223;
    wire N__32222;
    wire N__32221;
    wire N__32220;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32204;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32132;
    wire N__32129;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32119;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32092;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32073;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32012;
    wire N__32011;
    wire N__32008;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31962;
    wire N__31959;
    wire N__31956;
    wire N__31955;
    wire N__31952;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31904;
    wire N__31901;
    wire N__31898;
    wire N__31895;
    wire N__31892;
    wire N__31887;
    wire N__31884;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31874;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31814;
    wire N__31813;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31794;
    wire N__31791;
    wire N__31790;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31779;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31755;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31724;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31709;
    wire N__31704;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31687;
    wire N__31682;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31641;
    wire N__31638;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31611;
    wire N__31608;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31578;
    wire N__31575;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31558;
    wire N__31555;
    wire N__31552;
    wire N__31549;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31529;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31509;
    wire N__31506;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31479;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31443;
    wire N__31440;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31420;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31370;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31278;
    wire N__31277;
    wire N__31276;
    wire N__31275;
    wire N__31274;
    wire N__31271;
    wire N__31270;
    wire N__31269;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31261;
    wire N__31260;
    wire N__31259;
    wire N__31256;
    wire N__31255;
    wire N__31254;
    wire N__31253;
    wire N__31252;
    wire N__31249;
    wire N__31244;
    wire N__31231;
    wire N__31230;
    wire N__31227;
    wire N__31226;
    wire N__31223;
    wire N__31222;
    wire N__31221;
    wire N__31220;
    wire N__31217;
    wire N__31216;
    wire N__31213;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31205;
    wire N__31202;
    wire N__31199;
    wire N__31196;
    wire N__31189;
    wire N__31186;
    wire N__31181;
    wire N__31172;
    wire N__31163;
    wire N__31154;
    wire N__31143;
    wire N__31140;
    wire N__31139;
    wire N__31138;
    wire N__31135;
    wire N__31132;
    wire N__31129;
    wire N__31126;
    wire N__31123;
    wire N__31118;
    wire N__31113;
    wire N__31112;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31092;
    wire N__31091;
    wire N__31088;
    wire N__31085;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31067;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31050;
    wire N__31049;
    wire N__31048;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31013;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30920;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30854;
    wire N__30851;
    wire N__30848;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30833;
    wire N__30830;
    wire N__30827;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30815;
    wire N__30812;
    wire N__30811;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30792;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30771;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30712;
    wire N__30709;
    wire N__30706;
    wire N__30703;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30671;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30628;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30582;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30569;
    wire N__30566;
    wire N__30563;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30533;
    wire N__30532;
    wire N__30529;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30511;
    wire N__30510;
    wire N__30507;
    wire N__30502;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30408;
    wire N__30405;
    wire N__30402;
    wire N__30399;
    wire N__30398;
    wire N__30397;
    wire N__30392;
    wire N__30389;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30354;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30338;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30249;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30146;
    wire N__30143;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30132;
    wire N__30129;
    wire N__30124;
    wire N__30123;
    wire N__30120;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30101;
    wire N__30096;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30066;
    wire N__30063;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30039;
    wire N__30036;
    wire N__30035;
    wire N__30032;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30022;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29999;
    wire N__29996;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29942;
    wire N__29939;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29929;
    wire N__29922;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29907;
    wire N__29904;
    wire N__29901;
    wire N__29898;
    wire N__29895;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29798;
    wire N__29797;
    wire N__29794;
    wire N__29789;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29774;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29727;
    wire N__29724;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29702;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29691;
    wire N__29690;
    wire N__29689;
    wire N__29688;
    wire N__29687;
    wire N__29686;
    wire N__29685;
    wire N__29684;
    wire N__29683;
    wire N__29682;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29678;
    wire N__29677;
    wire N__29676;
    wire N__29675;
    wire N__29674;
    wire N__29673;
    wire N__29672;
    wire N__29671;
    wire N__29670;
    wire N__29669;
    wire N__29666;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29587;
    wire N__29578;
    wire N__29569;
    wire N__29560;
    wire N__29551;
    wire N__29544;
    wire N__29537;
    wire N__29534;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29497;
    wire N__29492;
    wire N__29489;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29477;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29467;
    wire N__29462;
    wire N__29459;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29338;
    wire N__29333;
    wire N__29330;
    wire N__29329;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29301;
    wire N__29298;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29276;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29249;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29232;
    wire N__29229;
    wire N__29228;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29204;
    wire N__29201;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29191;
    wire N__29188;
    wire N__29181;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29127;
    wire N__29126;
    wire N__29125;
    wire N__29124;
    wire N__29123;
    wire N__29122;
    wire N__29121;
    wire N__29120;
    wire N__29117;
    wire N__29116;
    wire N__29113;
    wire N__29112;
    wire N__29111;
    wire N__29108;
    wire N__29107;
    wire N__29106;
    wire N__29105;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29095;
    wire N__29094;
    wire N__29089;
    wire N__29084;
    wire N__29075;
    wire N__29068;
    wire N__29057;
    wire N__29048;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29021;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28965;
    wire N__28964;
    wire N__28961;
    wire N__28958;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28937;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28929;
    wire N__28926;
    wire N__28921;
    wire N__28918;
    wire N__28917;
    wire N__28914;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28869;
    wire N__28868;
    wire N__28867;
    wire N__28864;
    wire N__28859;
    wire N__28856;
    wire N__28851;
    wire N__28848;
    wire N__28847;
    wire N__28844;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28832;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28820;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28804;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28790;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28712;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28647;
    wire N__28644;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28553;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28523;
    wire N__28522;
    wire N__28519;
    wire N__28514;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28340;
    wire N__28337;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28319;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28218;
    wire N__28215;
    wire N__28214;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28206;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28180;
    wire N__28175;
    wire N__28172;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28113;
    wire N__28110;
    wire N__28109;
    wire N__28108;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28083;
    wire N__28082;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28031;
    wire N__28028;
    wire N__28027;
    wire N__28024;
    wire N__28019;
    wire N__28016;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27974;
    wire N__27971;
    wire N__27970;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27884;
    wire N__27879;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27867;
    wire N__27864;
    wire N__27863;
    wire N__27858;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27846;
    wire N__27843;
    wire N__27842;
    wire N__27839;
    wire N__27834;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27815;
    wire N__27810;
    wire N__27807;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27606;
    wire N__27605;
    wire N__27602;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27582;
    wire N__27581;
    wire N__27580;
    wire N__27577;
    wire N__27576;
    wire N__27573;
    wire N__27572;
    wire N__27569;
    wire N__27568;
    wire N__27567;
    wire N__27558;
    wire N__27553;
    wire N__27552;
    wire N__27551;
    wire N__27550;
    wire N__27547;
    wire N__27546;
    wire N__27545;
    wire N__27544;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27518;
    wire N__27515;
    wire N__27510;
    wire N__27505;
    wire N__27498;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27396;
    wire N__27393;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27356;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27275;
    wire N__27272;
    wire N__27271;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27131;
    wire N__27128;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27115;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27089;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27063;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27047;
    wire N__27046;
    wire N__27043;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26859;
    wire N__26856;
    wire N__26855;
    wire N__26854;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26831;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26804;
    wire N__26803;
    wire N__26802;
    wire N__26801;
    wire N__26800;
    wire N__26799;
    wire N__26798;
    wire N__26797;
    wire N__26796;
    wire N__26795;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26781;
    wire N__26778;
    wire N__26777;
    wire N__26772;
    wire N__26769;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26737;
    wire N__26732;
    wire N__26725;
    wire N__26720;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26654;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26606;
    wire N__26605;
    wire N__26600;
    wire N__26597;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26565;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26504;
    wire N__26501;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26478;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26468;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26432;
    wire N__26431;
    wire N__26428;
    wire N__26423;
    wire N__26418;
    wire N__26417;
    wire N__26416;
    wire N__26413;
    wire N__26408;
    wire N__26405;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26354;
    wire N__26353;
    wire N__26350;
    wire N__26349;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26334;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26309;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26293;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26277;
    wire N__26276;
    wire N__26275;
    wire N__26272;
    wire N__26267;
    wire N__26264;
    wire N__26259;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26249;
    wire N__26248;
    wire N__26245;
    wire N__26240;
    wire N__26237;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26209;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26187;
    wire N__26182;
    wire N__26175;
    wire N__26174;
    wire N__26171;
    wire N__26170;
    wire N__26167;
    wire N__26162;
    wire N__26161;
    wire N__26156;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26129;
    wire N__26128;
    wire N__26127;
    wire N__26126;
    wire N__26123;
    wire N__26114;
    wire N__26109;
    wire N__26106;
    wire N__26103;
    wire N__26100;
    wire N__26097;
    wire N__26094;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26074;
    wire N__26073;
    wire N__26070;
    wire N__26069;
    wire N__26068;
    wire N__26065;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26046;
    wire N__26041;
    wire N__26034;
    wire N__26033;
    wire N__26030;
    wire N__26029;
    wire N__26026;
    wire N__26025;
    wire N__26022;
    wire N__26017;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__26001;
    wire N__25996;
    wire N__25989;
    wire N__25986;
    wire N__25985;
    wire N__25984;
    wire N__25979;
    wire N__25978;
    wire N__25975;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25954;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25940;
    wire N__25939;
    wire N__25938;
    wire N__25935;
    wire N__25928;
    wire N__25927;
    wire N__25926;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25914;
    wire N__25911;
    wire N__25904;
    wire N__25899;
    wire N__25898;
    wire N__25897;
    wire N__25896;
    wire N__25895;
    wire N__25894;
    wire N__25893;
    wire N__25890;
    wire N__25885;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25857;
    wire N__25856;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25830;
    wire N__25829;
    wire N__25828;
    wire N__25827;
    wire N__25824;
    wire N__25819;
    wire N__25816;
    wire N__25809;
    wire N__25808;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25796;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25769;
    wire N__25766;
    wire N__25761;
    wire N__25758;
    wire N__25757;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25680;
    wire N__25677;
    wire N__25676;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25599;
    wire N__25596;
    wire N__25595;
    wire N__25594;
    wire N__25589;
    wire N__25586;
    wire N__25581;
    wire N__25580;
    wire N__25579;
    wire N__25576;
    wire N__25571;
    wire N__25568;
    wire N__25563;
    wire N__25562;
    wire N__25561;
    wire N__25560;
    wire N__25559;
    wire N__25554;
    wire N__25551;
    wire N__25546;
    wire N__25539;
    wire N__25536;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25524;
    wire N__25523;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25515;
    wire N__25514;
    wire N__25511;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25482;
    wire N__25481;
    wire N__25478;
    wire N__25477;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25463;
    wire N__25460;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25441;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25415;
    wire N__25412;
    wire N__25411;
    wire N__25408;
    wire N__25403;
    wire N__25400;
    wire N__25395;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25367;
    wire N__25366;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25358;
    wire N__25357;
    wire N__25352;
    wire N__25345;
    wire N__25342;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25328;
    wire N__25327;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25291;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25239;
    wire N__25238;
    wire N__25237;
    wire N__25236;
    wire N__25235;
    wire N__25234;
    wire N__25233;
    wire N__25232;
    wire N__25231;
    wire N__25230;
    wire N__25229;
    wire N__25228;
    wire N__25227;
    wire N__25226;
    wire N__25225;
    wire N__25224;
    wire N__25221;
    wire N__25220;
    wire N__25219;
    wire N__25218;
    wire N__25217;
    wire N__25216;
    wire N__25213;
    wire N__25208;
    wire N__25201;
    wire N__25194;
    wire N__25185;
    wire N__25180;
    wire N__25179;
    wire N__25178;
    wire N__25177;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25166;
    wire N__25165;
    wire N__25158;
    wire N__25157;
    wire N__25156;
    wire N__25155;
    wire N__25152;
    wire N__25143;
    wire N__25140;
    wire N__25131;
    wire N__25126;
    wire N__25123;
    wire N__25118;
    wire N__25117;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25095;
    wire N__25088;
    wire N__25083;
    wire N__25068;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25025;
    wire N__25024;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25010;
    wire N__25007;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24983;
    wire N__24980;
    wire N__24979;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24965;
    wire N__24962;
    wire N__24957;
    wire N__24956;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24945;
    wire N__24944;
    wire N__24943;
    wire N__24942;
    wire N__24941;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24920;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24908;
    wire N__24907;
    wire N__24904;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24884;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24764;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24696;
    wire N__24695;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24678;
    wire N__24675;
    wire N__24674;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24640;
    wire N__24635;
    wire N__24632;
    wire N__24627;
    wire N__24626;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24606;
    wire N__24603;
    wire N__24602;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24582;
    wire N__24581;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24561;
    wire N__24560;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24543;
    wire N__24540;
    wire N__24539;
    wire N__24538;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24515;
    wire N__24514;
    wire N__24513;
    wire N__24512;
    wire N__24511;
    wire N__24510;
    wire N__24509;
    wire N__24508;
    wire N__24507;
    wire N__24506;
    wire N__24505;
    wire N__24504;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24458;
    wire N__24451;
    wire N__24450;
    wire N__24443;
    wire N__24434;
    wire N__24429;
    wire N__24426;
    wire N__24417;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24372;
    wire N__24371;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24344;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24324;
    wire N__24321;
    wire N__24320;
    wire N__24319;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24307;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24287;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24254;
    wire N__24251;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24241;
    wire N__24240;
    wire N__24237;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24213;
    wire N__24212;
    wire N__24209;
    wire N__24208;
    wire N__24205;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24189;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24158;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24134;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24104;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24096;
    wire N__24093;
    wire N__24092;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24053;
    wire N__24052;
    wire N__24049;
    wire N__24048;
    wire N__24045;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24013;
    wire N__24010;
    wire N__24003;
    wire N__24000;
    wire N__23999;
    wire N__23998;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23955;
    wire N__23952;
    wire N__23951;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23940;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23901;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23889;
    wire N__23886;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23867;
    wire N__23866;
    wire N__23865;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23844;
    wire N__23841;
    wire N__23832;
    wire N__23829;
    wire N__23828;
    wire N__23827;
    wire N__23826;
    wire N__23823;
    wire N__23820;
    wire N__23817;
    wire N__23814;
    wire N__23813;
    wire N__23810;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23791;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23627;
    wire N__23624;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23604;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23586;
    wire N__23583;
    wire N__23582;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23569;
    wire N__23562;
    wire N__23559;
    wire N__23558;
    wire N__23555;
    wire N__23554;
    wire N__23553;
    wire N__23552;
    wire N__23549;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23533;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23493;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23482;
    wire N__23481;
    wire N__23480;
    wire N__23479;
    wire N__23478;
    wire N__23477;
    wire N__23476;
    wire N__23475;
    wire N__23474;
    wire N__23473;
    wire N__23472;
    wire N__23471;
    wire N__23470;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23458;
    wire N__23453;
    wire N__23450;
    wire N__23445;
    wire N__23440;
    wire N__23433;
    wire N__23428;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23331;
    wire N__23328;
    wire N__23327;
    wire N__23324;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23304;
    wire N__23303;
    wire N__23298;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23261;
    wire N__23260;
    wire N__23259;
    wire N__23256;
    wire N__23251;
    wire N__23250;
    wire N__23249;
    wire N__23248;
    wire N__23245;
    wire N__23244;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23205;
    wire N__23204;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23187;
    wire N__23184;
    wire N__23183;
    wire N__23182;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23170;
    wire N__23169;
    wire N__23168;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23142;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23111;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23087;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23069;
    wire N__23064;
    wire N__23063;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23046;
    wire N__23043;
    wire N__23042;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23003;
    wire N__23002;
    wire N__23001;
    wire N__23000;
    wire N__22999;
    wire N__22998;
    wire N__22997;
    wire N__22996;
    wire N__22995;
    wire N__22994;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22950;
    wire N__22943;
    wire N__22936;
    wire N__22929;
    wire N__22924;
    wire N__22917;
    wire N__22914;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22857;
    wire N__22856;
    wire N__22855;
    wire N__22854;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22822;
    wire N__22817;
    wire N__22814;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22787;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22772;
    wire N__22769;
    wire N__22764;
    wire N__22763;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22746;
    wire N__22743;
    wire N__22742;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22724;
    wire N__22721;
    wire N__22716;
    wire N__22715;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22691;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22676;
    wire N__22673;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22654;
    wire N__22649;
    wire N__22646;
    wire N__22641;
    wire N__22638;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22630;
    wire N__22625;
    wire N__22622;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22607;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22592;
    wire N__22589;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22577;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22560;
    wire N__22557;
    wire N__22556;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22539;
    wire N__22536;
    wire N__22535;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22515;
    wire N__22512;
    wire N__22511;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22491;
    wire N__22488;
    wire N__22487;
    wire N__22484;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22467;
    wire N__22464;
    wire N__22463;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22448;
    wire N__22445;
    wire N__22440;
    wire N__22437;
    wire N__22436;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22419;
    wire N__22416;
    wire N__22415;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22395;
    wire N__22394;
    wire N__22393;
    wire N__22392;
    wire N__22391;
    wire N__22390;
    wire N__22389;
    wire N__22388;
    wire N__22387;
    wire N__22386;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22347;
    wire N__22340;
    wire N__22333;
    wire N__22326;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22303;
    wire N__22302;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22259;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22239;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22221;
    wire N__22218;
    wire N__22217;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22200;
    wire N__22197;
    wire N__22196;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22179;
    wire N__22176;
    wire N__22175;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22062;
    wire N__22059;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22026;
    wire N__22023;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21984;
    wire N__21983;
    wire N__21982;
    wire N__21981;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21973;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21965;
    wire N__21962;
    wire N__21955;
    wire N__21950;
    wire N__21945;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21929;
    wire N__21926;
    wire N__21925;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21899;
    wire N__21896;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21827;
    wire N__21826;
    wire N__21825;
    wire N__21822;
    wire N__21821;
    wire N__21820;
    wire N__21817;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21809;
    wire N__21804;
    wire N__21801;
    wire N__21790;
    wire N__21787;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21761;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21725;
    wire N__21724;
    wire N__21721;
    wire N__21716;
    wire N__21713;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21698;
    wire N__21697;
    wire N__21694;
    wire N__21689;
    wire N__21686;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21671;
    wire N__21670;
    wire N__21667;
    wire N__21662;
    wire N__21659;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21605;
    wire N__21602;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21560;
    wire N__21557;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21383;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21375;
    wire N__21372;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21356;
    wire N__21351;
    wire N__21348;
    wire N__21347;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21327;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21297;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21269;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21258;
    wire N__21255;
    wire N__21250;
    wire N__21247;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21090;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21029;
    wire N__21028;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21012;
    wire N__21009;
    wire N__21008;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20991;
    wire N__20988;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20958;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20946;
    wire N__20943;
    wire N__20942;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20925;
    wire N__20922;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20910;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20898;
    wire N__20897;
    wire N__20896;
    wire N__20895;
    wire N__20894;
    wire N__20893;
    wire N__20892;
    wire N__20891;
    wire N__20890;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20854;
    wire N__20849;
    wire N__20842;
    wire N__20835;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20778;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20742;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20727;
    wire N__20724;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20712;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20694;
    wire N__20691;
    wire N__20690;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20673;
    wire N__20670;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20658;
    wire N__20655;
    wire N__20654;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20637;
    wire N__20634;
    wire N__20633;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20616;
    wire N__20613;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20598;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20573;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20555;
    wire N__20550;
    wire N__20549;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20528;
    wire N__20523;
    wire N__20520;
    wire N__20519;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20501;
    wire N__20496;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20480;
    wire N__20477;
    wire N__20476;
    wire N__20475;
    wire N__20474;
    wire N__20471;
    wire N__20470;
    wire N__20469;
    wire N__20468;
    wire N__20467;
    wire N__20462;
    wire N__20453;
    wire N__20448;
    wire N__20445;
    wire N__20436;
    wire N__20433;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20342;
    wire N__20341;
    wire N__20338;
    wire N__20333;
    wire N__20330;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20291;
    wire N__20290;
    wire N__20287;
    wire N__20282;
    wire N__20279;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20177;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20157;
    wire N__20154;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20139;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20052;
    wire N__20049;
    wire N__20048;
    wire N__20047;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20030;
    wire N__20027;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20009;
    wire N__20006;
    wire N__20005;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19988;
    wire N__19987;
    wire N__19984;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19961;
    wire N__19960;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19928;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19908;
    wire N__19907;
    wire N__19902;
    wire N__19899;
    wire N__19898;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19881;
    wire N__19880;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19772;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19755;
    wire N__19752;
    wire N__19751;
    wire N__19746;
    wire N__19743;
    wire N__19742;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19722;
    wire N__19719;
    wire N__19718;
    wire N__19713;
    wire N__19710;
    wire N__19709;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19689;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19607;
    wire N__19604;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19520;
    wire N__19519;
    wire N__19518;
    wire N__19515;
    wire N__19514;
    wire N__19513;
    wire N__19510;
    wire N__19509;
    wire N__19506;
    wire N__19505;
    wire N__19502;
    wire N__19501;
    wire N__19500;
    wire N__19495;
    wire N__19484;
    wire N__19477;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19442;
    wire N__19439;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19422;
    wire N__19419;
    wire N__19418;
    wire N__19417;
    wire N__19414;
    wire N__19409;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19388;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19373;
    wire N__19370;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19322;
    wire N__19319;
    wire N__19318;
    wire N__19315;
    wire N__19310;
    wire N__19307;
    wire N__19302;
    wire N__19299;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19238;
    wire N__19233;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19221;
    wire N__19218;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19143;
    wire N__19140;
    wire N__19139;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19122;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19088;
    wire N__19085;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19070;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19046;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18996;
    wire N__18993;
    wire N__18992;
    wire N__18989;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18969;
    wire N__18966;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18944;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18926;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18902;
    wire N__18899;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18879;
    wire N__18876;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18868;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18854;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18842;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18827;
    wire N__18822;
    wire N__18819;
    wire N__18818;
    wire N__18815;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18788;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18747;
    wire N__18744;
    wire N__18743;
    wire N__18740;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18710;
    wire N__18707;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18680;
    wire N__18677;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18650;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18635;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18620;
    wire N__18617;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18590;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18580;
    wire N__18577;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18563;
    wire N__18560;
    wire N__18559;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18533;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18513;
    wire N__18510;
    wire N__18509;
    wire N__18506;
    wire N__18505;
    wire N__18502;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18486;
    wire N__18483;
    wire N__18480;
    wire N__18477;
    wire N__18474;
    wire N__18471;
    wire N__18468;
    wire N__18467;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18426;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18347;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18315;
    wire N__18312;
    wire N__18309;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18047;
    wire N__18042;
    wire N__18039;
    wire N__18038;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17988;
    wire N__17985;
    wire N__17982;
    wire N__17981;
    wire N__17976;
    wire N__17973;
    wire N__17972;
    wire N__17967;
    wire N__17964;
    wire N__17963;
    wire N__17958;
    wire N__17955;
    wire N__17954;
    wire N__17949;
    wire N__17946;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17934;
    wire N__17933;
    wire N__17928;
    wire N__17925;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17910;
    wire N__17907;
    wire N__17904;
    wire N__17901;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17886;
    wire N__17883;
    wire N__17880;
    wire N__17877;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17826;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17802;
    wire N__17799;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17784;
    wire N__17781;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17766;
    wire N__17763;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17748;
    wire N__17745;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17730;
    wire N__17727;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17712;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17688;
    wire N__17685;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17670;
    wire N__17667;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17655;
    wire N__17652;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17640;
    wire N__17637;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17625;
    wire N__17622;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17589;
    wire N__17586;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17571;
    wire N__17568;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17556;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17544;
    wire N__17543;
    wire N__17538;
    wire N__17535;
    wire N__17534;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17517;
    wire N__17514;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17499;
    wire N__17496;
    wire N__17495;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17463;
    wire N__17462;
    wire N__17457;
    wire N__17454;
    wire N__17453;
    wire N__17448;
    wire N__17445;
    wire N__17444;
    wire N__17439;
    wire N__17436;
    wire N__17435;
    wire N__17430;
    wire N__17427;
    wire N__17426;
    wire N__17421;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17406;
    wire N__17403;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire neo_pixel_transmitter_t0_0;
    wire neo_pixel_transmitter_t0_21;
    wire neo_pixel_transmitter_t0_7;
    wire neo_pixel_transmitter_t0_12;
    wire neo_pixel_transmitter_t0_4;
    wire neo_pixel_transmitter_t0_9;
    wire neopxl_color_prev_12;
    wire n24_adj_801_cascade_;
    wire n12414;
    wire neopxl_color_prev_6;
    wire neo_pixel_transmitter_t0_18;
    wire neo_pixel_transmitter_t0_20;
    wire neo_pixel_transmitter_t0_24;
    wire neo_pixel_transmitter_t0_31;
    wire n15_adj_841;
    wire n14_adj_842;
    wire delay_counter_0;
    wire bfn_1_22_0_;
    wire delay_counter_1;
    wire n10582;
    wire delay_counter_2;
    wire n10583;
    wire delay_counter_3;
    wire n10584;
    wire delay_counter_4;
    wire n10585;
    wire delay_counter_5;
    wire n10586;
    wire delay_counter_6;
    wire n10587;
    wire delay_counter_7;
    wire n10588;
    wire n10589;
    wire delay_counter_8;
    wire bfn_1_23_0_;
    wire delay_counter_9;
    wire n10590;
    wire delay_counter_10;
    wire n10591;
    wire delay_counter_11;
    wire n10592;
    wire delay_counter_12;
    wire n10593;
    wire delay_counter_13;
    wire n10594;
    wire delay_counter_14;
    wire n10595;
    wire n10596;
    wire n10597;
    wire bfn_1_24_0_;
    wire n10598;
    wire n10599;
    wire n10600;
    wire n10601;
    wire n10602;
    wire n10603;
    wire delay_counter_23;
    wire n10604;
    wire n10605;
    wire bfn_1_25_0_;
    wire delay_counter_25;
    wire n10606;
    wire n10607;
    wire delay_counter_27;
    wire n10608;
    wire n10609;
    wire n10610;
    wire delay_counter_30;
    wire n10611;
    wire n10612;
    wire neo_pixel_transmitter_t0_23;
    wire neo_pixel_transmitter_t0_15;
    wire neo_pixel_transmitter_t0_8;
    wire neo_pixel_transmitter_t0_2;
    wire neo_pixel_transmitter_t0_6;
    wire neo_pixel_transmitter_t0_17;
    wire neo_pixel_transmitter_t0_22;
    wire neo_pixel_transmitter_t0_10;
    wire \nx.n33 ;
    wire bfn_2_19_0_;
    wire \nx.n10669 ;
    wire \nx.n31_adj_711 ;
    wire \nx.n10670 ;
    wire \nx.n10671 ;
    wire \nx.n29_adj_714 ;
    wire \nx.n10672 ;
    wire \nx.n10673 ;
    wire \nx.n27_adj_720 ;
    wire \nx.n10674 ;
    wire \nx.n26_adj_722 ;
    wire \nx.n10675 ;
    wire \nx.n10676 ;
    wire \nx.n25_adj_724 ;
    wire bfn_2_20_0_;
    wire \nx.n24_adj_734 ;
    wire \nx.n10677 ;
    wire \nx.n23 ;
    wire \nx.n10678 ;
    wire \nx.n10679 ;
    wire \nx.one_wire_N_599_11 ;
    wire \nx.n21_adj_737 ;
    wire \nx.n10680 ;
    wire \nx.n13173 ;
    wire \nx.n10681 ;
    wire \nx.n13175 ;
    wire \nx.n10682 ;
    wire \nx.n10683 ;
    wire \nx.n10683_THRU_CRY_0_THRU_CO ;
    wire \nx.n13177 ;
    wire \nx.n18_adj_723 ;
    wire bfn_2_21_0_;
    wire \nx.n13179 ;
    wire \nx.n10684 ;
    wire \nx.n13181 ;
    wire \nx.n16_adj_672 ;
    wire \nx.n10685 ;
    wire \nx.n13183 ;
    wire \nx.n15 ;
    wire \nx.n10686 ;
    wire \nx.n13185 ;
    wire \nx.n10687 ;
    wire \nx.n13187 ;
    wire \nx.n13 ;
    wire \nx.n10688 ;
    wire \nx.n10689 ;
    wire \nx.n10689_THRU_CRY_0_THRU_CO ;
    wire \nx.n10689_THRU_CRY_1_THRU_CO ;
    wire \nx.n13189 ;
    wire \nx.n12 ;
    wire bfn_2_22_0_;
    wire \nx.n13191 ;
    wire \nx.n11 ;
    wire \nx.n10690 ;
    wire \nx.n13193 ;
    wire \nx.n10 ;
    wire \nx.n10691 ;
    wire \nx.n13195 ;
    wire \nx.n9 ;
    wire \nx.n10692 ;
    wire \nx.n13197 ;
    wire \nx.n10693 ;
    wire \nx.n13199 ;
    wire \nx.n10694 ;
    wire \nx.n10695 ;
    wire GNDG0;
    wire \nx.n10695_THRU_CRY_0_THRU_CO ;
    wire \nx.n10695_THRU_CRY_1_THRU_CO ;
    wire \nx.n13201 ;
    wire bfn_2_23_0_;
    wire \nx.n13203 ;
    wire \nx.n10696 ;
    wire \nx.n13205 ;
    wire \nx.n4_adj_710 ;
    wire \nx.n10697 ;
    wire \nx.n13207 ;
    wire \nx.n10698 ;
    wire \nx.n2 ;
    wire \nx.n13209 ;
    wire \nx.n10699 ;
    wire \nx.n6 ;
    wire neo_pixel_transmitter_t0_27;
    wire bfn_2_25_0_;
    wire \nx.n10773 ;
    wire \nx.n10774 ;
    wire \nx.n10775 ;
    wire \nx.n10776 ;
    wire \nx.n10777 ;
    wire \nx.n10778 ;
    wire \nx.n10779 ;
    wire \nx.n10780 ;
    wire bfn_2_26_0_;
    wire \nx.n10781 ;
    wire \nx.n10782 ;
    wire \nx.n1469 ;
    wire neo_pixel_transmitter_t0_14;
    wire \nx.n19_adj_725 ;
    wire \nx.n11834_cascade_ ;
    wire timer_0;
    wire bfn_3_18_0_;
    wire \nx.n10707 ;
    wire timer_2;
    wire \nx.n10708 ;
    wire \nx.n10709 ;
    wire timer_4;
    wire \nx.n10710 ;
    wire \nx.n10711 ;
    wire timer_6;
    wire \nx.n10712 ;
    wire timer_7;
    wire \nx.n10713 ;
    wire \nx.n10714 ;
    wire timer_8;
    wire bfn_3_19_0_;
    wire timer_9;
    wire \nx.n10715 ;
    wire timer_10;
    wire \nx.n10716 ;
    wire \nx.n10717 ;
    wire timer_12;
    wire \nx.n10718 ;
    wire \nx.n10719 ;
    wire timer_14;
    wire \nx.n10720 ;
    wire timer_15;
    wire \nx.n10721 ;
    wire \nx.n10722 ;
    wire bfn_3_20_0_;
    wire timer_17;
    wire \nx.n10723 ;
    wire timer_18;
    wire \nx.n10724 ;
    wire \nx.n10725 ;
    wire timer_20;
    wire \nx.n10726 ;
    wire timer_21;
    wire \nx.n10727 ;
    wire timer_22;
    wire \nx.n10728 ;
    wire timer_23;
    wire \nx.n10729 ;
    wire \nx.n10730 ;
    wire timer_24;
    wire bfn_3_21_0_;
    wire \nx.n10731 ;
    wire \nx.n10732 ;
    wire timer_27;
    wire \nx.n10733 ;
    wire \nx.n10734 ;
    wire \nx.n10735 ;
    wire \nx.n10736 ;
    wire \nx.n10737 ;
    wire timer_31;
    wire n11826_cascade_;
    wire pin_oe_1;
    wire delay_counter_17;
    wire delay_counter_15;
    wire n12382;
    wire n11828_cascade_;
    wire pin_oe_5;
    wire timer_16;
    wire neo_pixel_transmitter_t0_16;
    wire \nx.n17 ;
    wire \nx.n1309_cascade_ ;
    wire delay_counter_21;
    wire delay_counter_29;
    wire n12379;
    wire \nx.n12_adj_669 ;
    wire \nx.n1308_cascade_ ;
    wire \nx.n1334_cascade_ ;
    wire \nx.n1403_cascade_ ;
    wire \nx.n1402 ;
    wire \nx.n16_adj_727_cascade_ ;
    wire \nx.n1471 ;
    wire \nx.n1473 ;
    wire \nx.n1406 ;
    wire \nx.n1404 ;
    wire \nx.n13_adj_729 ;
    wire \nx.n18_adj_728 ;
    wire \nx.n1405 ;
    wire \nx.n1433_cascade_ ;
    wire \nx.n1472 ;
    wire \nx.n1470 ;
    wire \nx.n1403 ;
    wire \nx.n1502_cascade_ ;
    wire \nx.n1474 ;
    wire \nx.n1407 ;
    wire \nx.n1476 ;
    wire \nx.n1409 ;
    wire \nx.n1468 ;
    wire \nx.n1475 ;
    wire \nx.n1408 ;
    wire \nx.n1507_cascade_ ;
    wire \nx.n18_adj_731_cascade_ ;
    wire \nx.n20_adj_733_cascade_ ;
    wire \nx.n16_adj_732 ;
    wire \nx.n1532_cascade_ ;
    wire \nx.n1477 ;
    wire \nx.n1433 ;
    wire \nx.n1509_cascade_ ;
    wire \nx.n9729 ;
    wire \nx.n46_adj_779 ;
    wire \nx.n3 ;
    wire \nx.n7_adj_764_cascade_ ;
    wire \nx.n11864_cascade_ ;
    wire \nx.n7_adj_667 ;
    wire \nx.n103 ;
    wire \nx.n11892 ;
    wire \nx.n30_adj_712 ;
    wire \nx.n32 ;
    wire \nx.n28_adj_715 ;
    wire timer_5;
    wire neo_pixel_transmitter_t0_5;
    wire timer_1;
    wire neo_pixel_transmitter_t0_1;
    wire timer_3;
    wire neo_pixel_transmitter_t0_3;
    wire \nx.n16_adj_785 ;
    wire \nx.one_wire_N_599_4 ;
    wire \nx.n6_adj_786_cascade_ ;
    wire \nx.one_wire_N_599_5 ;
    wire \nx.n13659 ;
    wire \nx.one_wire_N_599_7 ;
    wire \nx.one_wire_N_599_8 ;
    wire \nx.one_wire_N_599_6 ;
    wire \nx.n13211 ;
    wire \nx.one_wire_N_599_10 ;
    wire \nx.one_wire_N_599_9 ;
    wire \nx.n13217_cascade_ ;
    wire \nx.n7608 ;
    wire \nx.n20_adj_726 ;
    wire timer_13;
    wire neo_pixel_transmitter_t0_13;
    wire timer_25;
    wire timer_19;
    wire pin_in_7;
    wire pin_in_6;
    wire timer_29;
    wire neo_pixel_transmitter_t0_29;
    wire neo_pixel_transmitter_t0_25;
    wire \nx.n8 ;
    wire \nx.n1205_cascade_ ;
    wire \nx.n11_adj_674 ;
    wire \nx.n1235_cascade_ ;
    wire \nx.n1203_cascade_ ;
    wire \nx.n13_adj_675 ;
    wire \nx.n1377 ;
    wire bfn_4_23_0_;
    wire \nx.n1309 ;
    wire \nx.n1376 ;
    wire \nx.n10764 ;
    wire \nx.n1308 ;
    wire \nx.n1375 ;
    wire \nx.n10765 ;
    wire \nx.n1374 ;
    wire \nx.n10766 ;
    wire \nx.n1306 ;
    wire \nx.n1373 ;
    wire \nx.n10767 ;
    wire \nx.n1372 ;
    wire \nx.n10768 ;
    wire \nx.n1371 ;
    wire \nx.n10769 ;
    wire \nx.n1303 ;
    wire \nx.n1370 ;
    wire \nx.n10770 ;
    wire \nx.n10771 ;
    wire bfn_4_24_0_;
    wire \nx.n10772 ;
    wire \nx.n1400 ;
    wire delay_counter_18;
    wire delay_counter_16;
    wire n6_adj_843;
    wire \nx.n1304 ;
    wire \nx.n1305 ;
    wire \nx.n10_adj_668_cascade_ ;
    wire \nx.n1307 ;
    wire \nx.n16 ;
    wire \nx.n1369 ;
    wire \nx.n1334 ;
    wire \nx.n1401 ;
    wire n22_adj_795;
    wire \nx.n1631_cascade_ ;
    wire \nx.n15_adj_676_cascade_ ;
    wire \nx.n22 ;
    wire \nx.n47_adj_780 ;
    wire \nx.n18 ;
    wire delay_counter_28;
    wire delay_counter_24;
    wire delay_counter_22;
    wire delay_counter_26;
    wire bfn_4_26_0_;
    wire \nx.n1509 ;
    wire \nx.n13604 ;
    wire \nx.n10783 ;
    wire \nx.n1508 ;
    wire \nx.n10784 ;
    wire \nx.n1507 ;
    wire \nx.n10785 ;
    wire \nx.n1506 ;
    wire \nx.n10786 ;
    wire \nx.n1505 ;
    wire \nx.n10787 ;
    wire \nx.n1504 ;
    wire \nx.n10788 ;
    wire \nx.n1503 ;
    wire \nx.n10789 ;
    wire \nx.n10790 ;
    wire \nx.n1502 ;
    wire bfn_4_27_0_;
    wire \nx.n1501 ;
    wire \nx.n10791 ;
    wire \nx.n1500 ;
    wire \nx.n10792 ;
    wire \nx.n1499 ;
    wire \nx.n1532 ;
    wire \nx.n10793 ;
    wire \nx.n45_adj_781 ;
    wire \nx.n19 ;
    wire pin_in_10;
    wire pin_in_11;
    wire pin_oe_6;
    wire pin_in_9;
    wire pin_in_8;
    wire n13649;
    wire timer_30;
    wire neo_pixel_transmitter_t0_30;
    wire \nx.n11946 ;
    wire \nx.n13445 ;
    wire \nx.n11948_cascade_ ;
    wire pin_in_2;
    wire pin_in_3;
    wire n13379_cascade_;
    wire \nx.n13438 ;
    wire \nx.one_wire_N_599_3 ;
    wire \nx.n11908_cascade_ ;
    wire \nx.n11926 ;
    wire \nx.n11926_cascade_ ;
    wire n7671_cascade_;
    wire \nx.one_wire_N_599_2 ;
    wire \nx.n4_adj_771 ;
    wire \nx.n9747 ;
    wire \nx.n12381 ;
    wire timer_11;
    wire pin_in_0;
    wire pin_in_1;
    wire n13378;
    wire pin_in_4;
    wire pin_in_5;
    wire n13382;
    wire n13381_cascade_;
    wire n13613;
    wire neo_pixel_transmitter_t0_11;
    wire \nx.n22_adj_749 ;
    wire neo_pixel_transmitter_t0_19;
    wire \nx.n14 ;
    wire \nx.n1109_cascade_ ;
    wire \nx.n9737_cascade_ ;
    wire \nx.n12_adj_673_cascade_ ;
    wire \nx.n1177 ;
    wire bfn_5_21_0_;
    wire \nx.n1109 ;
    wire \nx.n1176 ;
    wire \nx.n10749 ;
    wire \nx.n1108 ;
    wire \nx.n1175 ;
    wire \nx.n10750 ;
    wire \nx.n1174 ;
    wire \nx.n10751 ;
    wire \nx.n1106 ;
    wire \nx.n1173 ;
    wire \nx.n10752 ;
    wire \nx.n1172 ;
    wire \nx.n10753 ;
    wire \nx.n1104 ;
    wire \nx.n1171 ;
    wire \nx.n10754 ;
    wire \nx.n1136 ;
    wire \nx.n10755 ;
    wire \nx.n1277 ;
    wire bfn_5_22_0_;
    wire \nx.n1209 ;
    wire \nx.n1276 ;
    wire \nx.n10756 ;
    wire \nx.n1208 ;
    wire \nx.n1275 ;
    wire \nx.n10757 ;
    wire \nx.n1207 ;
    wire \nx.n1274 ;
    wire \nx.n10758 ;
    wire \nx.n1206 ;
    wire \nx.n1273 ;
    wire \nx.n10759 ;
    wire \nx.n1205 ;
    wire \nx.n1272 ;
    wire \nx.n10760 ;
    wire \nx.n1204 ;
    wire \nx.n1271 ;
    wire \nx.n10761 ;
    wire \nx.n10762 ;
    wire \nx.n10763 ;
    wire \nx.n1202 ;
    wire bfn_5_23_0_;
    wire \nx.n1301 ;
    wire delay_counter_19;
    wire delay_counter_20;
    wire n4;
    wire \nx.n1203 ;
    wire \nx.n1235 ;
    wire \nx.n1270 ;
    wire \nx.n1302 ;
    wire \nx.n49_adj_784_cascade_ ;
    wire \nx.n54 ;
    wire n7664;
    wire \nx.n30_adj_777_cascade_ ;
    wire \nx.n43_adj_783 ;
    wire bfn_5_25_0_;
    wire \nx.n1609 ;
    wire \nx.n13602 ;
    wire \nx.n10794 ;
    wire \nx.n1608 ;
    wire \nx.n10795 ;
    wire \nx.n1607 ;
    wire \nx.n10796 ;
    wire \nx.n1606 ;
    wire \nx.n10797 ;
    wire \nx.n1605 ;
    wire \nx.n10798 ;
    wire \nx.n1604 ;
    wire \nx.n10799 ;
    wire \nx.n1603 ;
    wire \nx.n10800 ;
    wire \nx.n10801 ;
    wire \nx.n1602 ;
    wire bfn_5_26_0_;
    wire \nx.n1601 ;
    wire \nx.n10802 ;
    wire \nx.n1600 ;
    wire \nx.n10803 ;
    wire \nx.n1599 ;
    wire \nx.n10804 ;
    wire \nx.n1598 ;
    wire \nx.n1631 ;
    wire \nx.n10805 ;
    wire bfn_5_27_0_;
    wire \nx.n1709 ;
    wire \nx.n10806 ;
    wire \nx.n1708 ;
    wire \nx.n10807 ;
    wire \nx.n1707 ;
    wire \nx.n10808 ;
    wire \nx.n10809 ;
    wire \nx.n10810 ;
    wire \nx.n1704 ;
    wire \nx.n10811 ;
    wire \nx.n10812 ;
    wire \nx.n10813 ;
    wire bfn_5_28_0_;
    wire \nx.n1701 ;
    wire \nx.n10814 ;
    wire \nx.n10815 ;
    wire \nx.n10816 ;
    wire \nx.n10817 ;
    wire \nx.n10818 ;
    wire \nx.n1703 ;
    wire \nx.n1706 ;
    wire \nx.n1705 ;
    wire \nx.n1700 ;
    wire \nx.n16_adj_766 ;
    wire \nx.n1702 ;
    wire \nx.n22_adj_774_cascade_ ;
    wire \nx.n1698 ;
    wire \nx.n1699 ;
    wire \nx.n1697 ;
    wire \nx.n24_adj_776_cascade_ ;
    wire \nx.n20_adj_775 ;
    wire \nx.n1730 ;
    wire \nx.n1730_cascade_ ;
    wire \nx.n13601 ;
    wire n11972;
    wire \nx.n13514 ;
    wire \nx.n13513 ;
    wire \nx.n7598 ;
    wire \nx.n11113 ;
    wire \nx.n7598_cascade_ ;
    wire timer_26;
    wire neo_pixel_transmitter_t0_26;
    wire \nx.n7 ;
    wire \nx.n10_adj_760 ;
    wire n12_adj_844;
    wire \nx.start ;
    wire \nx.n11908 ;
    wire \nx.n7564 ;
    wire update_color;
    wire \nx.n13436_cascade_ ;
    wire \nx.n3901 ;
    wire state_1_adj_791;
    wire \nx.n3901_cascade_ ;
    wire \nx.n13435 ;
    wire \nx.n1077 ;
    wire bfn_6_20_0_;
    wire \nx.n1076 ;
    wire \nx.n10743 ;
    wire \nx.n10744 ;
    wire \nx.n1074 ;
    wire \nx.n10745 ;
    wire \nx.n10746 ;
    wire \nx.n1072 ;
    wire \nx.n10747 ;
    wire \nx.n10748 ;
    wire \nx.n1103 ;
    wire \nx.n5 ;
    wire \nx.n1007 ;
    wire \nx.n1075 ;
    wire \nx.n1107 ;
    wire \nx.n1005 ;
    wire \nx.n1005_cascade_ ;
    wire \nx.n1009 ;
    wire \nx.n7_adj_690_cascade_ ;
    wire \nx.n1037 ;
    wire \nx.n1037_cascade_ ;
    wire \nx.n1073 ;
    wire \nx.n1105 ;
    wire \nx.n7899_cascade_ ;
    wire \nx.n740 ;
    wire \nx.n740_cascade_ ;
    wire \nx.n11866_cascade_ ;
    wire \nx.n838_cascade_ ;
    wire n18_adj_815;
    wire delay_counter_31;
    wire n19_adj_814;
    wire n17_adj_816;
    wire bfn_6_23_0_;
    wire \nx.n10613 ;
    wire \nx.n10614 ;
    wire \nx.n10615 ;
    wire \nx.n10616 ;
    wire \nx.n10617 ;
    wire \nx.n10618 ;
    wire \nx.n10619 ;
    wire \nx.n10620 ;
    wire bfn_6_24_0_;
    wire \nx.n10621 ;
    wire \nx.n10622 ;
    wire \nx.n10623 ;
    wire \nx.n10624 ;
    wire \nx.n10625 ;
    wire \nx.n10626 ;
    wire \nx.n10627 ;
    wire \nx.n10628 ;
    wire bfn_6_25_0_;
    wire \nx.n10629 ;
    wire \nx.n10630 ;
    wire \nx.bit_ctr_19 ;
    wire \nx.n10631 ;
    wire \nx.bit_ctr_20 ;
    wire \nx.n10632 ;
    wire \nx.bit_ctr_21 ;
    wire \nx.n10633 ;
    wire \nx.n10634 ;
    wire \nx.bit_ctr_23 ;
    wire \nx.n10635 ;
    wire \nx.n10636 ;
    wire \nx.bit_ctr_24 ;
    wire bfn_6_26_0_;
    wire \nx.bit_ctr_25 ;
    wire \nx.n10637 ;
    wire \nx.n10638 ;
    wire \nx.n10639 ;
    wire \nx.n10640 ;
    wire \nx.n10641 ;
    wire \nx.n10642 ;
    wire \nx.n10643 ;
    wire \nx.n7657 ;
    wire \nx.n7994 ;
    wire bfn_6_27_0_;
    wire \nx.n10819 ;
    wire \nx.n10820 ;
    wire \nx.n1807 ;
    wire \nx.n10821 ;
    wire \nx.n1806 ;
    wire \nx.n10822 ;
    wire \nx.n10823 ;
    wire \nx.n1804 ;
    wire \nx.n10824 ;
    wire \nx.n10825 ;
    wire \nx.n10826 ;
    wire \nx.n1802 ;
    wire bfn_6_28_0_;
    wire \nx.n1801 ;
    wire \nx.n10827 ;
    wire \nx.n10828 ;
    wire \nx.n10829 ;
    wire \nx.n10830 ;
    wire \nx.n1797 ;
    wire \nx.n10831 ;
    wire \nx.n10832 ;
    wire \nx.bit_ctr_18 ;
    wire \nx.n48_adj_778 ;
    wire \nx.n18_adj_716 ;
    wire \nx.n1799 ;
    wire \nx.n1805 ;
    wire \nx.n24_adj_717 ;
    wire \nx.n1798 ;
    wire \nx.n1808 ;
    wire \nx.n26_adj_719_cascade_ ;
    wire \nx.n1809 ;
    wire \nx.n1803 ;
    wire \nx.n1800 ;
    wire \nx.n9717_cascade_ ;
    wire \nx.n1796 ;
    wire \nx.n22_adj_718 ;
    wire \nx.n1829 ;
    wire \nx.n13605 ;
    wire pin_oe_7;
    wire \nx.neo_pixel_transmitter_done ;
    wire NEOPXL_c;
    wire \nx.n11988 ;
    wire \nx.n12451 ;
    wire \nx.bit_ctr_1 ;
    wire \nx.n13364 ;
    wire \nx.n11156_cascade_ ;
    wire \nx.n13363 ;
    wire \nx.n13619_cascade_ ;
    wire \nx.n11156 ;
    wire n11966;
    wire pin_oe_2;
    wire \nx.n13372 ;
    wire timer_28;
    wire n11353;
    wire neo_pixel_transmitter_t0_28;
    wire n9_adj_847;
    wire current_pin_7__N_153;
    wire neopxl_color_prev_14;
    wire neopxl_color_13;
    wire neopxl_color_prev_13;
    wire n11_adj_845;
    wire neopxl_color_prev_4;
    wire neopxl_color_14;
    wire \nx.n11941 ;
    wire \nx.n1008 ;
    wire \nx.n1006 ;
    wire \nx.n12837_cascade_ ;
    wire \nx.n905_cascade_ ;
    wire \nx.n12839 ;
    wire \nx.n11174 ;
    wire \nx.n11174_cascade_ ;
    wire \nx.bit_ctr_26 ;
    wire \nx.n977 ;
    wire bfn_7_22_0_;
    wire \nx.n7497 ;
    wire \nx.n976 ;
    wire \nx.n10738 ;
    wire \nx.n7899 ;
    wire \nx.n975 ;
    wire \nx.n10739 ;
    wire \nx.n974 ;
    wire \nx.n10740 ;
    wire \nx.n906 ;
    wire \nx.n973 ;
    wire \nx.n10741 ;
    wire \nx.n13594 ;
    wire \nx.n905 ;
    wire \nx.n10742 ;
    wire \nx.n4 ;
    wire \nx.n807 ;
    wire \nx.n11866 ;
    wire \nx.n838 ;
    wire \nx.n11868 ;
    wire \nx.bit_ctr_17 ;
    wire \nx.bit_ctr_22 ;
    wire \nx.n44_adj_782 ;
    wire \nx.n11912_cascade_ ;
    wire \nx.n58 ;
    wire \nx.bit_ctr_29 ;
    wire \nx.bit_ctr_30 ;
    wire \nx.bit_ctr_31 ;
    wire \nx.n9803 ;
    wire \nx.bit_ctr_27 ;
    wire \nx.bit_ctr_28 ;
    wire \nx.n11912 ;
    wire \nx.n708 ;
    wire \nx.n5703 ;
    wire n10_adj_846;
    wire neopxl_color_prev_7;
    wire neopxl_color_15;
    wire neopxl_color_prev_15;
    wire neopxl_color_6;
    wire \nx.bit_ctr_0 ;
    wire \nx.n13373 ;
    wire neopxl_color_7;
    wire n22_adj_793;
    wire \nx.n26_cascade_ ;
    wire \nx.n20 ;
    wire \nx.n28_adj_679_cascade_ ;
    wire \nx.n16_adj_678 ;
    wire \nx.n1928_cascade_ ;
    wire \nx.bit_ctr_16 ;
    wire \nx.n1977 ;
    wire bfn_7_27_0_;
    wire \nx.n1909 ;
    wire \nx.n1976 ;
    wire \nx.n10833 ;
    wire \nx.n1908 ;
    wire \nx.n1975 ;
    wire \nx.n10834 ;
    wire \nx.n1907 ;
    wire \nx.n1974 ;
    wire \nx.n10835 ;
    wire \nx.n1906 ;
    wire \nx.n1973 ;
    wire \nx.n10836 ;
    wire \nx.n10837 ;
    wire \nx.n10838 ;
    wire \nx.n10839 ;
    wire \nx.n10840 ;
    wire bfn_7_28_0_;
    wire \nx.n10841 ;
    wire \nx.n10842 ;
    wire \nx.n10843 ;
    wire \nx.n10844 ;
    wire \nx.n10845 ;
    wire \nx.n10846 ;
    wire \nx.n1895 ;
    wire \nx.n10847 ;
    wire \nx.n24 ;
    wire \nx.n1963 ;
    wire \nx.n1896 ;
    wire \nx.n1995_cascade_ ;
    wire \nx.n1965 ;
    wire \nx.n1898 ;
    wire \nx.n1964 ;
    wire \nx.n1897 ;
    wire \nx.n1971 ;
    wire \nx.n1904 ;
    wire n13360;
    wire n13361_cascade_;
    wire LED_c;
    wire neopxl_color_12;
    wire \nx.n59 ;
    wire \nx.n61_cascade_ ;
    wire \nx.n11153 ;
    wire \nx.bit_ctr_2 ;
    wire state_3_N_448_1;
    wire \nx.color_bit_N_642_4 ;
    wire \nx.n13622 ;
    wire state_0_adj_792;
    wire n7671;
    wire \nx.n7983 ;
    wire \nx.n12817 ;
    wire \nx.n12819_cascade_ ;
    wire \nx.n12821 ;
    wire \nx.n3009_cascade_ ;
    wire \nx.n2791_cascade_ ;
    wire bfn_9_21_0_;
    wire \nx.n2876 ;
    wire \nx.n11004 ;
    wire \nx.n2875 ;
    wire \nx.n11005 ;
    wire \nx.n11006 ;
    wire \nx.n11007 ;
    wire \nx.n11008 ;
    wire \nx.n11009 ;
    wire \nx.n11010 ;
    wire \nx.n11011 ;
    wire bfn_9_22_0_;
    wire \nx.n11012 ;
    wire \nx.n11013 ;
    wire \nx.n11014 ;
    wire \nx.n11015 ;
    wire \nx.n11016 ;
    wire \nx.n11017 ;
    wire \nx.n11018 ;
    wire \nx.n11019 ;
    wire bfn_9_23_0_;
    wire \nx.n11020 ;
    wire \nx.n2859 ;
    wire \nx.n11021 ;
    wire \nx.n2791 ;
    wire \nx.n2858 ;
    wire \nx.n11022 ;
    wire \nx.n11023 ;
    wire \nx.n2856 ;
    wire \nx.n11024 ;
    wire \nx.n11025 ;
    wire \nx.n11026 ;
    wire \nx.n11027 ;
    wire bfn_9_24_0_;
    wire \nx.n2792 ;
    wire neopxl_color_prev_5;
    wire neopxl_color_5;
    wire n22;
    wire \nx.n1966 ;
    wire \nx.n1899 ;
    wire \nx.n1967 ;
    wire \nx.n1900 ;
    wire \nx.n1970 ;
    wire \nx.n1903 ;
    wire \nx.n1972 ;
    wire \nx.n1905 ;
    wire bfn_9_26_0_;
    wire \nx.n10848 ;
    wire \nx.n10849 ;
    wire \nx.n10850 ;
    wire \nx.n10851 ;
    wire \nx.n10852 ;
    wire \nx.n10853 ;
    wire \nx.n10854 ;
    wire \nx.n10855 ;
    wire bfn_9_27_0_;
    wire \nx.n10856 ;
    wire \nx.n10857 ;
    wire \nx.n10858 ;
    wire \nx.n10859 ;
    wire \nx.n10860 ;
    wire \nx.n10861 ;
    wire \nx.n10862 ;
    wire \nx.n10863 ;
    wire \nx.n1994 ;
    wire bfn_9_28_0_;
    wire \nx.n1995 ;
    wire \nx.n2062 ;
    wire \nx.n2094_cascade_ ;
    wire \nx.n1901 ;
    wire \nx.n1968 ;
    wire \nx.n1969 ;
    wire \nx.n1902 ;
    wire \nx.n1928 ;
    wire \nx.n2068 ;
    wire \nx.n2001_cascade_ ;
    wire \nx.n2067 ;
    wire \nx.n2099_cascade_ ;
    wire n26_adj_798;
    wire bfn_9_29_0_;
    wire n25;
    wire n10644;
    wire n24;
    wire n10645;
    wire n23;
    wire n10646;
    wire n22_adj_799;
    wire n10647;
    wire n21;
    wire n10648;
    wire n20;
    wire n10649;
    wire n19_adj_800;
    wire n10650;
    wire n10651;
    wire n18;
    wire bfn_9_30_0_;
    wire n17;
    wire n10652;
    wire n16;
    wire n10653;
    wire n15;
    wire n10654;
    wire n14_adj_802;
    wire n10655;
    wire n13;
    wire n10656;
    wire n12;
    wire n10657;
    wire n11;
    wire n10658;
    wire n10659;
    wire n10_adj_806;
    wire bfn_9_31_0_;
    wire n9_adj_807;
    wire n10660;
    wire n8;
    wire n10661;
    wire n7_adj_808;
    wire n10662;
    wire n6_adj_809;
    wire n10663;
    wire blink_counter_21;
    wire n10664;
    wire blink_counter_22;
    wire n10665;
    wire blink_counter_23;
    wire n10666;
    wire n10667;
    wire blink_counter_24;
    wire bfn_9_32_0_;
    wire n10668;
    wire blink_counter_25;
    wire \nx.n45_adj_754_cascade_ ;
    wire \nx.n12809_cascade_ ;
    wire \nx.n12811_cascade_ ;
    wire \nx.n12813_cascade_ ;
    wire \nx.n12815 ;
    wire \nx.n43_adj_753 ;
    wire \nx.n46_cascade_ ;
    wire \nx.n13_adj_743_cascade_ ;
    wire \nx.n12775 ;
    wire \nx.n12787_cascade_ ;
    wire \nx.n12803 ;
    wire \nx.n35_adj_738 ;
    wire \nx.n2987_cascade_ ;
    wire \nx.n41_cascade_ ;
    wire \nx.n39_adj_671 ;
    wire \nx.n50_cascade_ ;
    wire \nx.n2877 ;
    wire \nx.n2857 ;
    wire \nx.n2790 ;
    wire \nx.n2889_cascade_ ;
    wire \nx.n2868 ;
    wire \nx.n2801 ;
    wire \nx.n2808 ;
    wire \nx.n40_adj_705_cascade_ ;
    wire \nx.n44_adj_721_cascade_ ;
    wire \nx.n2862 ;
    wire \nx.n2819_cascade_ ;
    wire \nx.n2874 ;
    wire \nx.n42_adj_730 ;
    wire \nx.n2807 ;
    wire \nx.n2809 ;
    wire \nx.n2809_cascade_ ;
    wire \nx.bit_ctr_7 ;
    wire \nx.n30_adj_704 ;
    wire \nx.n2802 ;
    wire \nx.n2869 ;
    wire \nx.n2802_cascade_ ;
    wire \nx.n2795 ;
    wire \nx.n2720_cascade_ ;
    wire \nx.n2788_cascade_ ;
    wire \nx.n2789 ;
    wire \nx.n26_adj_706_cascade_ ;
    wire \nx.n38_adj_713 ;
    wire \nx.n43_adj_735 ;
    wire \nx.n2777 ;
    wire bfn_10_23_0_;
    wire \nx.n2776 ;
    wire \nx.n10981 ;
    wire \nx.n2775 ;
    wire \nx.n10982 ;
    wire \nx.n10983 ;
    wire \nx.n2773 ;
    wire \nx.n10984 ;
    wire \nx.n2772 ;
    wire \nx.n10985 ;
    wire \nx.n2771 ;
    wire \nx.n10986 ;
    wire \nx.n2770 ;
    wire \nx.n10987 ;
    wire \nx.n10988 ;
    wire \nx.n2769 ;
    wire bfn_10_24_0_;
    wire \nx.n2768 ;
    wire \nx.n10989 ;
    wire \nx.n10990 ;
    wire \nx.n10991 ;
    wire \nx.n10992 ;
    wire \nx.n10993 ;
    wire \nx.n2763 ;
    wire \nx.n10994 ;
    wire \nx.n2762 ;
    wire \nx.n10995 ;
    wire \nx.n10996 ;
    wire \nx.n2761 ;
    wire bfn_10_25_0_;
    wire \nx.n2760 ;
    wire \nx.n10997 ;
    wire \nx.n2759 ;
    wire \nx.n10998 ;
    wire \nx.n2758 ;
    wire \nx.n10999 ;
    wire \nx.n2757 ;
    wire \nx.n11000 ;
    wire \nx.n2756 ;
    wire \nx.n11001 ;
    wire \nx.n11002 ;
    wire \nx.n11003 ;
    wire \nx.n2786 ;
    wire \nx.n2070 ;
    wire \nx.n9709_cascade_ ;
    wire \nx.n25 ;
    wire \nx.n26_adj_681_cascade_ ;
    wire \nx.n2027_cascade_ ;
    wire \nx.n2074 ;
    wire \nx.n2001 ;
    wire \nx.n28_adj_680 ;
    wire \nx.n1999 ;
    wire \nx.n2066 ;
    wire \nx.n2007 ;
    wire \nx.n2003 ;
    wire \nx.n2000 ;
    wire \nx.n27 ;
    wire \nx.n2004 ;
    wire \nx.n2071 ;
    wire \nx.n2103_cascade_ ;
    wire \nx.n1998 ;
    wire \nx.n2065 ;
    wire \nx.n2073 ;
    wire \nx.n2006 ;
    wire \nx.n2105_cascade_ ;
    wire \nx.n2005 ;
    wire \nx.n2072 ;
    wire \nx.n2002 ;
    wire \nx.n2069 ;
    wire \nx.n2075 ;
    wire \nx.n2008 ;
    wire \nx.n2107_cascade_ ;
    wire \nx.n24_adj_684 ;
    wire \nx.n1997 ;
    wire \nx.n2064 ;
    wire \nx.n2096_cascade_ ;
    wire \nx.bit_ctr_15 ;
    wire \nx.n2077 ;
    wire \nx.n2109_cascade_ ;
    wire \nx.n2202_cascade_ ;
    wire \nx.n18_adj_682 ;
    wire \nx.n2193_cascade_ ;
    wire \nx.n2009 ;
    wire \nx.n2076 ;
    wire \nx.n2108_cascade_ ;
    wire \nx.n1996 ;
    wire \nx.n2027 ;
    wire \nx.n2063 ;
    wire \nx.n42_adj_739_cascade_ ;
    wire \nx.n32_adj_740_cascade_ ;
    wire \nx.n44_adj_741 ;
    wire \nx.n50_adj_742 ;
    wire \nx.n47 ;
    wire \nx.n49_cascade_ ;
    wire \nx.n48 ;
    wire \nx.n3116_cascade_ ;
    wire \nx.bit_ctr_5 ;
    wire bfn_11_18_0_;
    wire \nx.n3009 ;
    wire \nx.n13600 ;
    wire \nx.n11053 ;
    wire \nx.n3008 ;
    wire \nx.n11054 ;
    wire \nx.n3007 ;
    wire \nx.n11055 ;
    wire \nx.n11056 ;
    wire \nx.n11057 ;
    wire \nx.n11058 ;
    wire \nx.n11059 ;
    wire \nx.n11060 ;
    wire bfn_11_19_0_;
    wire \nx.n11061 ;
    wire \nx.n11062 ;
    wire \nx.n11063 ;
    wire \nx.n11064 ;
    wire \nx.n11065 ;
    wire \nx.n11066 ;
    wire \nx.n11067 ;
    wire \nx.n11068 ;
    wire bfn_11_20_0_;
    wire \nx.n11069 ;
    wire \nx.n11070 ;
    wire \nx.n11071 ;
    wire \nx.n11072 ;
    wire \nx.n11073 ;
    wire \nx.n11074 ;
    wire \nx.n2987 ;
    wire \nx.n11075 ;
    wire \nx.n11076 ;
    wire bfn_11_21_0_;
    wire \nx.n11077 ;
    wire \nx.n3017 ;
    wire \nx.n11078 ;
    wire \nx.n40_adj_670 ;
    wire \nx.n2996 ;
    wire \nx.n41_adj_736 ;
    wire \nx.n2998 ;
    wire \nx.n2765 ;
    wire \nx.n41_adj_688 ;
    wire \nx.n2767 ;
    wire \nx.n2854 ;
    wire \nx.n2886_cascade_ ;
    wire \nx.n2985 ;
    wire \nx.n2774 ;
    wire \nx.n2800 ;
    wire \nx.n2867 ;
    wire \nx.n2706 ;
    wire \nx.n2706_cascade_ ;
    wire \nx.n40_adj_687 ;
    wire \nx.n2755 ;
    wire \nx.n2787 ;
    wire \nx.n2699 ;
    wire \nx.n2766 ;
    wire \nx.n2699_cascade_ ;
    wire \nx.n2701 ;
    wire \nx.n2701_cascade_ ;
    wire \nx.n42_adj_683 ;
    wire \nx.n2698 ;
    wire \nx.bit_ctr_8 ;
    wire \nx.n2698_cascade_ ;
    wire \nx.n30 ;
    wire \nx.n2693 ;
    wire \nx.n2694 ;
    wire \nx.n2693_cascade_ ;
    wire \nx.n2696 ;
    wire \nx.n37_adj_677 ;
    wire \nx.n2709 ;
    wire bfn_11_25_0_;
    wire \nx.n10881 ;
    wire \nx.n10882 ;
    wire \nx.n10883 ;
    wire \nx.n10884 ;
    wire \nx.n10885 ;
    wire \nx.n10886 ;
    wire \nx.n10887 ;
    wire \nx.n10888 ;
    wire bfn_11_26_0_;
    wire \nx.n10889 ;
    wire \nx.n10890 ;
    wire \nx.n10891 ;
    wire \nx.n10892 ;
    wire \nx.n2264 ;
    wire \nx.n10893 ;
    wire \nx.n10894 ;
    wire \nx.n10895 ;
    wire \nx.n10896 ;
    wire bfn_11_27_0_;
    wire \nx.n10897 ;
    wire \nx.n10898 ;
    wire \nx.n2263 ;
    wire \nx.n2196_cascade_ ;
    wire \nx.n2193 ;
    wire \nx.n2260 ;
    wire \nx.n29 ;
    wire \nx.n28_adj_686 ;
    wire \nx.n27_adj_691 ;
    wire \nx.n30_adj_685 ;
    wire \nx.n2126_cascade_ ;
    wire \nx.n2199_cascade_ ;
    wire \nx.n31_cascade_ ;
    wire \nx.n28_adj_692 ;
    wire \nx.bit_ctr_14 ;
    wire \nx.n2177 ;
    wire bfn_11_29_0_;
    wire \nx.n2109 ;
    wire \nx.n2176 ;
    wire \nx.n10864 ;
    wire \nx.n2108 ;
    wire \nx.n2175 ;
    wire \nx.n10865 ;
    wire \nx.n2107 ;
    wire \nx.n2174 ;
    wire \nx.n10866 ;
    wire \nx.n2106 ;
    wire \nx.n2173 ;
    wire \nx.n10867 ;
    wire \nx.n2105 ;
    wire \nx.n2172 ;
    wire \nx.n10868 ;
    wire \nx.n2104 ;
    wire \nx.n2171 ;
    wire \nx.n10869 ;
    wire \nx.n2103 ;
    wire \nx.n2170 ;
    wire \nx.n10870 ;
    wire \nx.n10871 ;
    wire bfn_11_30_0_;
    wire \nx.n10872 ;
    wire \nx.n2100 ;
    wire \nx.n2167 ;
    wire \nx.n10873 ;
    wire \nx.n10874 ;
    wire \nx.n2098 ;
    wire \nx.n2165 ;
    wire \nx.n10875 ;
    wire \nx.n2097 ;
    wire \nx.n2164 ;
    wire \nx.n10876 ;
    wire \nx.n2096 ;
    wire \nx.n2163 ;
    wire \nx.n10877 ;
    wire \nx.n2095 ;
    wire \nx.n2162 ;
    wire \nx.n10878 ;
    wire \nx.n10879 ;
    wire \nx.n2094 ;
    wire \nx.n2161 ;
    wire bfn_11_31_0_;
    wire \nx.n2093 ;
    wire \nx.n10880 ;
    wire \nx.n2192 ;
    wire \nx.n21_adj_750_cascade_ ;
    wire \nx.bit_ctr_3 ;
    wire \nx.n12781_cascade_ ;
    wire \nx.n12801 ;
    wire \nx.n27_adj_744_cascade_ ;
    wire \nx.n3209 ;
    wire \nx.n25_adj_748_cascade_ ;
    wire \nx.n12785 ;
    wire \nx.n19_adj_745 ;
    wire \nx.n12777_cascade_ ;
    wire \nx.n12779 ;
    wire \nx.n39_adj_747_cascade_ ;
    wire \nx.n12789 ;
    wire \nx.n12799 ;
    wire \nx.n29_adj_746 ;
    wire \nx.n11_adj_751 ;
    wire \nx.n41_adj_752 ;
    wire \nx.n2989 ;
    wire \nx.n3000 ;
    wire \nx.n3001 ;
    wire \nx.n3001_cascade_ ;
    wire \nx.n44 ;
    wire \nx.n3003 ;
    wire \nx.n3005 ;
    wire \nx.n2863 ;
    wire \nx.n2895_cascade_ ;
    wire \nx.n2994 ;
    wire \nx.n2799 ;
    wire \nx.n2866 ;
    wire \nx.n2898_cascade_ ;
    wire \nx.n2997 ;
    wire \nx.n2997_cascade_ ;
    wire \nx.n45 ;
    wire \nx.n2988 ;
    wire \nx.n2855 ;
    wire \nx.n2788 ;
    wire \nx.n2764 ;
    wire \nx.n2697 ;
    wire \nx.n2720 ;
    wire \nx.n2796 ;
    wire \nx.n2597_cascade_ ;
    wire \nx.n2691 ;
    wire \nx.n2690 ;
    wire \nx.n2691_cascade_ ;
    wire \nx.n2692 ;
    wire \nx.n36 ;
    wire \nx.n2700 ;
    wire \nx.n2688 ;
    wire \nx.n2689 ;
    wire \nx.n34_cascade_ ;
    wire \nx.n38 ;
    wire \nx.n37 ;
    wire \nx.n39_cascade_ ;
    wire \nx.n2621_cascade_ ;
    wire \nx.n2707 ;
    wire \nx.bit_ctr_13 ;
    wire \nx.n2277 ;
    wire \nx.n2309_cascade_ ;
    wire \nx.n9697_cascade_ ;
    wire \nx.n2273 ;
    wire \nx.n2206 ;
    wire \nx.n2209 ;
    wire \nx.n2276 ;
    wire \nx.n2695 ;
    wire \nx.n2204 ;
    wire \nx.n2271 ;
    wire \nx.n2303_cascade_ ;
    wire \nx.n2269 ;
    wire \nx.n2202 ;
    wire \nx.n2203 ;
    wire \nx.n2270 ;
    wire \nx.n2302_cascade_ ;
    wire \nx.n2401_cascade_ ;
    wire \nx.n2274 ;
    wire \nx.n2207 ;
    wire \nx.n2208 ;
    wire \nx.n2275 ;
    wire \nx.n2272 ;
    wire \nx.n2205 ;
    wire \nx.n2391_cascade_ ;
    wire \nx.n30_adj_696_cascade_ ;
    wire \nx.n2266 ;
    wire \nx.n2199 ;
    wire \nx.n2267 ;
    wire \nx.n2299_cascade_ ;
    wire \nx.n2265 ;
    wire \nx.n2197 ;
    wire \nx.n2196 ;
    wire \nx.n30_adj_694 ;
    wire \nx.n22_adj_693 ;
    wire \nx.n21_cascade_ ;
    wire \nx.n34_adj_695 ;
    wire \nx.n2268 ;
    wire \nx.n2225_cascade_ ;
    wire neopxl_color_4;
    wire n22_adj_787;
    wire \nx.n2099 ;
    wire \nx.n2166 ;
    wire \nx.n2198 ;
    wire \nx.n2169 ;
    wire \nx.n2102 ;
    wire \nx.n2201 ;
    wire \nx.n2261 ;
    wire \nx.n2194 ;
    wire \nx.n2262 ;
    wire \nx.n2195 ;
    wire \nx.n2225 ;
    wire pin_oe_4;
    wire n11970_cascade_;
    wire pin_oe_0;
    wire n11968;
    wire \nx.bit_ctr_4 ;
    wire \nx.n3177 ;
    wire bfn_13_17_0_;
    wire \nx.n3109 ;
    wire \nx.n3176 ;
    wire \nx.n11079 ;
    wire \nx.n3108 ;
    wire \nx.n3175 ;
    wire \nx.n11080 ;
    wire \nx.n3107 ;
    wire \nx.n3174 ;
    wire \nx.n11081 ;
    wire \nx.n3106 ;
    wire \nx.n3173 ;
    wire \nx.n11082 ;
    wire \nx.n3105 ;
    wire \nx.n3172 ;
    wire \nx.n11083 ;
    wire \nx.n3104 ;
    wire \nx.n3171 ;
    wire \nx.n11084 ;
    wire \nx.n3103 ;
    wire \nx.n3170 ;
    wire \nx.n11085 ;
    wire \nx.n11086 ;
    wire \nx.n3102 ;
    wire \nx.n3169 ;
    wire bfn_13_18_0_;
    wire \nx.n3101 ;
    wire \nx.n3168 ;
    wire \nx.n11087 ;
    wire \nx.n3100 ;
    wire \nx.n3167 ;
    wire \nx.n11088 ;
    wire \nx.n3099 ;
    wire \nx.n3166 ;
    wire \nx.n11089 ;
    wire \nx.n3098 ;
    wire \nx.n3165 ;
    wire \nx.n11090 ;
    wire \nx.n3097 ;
    wire \nx.n3164 ;
    wire \nx.n11091 ;
    wire \nx.n3096 ;
    wire \nx.n3163 ;
    wire \nx.n11092 ;
    wire \nx.n3095 ;
    wire \nx.n3162 ;
    wire \nx.n11093 ;
    wire \nx.n11094 ;
    wire \nx.n3094 ;
    wire \nx.n3161 ;
    wire bfn_13_19_0_;
    wire \nx.n3093 ;
    wire \nx.n3160 ;
    wire \nx.n11095 ;
    wire \nx.n3092 ;
    wire \nx.n3159 ;
    wire \nx.n11096 ;
    wire \nx.n3091 ;
    wire \nx.n3158 ;
    wire \nx.n11097 ;
    wire \nx.n3090 ;
    wire \nx.n3157 ;
    wire \nx.n11098 ;
    wire \nx.n3089 ;
    wire \nx.n3156 ;
    wire \nx.n11099 ;
    wire \nx.n3088 ;
    wire \nx.n3155 ;
    wire \nx.n11100 ;
    wire \nx.n3087 ;
    wire \nx.n3154 ;
    wire \nx.n11101 ;
    wire \nx.n11102 ;
    wire \nx.n3086 ;
    wire \nx.n3153 ;
    wire bfn_13_20_0_;
    wire \nx.n3085 ;
    wire \nx.n3152 ;
    wire \nx.n11103 ;
    wire \nx.n3084 ;
    wire \nx.n3151 ;
    wire \nx.n11104 ;
    wire \nx.n3116 ;
    wire \nx.n3083 ;
    wire \nx.n11105 ;
    wire \nx.n13280 ;
    wire \nx.n2805 ;
    wire \nx.n2872 ;
    wire \nx.n2798 ;
    wire \nx.n2865 ;
    wire \nx.n2986 ;
    wire \nx.n2991 ;
    wire \nx.n2603_cascade_ ;
    wire \nx.n2702 ;
    wire \nx.n2803 ;
    wire \nx.n2870 ;
    wire \nx.n2501_cascade_ ;
    wire \nx.n2507_cascade_ ;
    wire \nx.n2398_cascade_ ;
    wire \nx.n31_adj_700 ;
    wire \nx.n32_adj_698 ;
    wire \nx.n33_adj_699 ;
    wire \nx.n34_adj_697 ;
    wire \nx.n2324_cascade_ ;
    wire \nx.bit_ctr_12 ;
    wire \nx.n2377 ;
    wire bfn_13_26_0_;
    wire \nx.n2309 ;
    wire \nx.n2376 ;
    wire \nx.n10899 ;
    wire \nx.n2308 ;
    wire \nx.n2375 ;
    wire \nx.n10900 ;
    wire \nx.n10901 ;
    wire \nx.n2306 ;
    wire \nx.n2373 ;
    wire \nx.n10902 ;
    wire \nx.n2305 ;
    wire \nx.n2372 ;
    wire \nx.n10903 ;
    wire \nx.n2304 ;
    wire \nx.n2371 ;
    wire \nx.n10904 ;
    wire \nx.n2303 ;
    wire \nx.n2370 ;
    wire \nx.n10905 ;
    wire \nx.n10906 ;
    wire \nx.n2302 ;
    wire \nx.n2369 ;
    wire bfn_13_27_0_;
    wire \nx.n10907 ;
    wire \nx.n2300 ;
    wire \nx.n2367 ;
    wire \nx.n10908 ;
    wire \nx.n2299 ;
    wire \nx.n2366 ;
    wire \nx.n10909 ;
    wire \nx.n10910 ;
    wire \nx.n10911 ;
    wire \nx.n2296 ;
    wire \nx.n2363 ;
    wire \nx.n10912 ;
    wire \nx.n10913 ;
    wire \nx.n10914 ;
    wire \nx.n2294 ;
    wire \nx.n2361 ;
    wire bfn_13_28_0_;
    wire \nx.n2293 ;
    wire \nx.n2360 ;
    wire \nx.n10915 ;
    wire \nx.n2292 ;
    wire \nx.n2359 ;
    wire \nx.n10916 ;
    wire \nx.n2291 ;
    wire \nx.n10917 ;
    wire \nx.n3006 ;
    wire \nx.n3004 ;
    wire \nx.n3006_cascade_ ;
    wire \nx.n43 ;
    wire \nx.n2999 ;
    wire \nx.n2797 ;
    wire \nx.n2864 ;
    wire \nx.n2896_cascade_ ;
    wire \nx.n43_adj_763_cascade_ ;
    wire \nx.n38_adj_762 ;
    wire \nx.n2806 ;
    wire \nx.n2873 ;
    wire \nx.bit_ctr_6 ;
    wire \nx.n2977 ;
    wire bfn_14_19_0_;
    wire \nx.n2909 ;
    wire \nx.n2976 ;
    wire \nx.n11028 ;
    wire \nx.n2908 ;
    wire \nx.n2975 ;
    wire \nx.n11029 ;
    wire \nx.n2907 ;
    wire \nx.n2974 ;
    wire \nx.n11030 ;
    wire \nx.n2906 ;
    wire \nx.n2973 ;
    wire \nx.n11031 ;
    wire \nx.n2905 ;
    wire \nx.n2972 ;
    wire \nx.n11032 ;
    wire \nx.n2971 ;
    wire \nx.n11033 ;
    wire \nx.n11034 ;
    wire \nx.n11035 ;
    wire \nx.n2902 ;
    wire \nx.n2969 ;
    wire bfn_14_20_0_;
    wire \nx.n2901 ;
    wire \nx.n2968 ;
    wire \nx.n11036 ;
    wire \nx.n2900 ;
    wire \nx.n2967 ;
    wire \nx.n11037 ;
    wire \nx.n2899 ;
    wire \nx.n2966 ;
    wire \nx.n11038 ;
    wire \nx.n2965 ;
    wire \nx.n11039 ;
    wire \nx.n2964 ;
    wire \nx.n11040 ;
    wire \nx.n11041 ;
    wire \nx.n2895 ;
    wire \nx.n2962 ;
    wire \nx.n11042 ;
    wire \nx.n11043 ;
    wire bfn_14_21_0_;
    wire \nx.n11044 ;
    wire \nx.n2959 ;
    wire \nx.n11045 ;
    wire \nx.n11046 ;
    wire \nx.n2957 ;
    wire \nx.n11047 ;
    wire \nx.n2889 ;
    wire \nx.n2956 ;
    wire \nx.n11048 ;
    wire \nx.n2888 ;
    wire \nx.n2955 ;
    wire \nx.n11049 ;
    wire \nx.n2887 ;
    wire \nx.n2954 ;
    wire \nx.n11050 ;
    wire \nx.n11051 ;
    wire \nx.n2886 ;
    wire \nx.n2953 ;
    wire bfn_14_22_0_;
    wire \nx.n2885 ;
    wire \nx.n11052 ;
    wire \nx.n2984 ;
    wire \nx.n27_adj_757 ;
    wire \nx.n36_adj_756 ;
    wire \nx.n2708 ;
    wire \nx.n2703 ;
    wire \nx.n39_adj_689 ;
    wire \nx.n25_adj_702_cascade_ ;
    wire \nx.n34_adj_701 ;
    wire \nx.n35_adj_708 ;
    wire \nx.n32_adj_703 ;
    wire \nx.n37_adj_709_cascade_ ;
    wire \nx.n31_adj_707 ;
    wire \nx.n2423_cascade_ ;
    wire \nx.n2374 ;
    wire \nx.bit_ctr_11 ;
    wire \nx.n2477 ;
    wire bfn_14_24_0_;
    wire \nx.n10918 ;
    wire \nx.n2408 ;
    wire \nx.n2475 ;
    wire \nx.n10919 ;
    wire \nx.n2407 ;
    wire \nx.n2474 ;
    wire \nx.n10920 ;
    wire \nx.n2406 ;
    wire \nx.n2473 ;
    wire \nx.n10921 ;
    wire \nx.n2405 ;
    wire \nx.n2472 ;
    wire \nx.n10922 ;
    wire \nx.n2404 ;
    wire \nx.n2471 ;
    wire \nx.n10923 ;
    wire \nx.n2403 ;
    wire \nx.n2470 ;
    wire \nx.n10924 ;
    wire \nx.n10925 ;
    wire \nx.n2402 ;
    wire \nx.n2469 ;
    wire bfn_14_25_0_;
    wire \nx.n2401 ;
    wire \nx.n2468 ;
    wire \nx.n10926 ;
    wire \nx.n10927 ;
    wire \nx.n2399 ;
    wire \nx.n2466 ;
    wire \nx.n10928 ;
    wire \nx.n10929 ;
    wire \nx.n10930 ;
    wire \nx.n10931 ;
    wire \nx.n10932 ;
    wire \nx.n10933 ;
    wire bfn_14_26_0_;
    wire \nx.n10934 ;
    wire \nx.n10935 ;
    wire \nx.n10936 ;
    wire \nx.n2390 ;
    wire \nx.n10937 ;
    wire pin_oe_18;
    wire \nx.n2295 ;
    wire \nx.n2362 ;
    wire \nx.n2297 ;
    wire \nx.n2364 ;
    wire \nx.n2298 ;
    wire \nx.n2365 ;
    wire \nx.n2168 ;
    wire \nx.n2101 ;
    wire \nx.n2126 ;
    wire \nx.n2200 ;
    wire \nx.n2301 ;
    wire \nx.n2368 ;
    wire n7602_cascade_;
    wire n7730_cascade_;
    wire pin_oe_9;
    wire pin_oe_10;
    wire n11960;
    wire n2618;
    wire pin_oe_3;
    wire n8_adj_825_cascade_;
    wire pin_out_9;
    wire n6_adj_813_cascade_;
    wire n11974;
    wire \nx.n2890 ;
    wire \nx.n30_adj_759 ;
    wire \nx.n39_adj_761 ;
    wire \nx.n42_adj_765 ;
    wire \nx.n45_adj_769_cascade_ ;
    wire \nx.n47_adj_770 ;
    wire \nx.n2896 ;
    wire \nx.n2918_cascade_ ;
    wire \nx.n2963 ;
    wire \nx.n2970 ;
    wire \nx.n3002 ;
    wire \nx.n2995 ;
    wire \nx.n3002_cascade_ ;
    wire \nx.n42 ;
    wire \nx.n2958 ;
    wire \nx.n2891 ;
    wire \nx.n2990 ;
    wire \nx.n2804 ;
    wire \nx.n2871 ;
    wire \nx.n2903 ;
    wire \nx.n2793 ;
    wire \nx.n2860 ;
    wire \nx.n2892 ;
    wire \nx.n2960 ;
    wire \nx.n2992 ;
    wire \nx.n2794 ;
    wire \nx.n2861 ;
    wire \nx.n2819 ;
    wire \nx.n2893 ;
    wire \nx.n2898 ;
    wire \nx.n2904 ;
    wire \nx.n2893_cascade_ ;
    wire \nx.n2897 ;
    wire \nx.n41_adj_768 ;
    wire \nx.n2894 ;
    wire \nx.n2918 ;
    wire \nx.n2961 ;
    wire \nx.n2993 ;
    wire \nx.n40 ;
    wire \nx.n2609_cascade_ ;
    wire \nx.n28 ;
    wire \nx.n2606_cascade_ ;
    wire \nx.n2705 ;
    wire \nx.n2704 ;
    wire \nx.n37_adj_772_cascade_ ;
    wire \nx.n39_adj_773 ;
    wire \nx.n2522_cascade_ ;
    wire \nx.n2592_cascade_ ;
    wire \nx.n35 ;
    wire \nx.n2391 ;
    wire \nx.n2458 ;
    wire \nx.n2490_cascade_ ;
    wire \nx.n22_adj_755 ;
    wire \nx.n2324 ;
    wire \nx.n2307 ;
    wire \nx.n13321 ;
    wire \nx.n2505_cascade_ ;
    wire \nx.n2476 ;
    wire \nx.n2409 ;
    wire \nx.n2400 ;
    wire \nx.n2467 ;
    wire \nx.n2396 ;
    wire \nx.n2463 ;
    wire \nx.n2495_cascade_ ;
    wire \nx.n34_adj_758 ;
    wire \nx.n2398 ;
    wire \nx.n2465 ;
    wire \nx.n2395 ;
    wire \nx.n2462 ;
    wire \nx.n2397 ;
    wire \nx.n2464 ;
    wire \nx.n2496_cascade_ ;
    wire \nx.n2394 ;
    wire \nx.n2461 ;
    wire pin_oe_22;
    wire \nx.n2392 ;
    wire \nx.n2459 ;
    wire \nx.n2491_cascade_ ;
    wire \nx.n33_adj_767 ;
    wire \nx.n2460 ;
    wire \nx.n2393 ;
    wire \nx.n2423 ;
    wire n7992;
    wire n7602;
    wire pin_oe_11;
    wire n9;
    wire n9_cascade_;
    wire n8_adj_820_cascade_;
    wire n6_adj_805_cascade_;
    wire n1788;
    wire n9488_cascade_;
    wire n7_adj_818_cascade_;
    wire n7_adj_821;
    wire pin_out_3;
    wire pin_out_2;
    wire n13355_cascade_;
    wire n13354;
    wire n7_adj_840_cascade_;
    wire pin_out_0;
    wire n8_adj_817;
    wire pin_out_1;
    wire n11952;
    wire pin_oe_8;
    wire \nx.bit_ctr_9 ;
    wire \nx.n2677 ;
    wire bfn_16_21_0_;
    wire \nx.n2609 ;
    wire \nx.n2676 ;
    wire \nx.n10959 ;
    wire \nx.n2608 ;
    wire \nx.n2675 ;
    wire \nx.n10960 ;
    wire \nx.n2607 ;
    wire \nx.n2674 ;
    wire \nx.n10961 ;
    wire \nx.n2606 ;
    wire \nx.n2673 ;
    wire \nx.n10962 ;
    wire \nx.n2605 ;
    wire \nx.n2672 ;
    wire \nx.n10963 ;
    wire \nx.n2604 ;
    wire \nx.n2671 ;
    wire \nx.n10964 ;
    wire \nx.n2603 ;
    wire \nx.n2670 ;
    wire \nx.n10965 ;
    wire \nx.n10966 ;
    wire \nx.n2602 ;
    wire \nx.n2669 ;
    wire bfn_16_22_0_;
    wire \nx.n2601 ;
    wire \nx.n2668 ;
    wire \nx.n10967 ;
    wire \nx.n2600 ;
    wire \nx.n2667 ;
    wire \nx.n10968 ;
    wire \nx.n2599 ;
    wire \nx.n2666 ;
    wire \nx.n10969 ;
    wire \nx.n2598 ;
    wire \nx.n2665 ;
    wire \nx.n10970 ;
    wire \nx.n2597 ;
    wire \nx.n2664 ;
    wire \nx.n10971 ;
    wire \nx.n2596 ;
    wire \nx.n2663 ;
    wire \nx.n10972 ;
    wire \nx.n2595 ;
    wire \nx.n2662 ;
    wire \nx.n10973 ;
    wire \nx.n10974 ;
    wire \nx.n2594 ;
    wire \nx.n2661 ;
    wire bfn_16_23_0_;
    wire \nx.n2593 ;
    wire \nx.n2660 ;
    wire \nx.n10975 ;
    wire \nx.n2592 ;
    wire \nx.n2659 ;
    wire \nx.n10976 ;
    wire \nx.n2591 ;
    wire \nx.n2658 ;
    wire \nx.n10977 ;
    wire \nx.n2590 ;
    wire \nx.n2657 ;
    wire \nx.n10978 ;
    wire \nx.n2656 ;
    wire \nx.n10979 ;
    wire \nx.n2621 ;
    wire \nx.n10980 ;
    wire \nx.n2687 ;
    wire \nx.n2589 ;
    wire \nx.bit_ctr_10 ;
    wire \nx.n2577 ;
    wire bfn_16_24_0_;
    wire \nx.n2509 ;
    wire \nx.n2576 ;
    wire \nx.n10938 ;
    wire \nx.n2508 ;
    wire \nx.n2575 ;
    wire \nx.n10939 ;
    wire \nx.n2507 ;
    wire \nx.n2574 ;
    wire \nx.n10940 ;
    wire \nx.n2506 ;
    wire \nx.n2573 ;
    wire \nx.n10941 ;
    wire \nx.n2505 ;
    wire \nx.n2572 ;
    wire \nx.n10942 ;
    wire \nx.n2504 ;
    wire \nx.n2571 ;
    wire \nx.n10943 ;
    wire \nx.n2503 ;
    wire \nx.n2570 ;
    wire \nx.n10944 ;
    wire \nx.n10945 ;
    wire \nx.n2502 ;
    wire \nx.n2569 ;
    wire bfn_16_25_0_;
    wire \nx.n2501 ;
    wire \nx.n2568 ;
    wire \nx.n10946 ;
    wire \nx.n2500 ;
    wire \nx.n2567 ;
    wire \nx.n10947 ;
    wire \nx.n2499 ;
    wire \nx.n2566 ;
    wire \nx.n10948 ;
    wire \nx.n2498 ;
    wire \nx.n2565 ;
    wire \nx.n10949 ;
    wire \nx.n2497 ;
    wire \nx.n2564 ;
    wire \nx.n10950 ;
    wire \nx.n2496 ;
    wire \nx.n2563 ;
    wire \nx.n10951 ;
    wire \nx.n2495 ;
    wire \nx.n2562 ;
    wire \nx.n10952 ;
    wire \nx.n10953 ;
    wire \nx.n2494 ;
    wire \nx.n2561 ;
    wire bfn_16_26_0_;
    wire \nx.n2493 ;
    wire \nx.n2560 ;
    wire \nx.n10954 ;
    wire \nx.n2492 ;
    wire \nx.n2559 ;
    wire \nx.n10955 ;
    wire \nx.n2491 ;
    wire \nx.n2558 ;
    wire \nx.n10956 ;
    wire \nx.n2490 ;
    wire \nx.n2557 ;
    wire \nx.n10957 ;
    wire CONSTANT_ONE_NET;
    wire \nx.n2489 ;
    wire \nx.n2522 ;
    wire \nx.n10958 ;
    wire \nx.n2588 ;
    wire pin_oe_12;
    wire n45;
    wire bfn_17_15_0_;
    wire n10700;
    wire n10701;
    wire n10702;
    wire n10703;
    wire n10704;
    wire n10705;
    wire n13603;
    wire n10706;
    wire n7681;
    wire n11824;
    wire bfn_17_17_0_;
    wire n10575;
    wire n10576;
    wire n10577;
    wire n10578;
    wire current_pin_5;
    wire n10579;
    wire current_pin_6;
    wire n10580;
    wire n10581;
    wire current_pin_7;
    wire n7985;
    wire n7635;
    wire n9_adj_824_cascade_;
    wire n8_adj_822_cascade_;
    wire pin_out_5;
    wire pin_out_4;
    wire n13357_cascade_;
    wire n13625;
    wire n6_adj_810_cascade_;
    wire n11874;
    wire n11823;
    wire n7;
    wire n7_adj_823_cascade_;
    wire pin_oe_19;
    wire pin_out_7;
    wire pin_out_6;
    wire n13358;
    wire n3762;
    wire n11964;
    wire pin_oe_16;
    wire n11820;
    wire counter_7;
    wire counter_0;
    wire counter_6;
    wire counter_1;
    wire n10_cascade_;
    wire counter_4;
    wire counter_5;
    wire counter_2;
    wire counter_3;
    wire n14;
    wire pin_out_11;
    wire n7_adj_827_cascade_;
    wire pin_out_10;
    wire n9675_cascade_;
    wire n8_adj_832;
    wire pin_out_22__N_216;
    wire pin_out_22__N_216_cascade_;
    wire n13370;
    wire n13369;
    wire n13640_cascade_;
    wire n13628;
    wire n13540;
    wire current_pin_4;
    wire n7_adj_797_cascade_;
    wire n13551;
    wire state_7_N_167_2;
    wire n26;
    wire n11825_cascade_;
    wire pin_oe_15;
    wire n1907;
    wire state_1;
    wire state_2;
    wire n8025;
    wire n11954_cascade_;
    wire pin_oe_20;
    wire n9488;
    wire n11821;
    wire n8_adj_826;
    wire pin_out_8;
    wire n11962_cascade_;
    wire pin_oe_14;
    wire n9_adj_812;
    wire n8_adj_828;
    wire n11958_cascade_;
    wire pin_oe_21;
    wire n13652;
    wire n13536_cascade_;
    wire n13616;
    wire n13542;
    wire n7_adj_831_cascade_;
    wire n6_adj_813;
    wire n7_adj_833_cascade_;
    wire n8_adj_836;
    wire n7_adj_811;
    wire n7_adj_835_cascade_;
    wire n6_adj_810;
    wire n7_adj_839_cascade_;
    wire pin_out_18;
    wire pin_out_19;
    wire n7_adj_797;
    wire n6;
    wire n6_adj_819;
    wire n8_adj_834_cascade_;
    wire pin_out_17;
    wire n13631;
    wire pin_out_16;
    wire n13634_cascade_;
    wire n13389;
    wire n7_adj_838;
    wire n7_adj_837;
    wire pin_out_21;
    wire pin_out_20;
    wire pin_out_22;
    wire n19_adj_790_cascade_;
    wire n13388;
    wire n13375_cascade_;
    wire n13637;
    wire n8_adj_829;
    wire pin_out_12;
    wire n9675;
    wire n7_adj_830;
    wire n11789;
    wire pin_out_13;
    wire pin_out_15;
    wire pin_out_14;
    wire n13376;
    wire n11956;
    wire pin_oe_13;
    wire current_pin_2;
    wire current_pin_3;
    wire n13465;
    wire pin_in_15;
    wire pin_in_14;
    wire pin_in_13;
    wire n13643_cascade_;
    wire pin_in_12;
    wire n13646;
    wire n11822;
    wire state_0;
    wire n7730;
    wire pin_oe_17;
    wire CLK_c;
    wire pin_in_22;
    wire n13352;
    wire pin_in_17;
    wire pin_in_16;
    wire n13610;
    wire pin_in_19;
    wire pin_in_18;
    wire current_pin_1;
    wire n13607;
    wire current_pin_0;
    wire pin_in_21;
    wire pin_in_20;
    wire n19_adj_789;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__47950),
            .DIN(N__47949),
            .DOUT(N__47948),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__47950),
            .PADOUT(N__47949),
            .PADIN(N__47948),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26619),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam NEOPXL_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam NEOPXL_pad_iopad.PULLUP=1'b0;
    IO_PAD NEOPXL_pad_iopad (
            .OE(N__47941),
            .DIN(N__47940),
            .DOUT(N__47939),
            .PACKAGEPIN(NEOPXL));
    defparam NEOPXL_pad_preio.PIN_TYPE=6'b011001;
    defparam NEOPXL_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO NEOPXL_pad_preio (
            .PADOEN(N__47941),
            .PADOUT(N__47940),
            .PADIN(N__47939),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__24873),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam pin0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin0_iopad.PULLUP=1'b1;
    IO_PAD pin0_iopad (
            .OE(N__47932),
            .DIN(N__47931),
            .DOUT(N__47930),
            .PACKAGEPIN(USBPU));
    defparam pin0_preio.PIN_TYPE=6'b101001;
    defparam pin0_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin0_preio (
            .PADOEN(N__47932),
            .PADOUT(N__47931),
            .PADIN(N__47930),
            .CLOCKENABLE(),
            .DIN0(pin_in_0),
            .DIN1(),
            .DOUT0(N__39036),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__32448));
    defparam pin1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin1_iopad.PULLUP=1'b1;
    IO_PAD pin1_iopad (
            .OE(N__47923),
            .DIN(N__47922),
            .DOUT(N__47921),
            .PACKAGEPIN(ENCODER0_A));
    defparam pin1_preio.PIN_TYPE=6'b101001;
    defparam pin1_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin1_preio (
            .PADOEN(N__47923),
            .PADOUT(N__47922),
            .PADIN(N__47921),
            .CLOCKENABLE(),
            .DIN0(pin_in_1),
            .DIN1(),
            .DOUT0(N__38997),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19020));
    defparam pin10_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin10_iopad.PULLUP=1'b1;
    IO_PAD pin10_iopad (
            .OE(N__47914),
            .DIN(N__47913),
            .DOUT(N__47912),
            .PACKAGEPIN(TX));
    defparam pin10_preio.PIN_TYPE=6'b101001;
    defparam pin10_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin10_preio (
            .PADOEN(N__47914),
            .PADOUT(N__47913),
            .PADIN(N__47912),
            .CLOCKENABLE(),
            .DIN0(pin_in_10),
            .DIN1(),
            .DOUT0(N__43026),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__36756));
    defparam pin11_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin11_iopad.PULLUP=1'b1;
    IO_PAD pin11_iopad (
            .OE(N__47905),
            .DIN(N__47904),
            .DOUT(N__47903),
            .PACKAGEPIN(RX));
    defparam pin11_preio.PIN_TYPE=6'b101001;
    defparam pin11_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin11_preio (
            .PADOEN(N__47905),
            .PADOUT(N__47904),
            .PADIN(N__47903),
            .CLOCKENABLE(),
            .DIN0(pin_in_11),
            .DIN1(),
            .DOUT0(N__43056),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38364));
    defparam pin12_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin12_iopad.PULLUP=1'b1;
    IO_PAD pin12_iopad (
            .OE(N__47896),
            .DIN(N__47895),
            .DOUT(N__47894),
            .PACKAGEPIN(CS_CLK));
    defparam pin12_preio.PIN_TYPE=6'b101001;
    defparam pin12_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin12_preio (
            .PADOEN(N__47896),
            .PADOUT(N__47895),
            .PADIN(N__47894),
            .CLOCKENABLE(),
            .DIN0(pin_in_12),
            .DIN1(),
            .DOUT0(N__46185),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__40779));
    defparam pin13_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin13_iopad.PULLUP=1'b1;
    IO_PAD pin13_iopad (
            .OE(N__47887),
            .DIN(N__47886),
            .DOUT(N__47885),
            .PACKAGEPIN(CS));
    defparam pin13_preio.PIN_TYPE=6'b101001;
    defparam pin13_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin13_preio (
            .PADOEN(N__47887),
            .PADOUT(N__47886),
            .PADIN(N__47885),
            .CLOCKENABLE(),
            .DIN0(pin_in_13),
            .DIN1(),
            .DOUT0(N__45819),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__45723));
    defparam pin14_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin14_iopad.PULLUP=1'b1;
    IO_PAD pin14_iopad (
            .OE(N__47878),
            .DIN(N__47877),
            .DOUT(N__47876),
            .PACKAGEPIN(CS_MISO));
    defparam pin14_preio.PIN_TYPE=6'b101001;
    defparam pin14_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin14_preio (
            .PADOEN(N__47878),
            .PADOUT(N__47877),
            .PADIN(N__47876),
            .CLOCKENABLE(),
            .DIN0(pin_in_14),
            .DIN1(),
            .DOUT0(N__45768),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__44247));
    defparam pin15_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin15_iopad.PULLUP=1'b1;
    IO_PAD pin15_iopad (
            .OE(N__47869),
            .DIN(N__47868),
            .DOUT(N__47867),
            .PACKAGEPIN(SCL));
    defparam pin15_preio.PIN_TYPE=6'b101001;
    defparam pin15_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin15_preio (
            .PADOEN(N__47869),
            .PADOUT(N__47868),
            .PADIN(N__47867),
            .CLOCKENABLE(),
            .DIN0(pin_in_15),
            .DIN1(),
            .DOUT0(N__45798),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__44004));
    defparam pin16_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin16_iopad.PULLUP=1'b1;
    IO_PAD pin16_iopad (
            .OE(N__47860),
            .DIN(N__47859),
            .DOUT(N__47858),
            .PACKAGEPIN(SDA));
    defparam pin16_preio.PIN_TYPE=6'b101001;
    defparam pin16_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin16_preio (
            .PADOEN(N__47860),
            .PADOUT(N__47859),
            .PADIN(N__47858),
            .CLOCKENABLE(),
            .DIN0(pin_in_16),
            .DIN1(),
            .DOUT0(N__44718),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__42834));
    defparam pin17_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin17_iopad.PULLUP=1'b1;
    IO_PAD pin17_iopad (
            .OE(N__47851),
            .DIN(N__47850),
            .DOUT(N__47849),
            .PACKAGEPIN(INLC));
    defparam pin17_preio.PIN_TYPE=6'b101001;
    defparam pin17_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin17_preio (
            .PADOEN(N__47851),
            .PADOUT(N__47850),
            .PADIN(N__47849),
            .CLOCKENABLE(),
            .DIN0(pin_in_17),
            .DIN1(),
            .DOUT0(N__44751),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__46950));
    defparam pin18_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin18_iopad.PULLUP=1'b1;
    IO_PAD pin18_iopad (
            .OE(N__47842),
            .DIN(N__47841),
            .DOUT(N__47840),
            .PACKAGEPIN(INHC));
    defparam pin18_preio.PIN_TYPE=6'b101001;
    defparam pin18_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin18_preio (
            .PADOEN(N__47842),
            .PADOUT(N__47841),
            .PADIN(N__47840),
            .CLOCKENABLE(),
            .DIN0(pin_in_18),
            .DIN1(),
            .DOUT0(N__44325),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__36339));
    defparam pin19_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin19_iopad.PULLUP=1'b1;
    IO_PAD pin19_iopad (
            .OE(N__47833),
            .DIN(N__47832),
            .DOUT(N__47831),
            .PACKAGEPIN(INLB));
    defparam pin19_preio.PIN_TYPE=6'b101001;
    defparam pin19_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin19_preio (
            .PADOEN(N__47833),
            .PADOUT(N__47832),
            .PADIN(N__47831),
            .CLOCKENABLE(),
            .DIN0(pin_in_19),
            .DIN1(),
            .DOUT0(N__44292),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__42990));
    defparam pin2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin2_iopad.PULLUP=1'b1;
    IO_PAD pin2_iopad (
            .OE(N__47824),
            .DIN(N__47823),
            .DOUT(N__47822),
            .PACKAGEPIN(ENCODER0_B));
    defparam pin2_preio.PIN_TYPE=6'b101001;
    defparam pin2_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin2_preio (
            .PADOEN(N__47824),
            .PADOUT(N__47823),
            .PADIN(N__47822),
            .CLOCKENABLE(),
            .DIN0(pin_in_2),
            .DIN1(),
            .DOUT0(N__38688),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__24792));
    defparam pin20_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin20_iopad.PULLUP=1'b1;
    IO_PAD pin20_iopad (
            .OE(N__47815),
            .DIN(N__47814),
            .DOUT(N__47813),
            .PACKAGEPIN(INHB));
    defparam pin20_preio.PIN_TYPE=6'b101001;
    defparam pin20_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin20_preio (
            .PADOEN(N__47815),
            .PADOUT(N__47814),
            .PADIN(N__47813),
            .CLOCKENABLE(),
            .DIN0(pin_in_20),
            .DIN1(),
            .DOUT0(N__44619),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__43455));
    defparam pin21_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin21_iopad.PULLUP=1'b1;
    IO_PAD pin21_iopad (
            .OE(N__47806),
            .DIN(N__47805),
            .DOUT(N__47804),
            .PACKAGEPIN(INLA));
    defparam pin21_preio.PIN_TYPE=6'b101001;
    defparam pin21_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin21_preio (
            .PADOEN(N__47806),
            .PADOUT(N__47805),
            .PADIN(N__47804),
            .CLOCKENABLE(),
            .DIN0(pin_in_21),
            .DIN1(),
            .DOUT0(N__44655),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__44187));
    defparam pin22_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin22_iopad.PULLUP=1'b1;
    IO_PAD pin22_iopad (
            .OE(N__47797),
            .DIN(N__47796),
            .DOUT(N__47795),
            .PACKAGEPIN(INHA));
    defparam pin22_preio.PIN_TYPE=6'b101001;
    defparam pin22_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin22_preio (
            .PADOEN(N__47797),
            .PADOUT(N__47796),
            .PADIN(N__47795),
            .CLOCKENABLE(),
            .DIN0(pin_in_22),
            .DIN1(),
            .DOUT0(N__44595),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38616));
    defparam pin3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin3_iopad.PULLUP=1'b1;
    IO_PAD pin3_iopad (
            .OE(N__47788),
            .DIN(N__47787),
            .DOUT(N__47786),
            .PACKAGEPIN(ENCODER1_A));
    defparam pin3_preio.PIN_TYPE=6'b101001;
    defparam pin3_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin3_preio (
            .PADOEN(N__47788),
            .PADOUT(N__47787),
            .PADIN(N__47786),
            .CLOCKENABLE(),
            .DIN0(pin_in_3),
            .DIN1(),
            .DOUT0(N__38721),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__36723));
    defparam pin4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin4_iopad.PULLUP=1'b1;
    IO_PAD pin4_iopad (
            .OE(N__47779),
            .DIN(N__47778),
            .DOUT(N__47777),
            .PACKAGEPIN(ENCODER1_B));
    defparam pin4_preio.PIN_TYPE=6'b101001;
    defparam pin4_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin4_preio (
            .PADOEN(N__47779),
            .PADOUT(N__47778),
            .PADIN(N__47777),
            .CLOCKENABLE(),
            .DIN0(pin_in_4),
            .DIN1(),
            .DOUT0(N__42705),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__32475));
    defparam pin5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin5_iopad.PULLUP=1'b1;
    IO_PAD pin5_iopad (
            .OE(N__47770),
            .DIN(N__47769),
            .DOUT(N__47768),
            .PACKAGEPIN(HALL1));
    defparam pin5_preio.PIN_TYPE=6'b101001;
    defparam pin5_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin5_preio (
            .PADOEN(N__47770),
            .PADOUT(N__47769),
            .PADIN(N__47768),
            .CLOCKENABLE(),
            .DIN0(pin_in_5),
            .DIN1(),
            .DOUT0(N__42735),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19167));
    defparam pin6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin6_iopad.PULLUP=1'b1;
    IO_PAD pin6_iopad (
            .OE(N__47761),
            .DIN(N__47760),
            .DOUT(N__47759),
            .PACKAGEPIN(HALL2));
    defparam pin6_preio.PIN_TYPE=6'b101001;
    defparam pin6_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin6_preio (
            .PADOEN(N__47761),
            .PADOUT(N__47760),
            .PADIN(N__47759),
            .CLOCKENABLE(),
            .DIN0(pin_in_6),
            .DIN1(),
            .DOUT0(N__42927),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21192));
    defparam pin7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin7_iopad.PULLUP=1'b1;
    IO_PAD pin7_iopad (
            .OE(N__47752),
            .DIN(N__47751),
            .DOUT(N__47750),
            .PACKAGEPIN(HALL3));
    defparam pin7_preio.PIN_TYPE=6'b101001;
    defparam pin7_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin7_preio (
            .PADOEN(N__47752),
            .PADOUT(N__47751),
            .PADIN(N__47750),
            .CLOCKENABLE(),
            .DIN0(pin_in_7),
            .DIN1(),
            .DOUT0(N__42966),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__24396));
    defparam pin8_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin8_iopad.PULLUP=1'b1;
    IO_PAD pin8_iopad (
            .OE(N__47743),
            .DIN(N__47742),
            .DOUT(N__47741),
            .PACKAGEPIN(FAULT_N));
    defparam pin8_preio.PIN_TYPE=6'b101001;
    defparam pin8_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin8_preio (
            .PADOEN(N__47743),
            .PADOUT(N__47742),
            .PADIN(N__47741),
            .CLOCKENABLE(),
            .DIN0(pin_in_8),
            .DIN1(),
            .DOUT0(N__43353),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__38952));
    defparam pin9_iopad.IO_STANDARD="SB_LVCMOS";
    defparam pin9_iopad.PULLUP=1'b1;
    IO_PAD pin9_iopad (
            .OE(N__47734),
            .DIN(N__47733),
            .DOUT(N__47732),
            .PACKAGEPIN(DE));
    defparam pin9_preio.PIN_TYPE=6'b101001;
    defparam pin9_preio.NEG_TRIGGER=1'b0;
    PRE_IO pin9_preio (
            .PADOEN(N__47734),
            .PADOUT(N__47733),
            .PADIN(N__47732),
            .CLOCKENABLE(),
            .DIN0(pin_in_9),
            .DIN1(),
            .DOUT0(N__36699),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__36777));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__47725),
            .DIN(N__47724),
            .DOUT(N__47723),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__47725),
            .PADOUT(N__47724),
            .PADIN(N__47723),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__11563 (
            .O(N__47706),
            .I(N__47703));
    LocalMux I__11562 (
            .O(N__47703),
            .I(N__47700));
    Odrv12 I__11561 (
            .O(N__47700),
            .I(n11822));
    CascadeMux I__11560 (
            .O(N__47697),
            .I(N__47690));
    CascadeMux I__11559 (
            .O(N__47696),
            .I(N__47687));
    CascadeMux I__11558 (
            .O(N__47695),
            .I(N__47684));
    CascadeMux I__11557 (
            .O(N__47694),
            .I(N__47681));
    InMux I__11556 (
            .O(N__47693),
            .I(N__47678));
    InMux I__11555 (
            .O(N__47690),
            .I(N__47669));
    InMux I__11554 (
            .O(N__47687),
            .I(N__47660));
    InMux I__11553 (
            .O(N__47684),
            .I(N__47654));
    InMux I__11552 (
            .O(N__47681),
            .I(N__47651));
    LocalMux I__11551 (
            .O(N__47678),
            .I(N__47648));
    CascadeMux I__11550 (
            .O(N__47677),
            .I(N__47643));
    CascadeMux I__11549 (
            .O(N__47676),
            .I(N__47638));
    CascadeMux I__11548 (
            .O(N__47675),
            .I(N__47632));
    CascadeMux I__11547 (
            .O(N__47674),
            .I(N__47628));
    InMux I__11546 (
            .O(N__47673),
            .I(N__47625));
    InMux I__11545 (
            .O(N__47672),
            .I(N__47621));
    LocalMux I__11544 (
            .O(N__47669),
            .I(N__47618));
    InMux I__11543 (
            .O(N__47668),
            .I(N__47611));
    InMux I__11542 (
            .O(N__47667),
            .I(N__47611));
    InMux I__11541 (
            .O(N__47666),
            .I(N__47611));
    InMux I__11540 (
            .O(N__47665),
            .I(N__47607));
    InMux I__11539 (
            .O(N__47664),
            .I(N__47604));
    CascadeMux I__11538 (
            .O(N__47663),
            .I(N__47601));
    LocalMux I__11537 (
            .O(N__47660),
            .I(N__47595));
    CascadeMux I__11536 (
            .O(N__47659),
            .I(N__47591));
    CascadeMux I__11535 (
            .O(N__47658),
            .I(N__47587));
    CascadeMux I__11534 (
            .O(N__47657),
            .I(N__47578));
    LocalMux I__11533 (
            .O(N__47654),
            .I(N__47570));
    LocalMux I__11532 (
            .O(N__47651),
            .I(N__47570));
    Span4Mux_h I__11531 (
            .O(N__47648),
            .I(N__47570));
    InMux I__11530 (
            .O(N__47647),
            .I(N__47563));
    InMux I__11529 (
            .O(N__47646),
            .I(N__47563));
    InMux I__11528 (
            .O(N__47643),
            .I(N__47563));
    InMux I__11527 (
            .O(N__47642),
            .I(N__47560));
    InMux I__11526 (
            .O(N__47641),
            .I(N__47555));
    InMux I__11525 (
            .O(N__47638),
            .I(N__47555));
    InMux I__11524 (
            .O(N__47637),
            .I(N__47550));
    InMux I__11523 (
            .O(N__47636),
            .I(N__47550));
    CascadeMux I__11522 (
            .O(N__47635),
            .I(N__47546));
    InMux I__11521 (
            .O(N__47632),
            .I(N__47543));
    CascadeMux I__11520 (
            .O(N__47631),
            .I(N__47540));
    InMux I__11519 (
            .O(N__47628),
            .I(N__47536));
    LocalMux I__11518 (
            .O(N__47625),
            .I(N__47533));
    InMux I__11517 (
            .O(N__47624),
            .I(N__47530));
    LocalMux I__11516 (
            .O(N__47621),
            .I(N__47523));
    Span4Mux_v I__11515 (
            .O(N__47618),
            .I(N__47523));
    LocalMux I__11514 (
            .O(N__47611),
            .I(N__47523));
    CascadeMux I__11513 (
            .O(N__47610),
            .I(N__47520));
    LocalMux I__11512 (
            .O(N__47607),
            .I(N__47509));
    LocalMux I__11511 (
            .O(N__47604),
            .I(N__47509));
    InMux I__11510 (
            .O(N__47601),
            .I(N__47506));
    CascadeMux I__11509 (
            .O(N__47600),
            .I(N__47503));
    CascadeMux I__11508 (
            .O(N__47599),
            .I(N__47499));
    InMux I__11507 (
            .O(N__47598),
            .I(N__47496));
    Span4Mux_h I__11506 (
            .O(N__47595),
            .I(N__47493));
    InMux I__11505 (
            .O(N__47594),
            .I(N__47490));
    InMux I__11504 (
            .O(N__47591),
            .I(N__47485));
    InMux I__11503 (
            .O(N__47590),
            .I(N__47475));
    InMux I__11502 (
            .O(N__47587),
            .I(N__47470));
    InMux I__11501 (
            .O(N__47586),
            .I(N__47470));
    InMux I__11500 (
            .O(N__47585),
            .I(N__47461));
    InMux I__11499 (
            .O(N__47584),
            .I(N__47461));
    InMux I__11498 (
            .O(N__47583),
            .I(N__47461));
    InMux I__11497 (
            .O(N__47582),
            .I(N__47461));
    InMux I__11496 (
            .O(N__47581),
            .I(N__47456));
    InMux I__11495 (
            .O(N__47578),
            .I(N__47453));
    CascadeMux I__11494 (
            .O(N__47577),
            .I(N__47450));
    Span4Mux_v I__11493 (
            .O(N__47570),
            .I(N__47447));
    LocalMux I__11492 (
            .O(N__47563),
            .I(N__47444));
    LocalMux I__11491 (
            .O(N__47560),
            .I(N__47437));
    LocalMux I__11490 (
            .O(N__47555),
            .I(N__47437));
    LocalMux I__11489 (
            .O(N__47550),
            .I(N__47437));
    InMux I__11488 (
            .O(N__47549),
            .I(N__47432));
    InMux I__11487 (
            .O(N__47546),
            .I(N__47432));
    LocalMux I__11486 (
            .O(N__47543),
            .I(N__47428));
    InMux I__11485 (
            .O(N__47540),
            .I(N__47425));
    InMux I__11484 (
            .O(N__47539),
            .I(N__47422));
    LocalMux I__11483 (
            .O(N__47536),
            .I(N__47415));
    Span4Mux_h I__11482 (
            .O(N__47533),
            .I(N__47415));
    LocalMux I__11481 (
            .O(N__47530),
            .I(N__47415));
    Span4Mux_h I__11480 (
            .O(N__47523),
            .I(N__47412));
    InMux I__11479 (
            .O(N__47520),
            .I(N__47407));
    InMux I__11478 (
            .O(N__47519),
            .I(N__47407));
    InMux I__11477 (
            .O(N__47518),
            .I(N__47402));
    InMux I__11476 (
            .O(N__47517),
            .I(N__47402));
    InMux I__11475 (
            .O(N__47516),
            .I(N__47397));
    InMux I__11474 (
            .O(N__47515),
            .I(N__47397));
    InMux I__11473 (
            .O(N__47514),
            .I(N__47394));
    Span4Mux_h I__11472 (
            .O(N__47509),
            .I(N__47391));
    LocalMux I__11471 (
            .O(N__47506),
            .I(N__47388));
    InMux I__11470 (
            .O(N__47503),
            .I(N__47385));
    InMux I__11469 (
            .O(N__47502),
            .I(N__47380));
    InMux I__11468 (
            .O(N__47499),
            .I(N__47380));
    LocalMux I__11467 (
            .O(N__47496),
            .I(N__47377));
    Span4Mux_v I__11466 (
            .O(N__47493),
            .I(N__47372));
    LocalMux I__11465 (
            .O(N__47490),
            .I(N__47372));
    CascadeMux I__11464 (
            .O(N__47489),
            .I(N__47369));
    CascadeMux I__11463 (
            .O(N__47488),
            .I(N__47364));
    LocalMux I__11462 (
            .O(N__47485),
            .I(N__47360));
    InMux I__11461 (
            .O(N__47484),
            .I(N__47355));
    InMux I__11460 (
            .O(N__47483),
            .I(N__47355));
    InMux I__11459 (
            .O(N__47482),
            .I(N__47350));
    InMux I__11458 (
            .O(N__47481),
            .I(N__47350));
    InMux I__11457 (
            .O(N__47480),
            .I(N__47347));
    InMux I__11456 (
            .O(N__47479),
            .I(N__47344));
    InMux I__11455 (
            .O(N__47478),
            .I(N__47341));
    LocalMux I__11454 (
            .O(N__47475),
            .I(N__47336));
    LocalMux I__11453 (
            .O(N__47470),
            .I(N__47336));
    LocalMux I__11452 (
            .O(N__47461),
            .I(N__47333));
    CascadeMux I__11451 (
            .O(N__47460),
            .I(N__47330));
    CascadeMux I__11450 (
            .O(N__47459),
            .I(N__47326));
    LocalMux I__11449 (
            .O(N__47456),
            .I(N__47318));
    LocalMux I__11448 (
            .O(N__47453),
            .I(N__47318));
    InMux I__11447 (
            .O(N__47450),
            .I(N__47315));
    Span4Mux_v I__11446 (
            .O(N__47447),
            .I(N__47308));
    Span4Mux_h I__11445 (
            .O(N__47444),
            .I(N__47308));
    Span4Mux_h I__11444 (
            .O(N__47437),
            .I(N__47308));
    LocalMux I__11443 (
            .O(N__47432),
            .I(N__47305));
    CascadeMux I__11442 (
            .O(N__47431),
            .I(N__47302));
    Span4Mux_v I__11441 (
            .O(N__47428),
            .I(N__47296));
    LocalMux I__11440 (
            .O(N__47425),
            .I(N__47277));
    LocalMux I__11439 (
            .O(N__47422),
            .I(N__47277));
    Sp12to4 I__11438 (
            .O(N__47415),
            .I(N__47277));
    Sp12to4 I__11437 (
            .O(N__47412),
            .I(N__47277));
    LocalMux I__11436 (
            .O(N__47407),
            .I(N__47277));
    LocalMux I__11435 (
            .O(N__47402),
            .I(N__47277));
    LocalMux I__11434 (
            .O(N__47397),
            .I(N__47277));
    LocalMux I__11433 (
            .O(N__47394),
            .I(N__47277));
    Sp12to4 I__11432 (
            .O(N__47391),
            .I(N__47277));
    Span4Mux_h I__11431 (
            .O(N__47388),
            .I(N__47272));
    LocalMux I__11430 (
            .O(N__47385),
            .I(N__47272));
    LocalMux I__11429 (
            .O(N__47380),
            .I(N__47269));
    Span4Mux_h I__11428 (
            .O(N__47377),
            .I(N__47264));
    Span4Mux_v I__11427 (
            .O(N__47372),
            .I(N__47264));
    InMux I__11426 (
            .O(N__47369),
            .I(N__47259));
    InMux I__11425 (
            .O(N__47368),
            .I(N__47259));
    InMux I__11424 (
            .O(N__47367),
            .I(N__47256));
    InMux I__11423 (
            .O(N__47364),
            .I(N__47251));
    InMux I__11422 (
            .O(N__47363),
            .I(N__47251));
    Span4Mux_h I__11421 (
            .O(N__47360),
            .I(N__47234));
    LocalMux I__11420 (
            .O(N__47355),
            .I(N__47234));
    LocalMux I__11419 (
            .O(N__47350),
            .I(N__47234));
    LocalMux I__11418 (
            .O(N__47347),
            .I(N__47234));
    LocalMux I__11417 (
            .O(N__47344),
            .I(N__47234));
    LocalMux I__11416 (
            .O(N__47341),
            .I(N__47234));
    Span4Mux_h I__11415 (
            .O(N__47336),
            .I(N__47234));
    Span4Mux_v I__11414 (
            .O(N__47333),
            .I(N__47234));
    InMux I__11413 (
            .O(N__47330),
            .I(N__47229));
    InMux I__11412 (
            .O(N__47329),
            .I(N__47229));
    InMux I__11411 (
            .O(N__47326),
            .I(N__47226));
    InMux I__11410 (
            .O(N__47325),
            .I(N__47221));
    InMux I__11409 (
            .O(N__47324),
            .I(N__47221));
    InMux I__11408 (
            .O(N__47323),
            .I(N__47218));
    Span4Mux_v I__11407 (
            .O(N__47318),
            .I(N__47215));
    LocalMux I__11406 (
            .O(N__47315),
            .I(N__47208));
    Span4Mux_v I__11405 (
            .O(N__47308),
            .I(N__47208));
    Span4Mux_h I__11404 (
            .O(N__47305),
            .I(N__47208));
    InMux I__11403 (
            .O(N__47302),
            .I(N__47199));
    InMux I__11402 (
            .O(N__47301),
            .I(N__47199));
    InMux I__11401 (
            .O(N__47300),
            .I(N__47199));
    InMux I__11400 (
            .O(N__47299),
            .I(N__47199));
    Sp12to4 I__11399 (
            .O(N__47296),
            .I(N__47194));
    Span12Mux_v I__11398 (
            .O(N__47277),
            .I(N__47194));
    Span4Mux_h I__11397 (
            .O(N__47272),
            .I(N__47183));
    Span4Mux_v I__11396 (
            .O(N__47269),
            .I(N__47183));
    Span4Mux_h I__11395 (
            .O(N__47264),
            .I(N__47183));
    LocalMux I__11394 (
            .O(N__47259),
            .I(N__47183));
    LocalMux I__11393 (
            .O(N__47256),
            .I(N__47183));
    LocalMux I__11392 (
            .O(N__47251),
            .I(N__47176));
    Span4Mux_v I__11391 (
            .O(N__47234),
            .I(N__47176));
    LocalMux I__11390 (
            .O(N__47229),
            .I(N__47176));
    LocalMux I__11389 (
            .O(N__47226),
            .I(state_0));
    LocalMux I__11388 (
            .O(N__47221),
            .I(state_0));
    LocalMux I__11387 (
            .O(N__47218),
            .I(state_0));
    Odrv4 I__11386 (
            .O(N__47215),
            .I(state_0));
    Odrv4 I__11385 (
            .O(N__47208),
            .I(state_0));
    LocalMux I__11384 (
            .O(N__47199),
            .I(state_0));
    Odrv12 I__11383 (
            .O(N__47194),
            .I(state_0));
    Odrv4 I__11382 (
            .O(N__47183),
            .I(state_0));
    Odrv4 I__11381 (
            .O(N__47176),
            .I(state_0));
    InMux I__11380 (
            .O(N__47157),
            .I(N__47150));
    InMux I__11379 (
            .O(N__47156),
            .I(N__47143));
    InMux I__11378 (
            .O(N__47155),
            .I(N__47140));
    InMux I__11377 (
            .O(N__47154),
            .I(N__47137));
    InMux I__11376 (
            .O(N__47153),
            .I(N__47134));
    LocalMux I__11375 (
            .O(N__47150),
            .I(N__47131));
    CascadeMux I__11374 (
            .O(N__47149),
            .I(N__47127));
    InMux I__11373 (
            .O(N__47148),
            .I(N__47116));
    InMux I__11372 (
            .O(N__47147),
            .I(N__47113));
    InMux I__11371 (
            .O(N__47146),
            .I(N__47110));
    LocalMux I__11370 (
            .O(N__47143),
            .I(N__47107));
    LocalMux I__11369 (
            .O(N__47140),
            .I(N__47102));
    LocalMux I__11368 (
            .O(N__47137),
            .I(N__47102));
    LocalMux I__11367 (
            .O(N__47134),
            .I(N__47099));
    Span4Mux_v I__11366 (
            .O(N__47131),
            .I(N__47096));
    InMux I__11365 (
            .O(N__47130),
            .I(N__47093));
    InMux I__11364 (
            .O(N__47127),
            .I(N__47090));
    InMux I__11363 (
            .O(N__47126),
            .I(N__47085));
    InMux I__11362 (
            .O(N__47125),
            .I(N__47085));
    InMux I__11361 (
            .O(N__47124),
            .I(N__47082));
    InMux I__11360 (
            .O(N__47123),
            .I(N__47079));
    InMux I__11359 (
            .O(N__47122),
            .I(N__47076));
    InMux I__11358 (
            .O(N__47121),
            .I(N__47073));
    InMux I__11357 (
            .O(N__47120),
            .I(N__47069));
    InMux I__11356 (
            .O(N__47119),
            .I(N__47066));
    LocalMux I__11355 (
            .O(N__47116),
            .I(N__47061));
    LocalMux I__11354 (
            .O(N__47113),
            .I(N__47061));
    LocalMux I__11353 (
            .O(N__47110),
            .I(N__47058));
    Span4Mux_h I__11352 (
            .O(N__47107),
            .I(N__47053));
    Span4Mux_v I__11351 (
            .O(N__47102),
            .I(N__47053));
    Span4Mux_h I__11350 (
            .O(N__47099),
            .I(N__47048));
    Span4Mux_h I__11349 (
            .O(N__47096),
            .I(N__47048));
    LocalMux I__11348 (
            .O(N__47093),
            .I(N__47043));
    LocalMux I__11347 (
            .O(N__47090),
            .I(N__47043));
    LocalMux I__11346 (
            .O(N__47085),
            .I(N__47040));
    LocalMux I__11345 (
            .O(N__47082),
            .I(N__47034));
    LocalMux I__11344 (
            .O(N__47079),
            .I(N__47031));
    LocalMux I__11343 (
            .O(N__47076),
            .I(N__47028));
    LocalMux I__11342 (
            .O(N__47073),
            .I(N__47025));
    InMux I__11341 (
            .O(N__47072),
            .I(N__47022));
    LocalMux I__11340 (
            .O(N__47069),
            .I(N__47019));
    LocalMux I__11339 (
            .O(N__47066),
            .I(N__47014));
    Span4Mux_v I__11338 (
            .O(N__47061),
            .I(N__47014));
    Span4Mux_h I__11337 (
            .O(N__47058),
            .I(N__47005));
    Span4Mux_v I__11336 (
            .O(N__47053),
            .I(N__47005));
    Span4Mux_h I__11335 (
            .O(N__47048),
            .I(N__47005));
    Span4Mux_h I__11334 (
            .O(N__47043),
            .I(N__47005));
    Span12Mux_v I__11333 (
            .O(N__47040),
            .I(N__47002));
    InMux I__11332 (
            .O(N__47039),
            .I(N__46999));
    InMux I__11331 (
            .O(N__47038),
            .I(N__46996));
    InMux I__11330 (
            .O(N__47037),
            .I(N__46993));
    Span4Mux_h I__11329 (
            .O(N__47034),
            .I(N__46990));
    Span4Mux_v I__11328 (
            .O(N__47031),
            .I(N__46985));
    Span4Mux_v I__11327 (
            .O(N__47028),
            .I(N__46985));
    Span12Mux_s9_h I__11326 (
            .O(N__47025),
            .I(N__46982));
    LocalMux I__11325 (
            .O(N__47022),
            .I(N__46975));
    Span4Mux_v I__11324 (
            .O(N__47019),
            .I(N__46975));
    Span4Mux_h I__11323 (
            .O(N__47014),
            .I(N__46975));
    Span4Mux_v I__11322 (
            .O(N__47005),
            .I(N__46972));
    Span12Mux_h I__11321 (
            .O(N__47002),
            .I(N__46969));
    LocalMux I__11320 (
            .O(N__46999),
            .I(n7730));
    LocalMux I__11319 (
            .O(N__46996),
            .I(n7730));
    LocalMux I__11318 (
            .O(N__46993),
            .I(n7730));
    Odrv4 I__11317 (
            .O(N__46990),
            .I(n7730));
    Odrv4 I__11316 (
            .O(N__46985),
            .I(n7730));
    Odrv12 I__11315 (
            .O(N__46982),
            .I(n7730));
    Odrv4 I__11314 (
            .O(N__46975),
            .I(n7730));
    Odrv4 I__11313 (
            .O(N__46972),
            .I(n7730));
    Odrv12 I__11312 (
            .O(N__46969),
            .I(n7730));
    IoInMux I__11311 (
            .O(N__46950),
            .I(N__46947));
    LocalMux I__11310 (
            .O(N__46947),
            .I(N__46944));
    Span4Mux_s3_v I__11309 (
            .O(N__46944),
            .I(N__46941));
    Sp12to4 I__11308 (
            .O(N__46941),
            .I(N__46938));
    Span12Mux_s11_h I__11307 (
            .O(N__46938),
            .I(N__46935));
    Span12Mux_v I__11306 (
            .O(N__46935),
            .I(N__46931));
    InMux I__11305 (
            .O(N__46934),
            .I(N__46928));
    Odrv12 I__11304 (
            .O(N__46931),
            .I(pin_oe_17));
    LocalMux I__11303 (
            .O(N__46928),
            .I(pin_oe_17));
    ClkMux I__11302 (
            .O(N__46923),
            .I(N__46668));
    ClkMux I__11301 (
            .O(N__46922),
            .I(N__46668));
    ClkMux I__11300 (
            .O(N__46921),
            .I(N__46668));
    ClkMux I__11299 (
            .O(N__46920),
            .I(N__46668));
    ClkMux I__11298 (
            .O(N__46919),
            .I(N__46668));
    ClkMux I__11297 (
            .O(N__46918),
            .I(N__46668));
    ClkMux I__11296 (
            .O(N__46917),
            .I(N__46668));
    ClkMux I__11295 (
            .O(N__46916),
            .I(N__46668));
    ClkMux I__11294 (
            .O(N__46915),
            .I(N__46668));
    ClkMux I__11293 (
            .O(N__46914),
            .I(N__46668));
    ClkMux I__11292 (
            .O(N__46913),
            .I(N__46668));
    ClkMux I__11291 (
            .O(N__46912),
            .I(N__46668));
    ClkMux I__11290 (
            .O(N__46911),
            .I(N__46668));
    ClkMux I__11289 (
            .O(N__46910),
            .I(N__46668));
    ClkMux I__11288 (
            .O(N__46909),
            .I(N__46668));
    ClkMux I__11287 (
            .O(N__46908),
            .I(N__46668));
    ClkMux I__11286 (
            .O(N__46907),
            .I(N__46668));
    ClkMux I__11285 (
            .O(N__46906),
            .I(N__46668));
    ClkMux I__11284 (
            .O(N__46905),
            .I(N__46668));
    ClkMux I__11283 (
            .O(N__46904),
            .I(N__46668));
    ClkMux I__11282 (
            .O(N__46903),
            .I(N__46668));
    ClkMux I__11281 (
            .O(N__46902),
            .I(N__46668));
    ClkMux I__11280 (
            .O(N__46901),
            .I(N__46668));
    ClkMux I__11279 (
            .O(N__46900),
            .I(N__46668));
    ClkMux I__11278 (
            .O(N__46899),
            .I(N__46668));
    ClkMux I__11277 (
            .O(N__46898),
            .I(N__46668));
    ClkMux I__11276 (
            .O(N__46897),
            .I(N__46668));
    ClkMux I__11275 (
            .O(N__46896),
            .I(N__46668));
    ClkMux I__11274 (
            .O(N__46895),
            .I(N__46668));
    ClkMux I__11273 (
            .O(N__46894),
            .I(N__46668));
    ClkMux I__11272 (
            .O(N__46893),
            .I(N__46668));
    ClkMux I__11271 (
            .O(N__46892),
            .I(N__46668));
    ClkMux I__11270 (
            .O(N__46891),
            .I(N__46668));
    ClkMux I__11269 (
            .O(N__46890),
            .I(N__46668));
    ClkMux I__11268 (
            .O(N__46889),
            .I(N__46668));
    ClkMux I__11267 (
            .O(N__46888),
            .I(N__46668));
    ClkMux I__11266 (
            .O(N__46887),
            .I(N__46668));
    ClkMux I__11265 (
            .O(N__46886),
            .I(N__46668));
    ClkMux I__11264 (
            .O(N__46885),
            .I(N__46668));
    ClkMux I__11263 (
            .O(N__46884),
            .I(N__46668));
    ClkMux I__11262 (
            .O(N__46883),
            .I(N__46668));
    ClkMux I__11261 (
            .O(N__46882),
            .I(N__46668));
    ClkMux I__11260 (
            .O(N__46881),
            .I(N__46668));
    ClkMux I__11259 (
            .O(N__46880),
            .I(N__46668));
    ClkMux I__11258 (
            .O(N__46879),
            .I(N__46668));
    ClkMux I__11257 (
            .O(N__46878),
            .I(N__46668));
    ClkMux I__11256 (
            .O(N__46877),
            .I(N__46668));
    ClkMux I__11255 (
            .O(N__46876),
            .I(N__46668));
    ClkMux I__11254 (
            .O(N__46875),
            .I(N__46668));
    ClkMux I__11253 (
            .O(N__46874),
            .I(N__46668));
    ClkMux I__11252 (
            .O(N__46873),
            .I(N__46668));
    ClkMux I__11251 (
            .O(N__46872),
            .I(N__46668));
    ClkMux I__11250 (
            .O(N__46871),
            .I(N__46668));
    ClkMux I__11249 (
            .O(N__46870),
            .I(N__46668));
    ClkMux I__11248 (
            .O(N__46869),
            .I(N__46668));
    ClkMux I__11247 (
            .O(N__46868),
            .I(N__46668));
    ClkMux I__11246 (
            .O(N__46867),
            .I(N__46668));
    ClkMux I__11245 (
            .O(N__46866),
            .I(N__46668));
    ClkMux I__11244 (
            .O(N__46865),
            .I(N__46668));
    ClkMux I__11243 (
            .O(N__46864),
            .I(N__46668));
    ClkMux I__11242 (
            .O(N__46863),
            .I(N__46668));
    ClkMux I__11241 (
            .O(N__46862),
            .I(N__46668));
    ClkMux I__11240 (
            .O(N__46861),
            .I(N__46668));
    ClkMux I__11239 (
            .O(N__46860),
            .I(N__46668));
    ClkMux I__11238 (
            .O(N__46859),
            .I(N__46668));
    ClkMux I__11237 (
            .O(N__46858),
            .I(N__46668));
    ClkMux I__11236 (
            .O(N__46857),
            .I(N__46668));
    ClkMux I__11235 (
            .O(N__46856),
            .I(N__46668));
    ClkMux I__11234 (
            .O(N__46855),
            .I(N__46668));
    ClkMux I__11233 (
            .O(N__46854),
            .I(N__46668));
    ClkMux I__11232 (
            .O(N__46853),
            .I(N__46668));
    ClkMux I__11231 (
            .O(N__46852),
            .I(N__46668));
    ClkMux I__11230 (
            .O(N__46851),
            .I(N__46668));
    ClkMux I__11229 (
            .O(N__46850),
            .I(N__46668));
    ClkMux I__11228 (
            .O(N__46849),
            .I(N__46668));
    ClkMux I__11227 (
            .O(N__46848),
            .I(N__46668));
    ClkMux I__11226 (
            .O(N__46847),
            .I(N__46668));
    ClkMux I__11225 (
            .O(N__46846),
            .I(N__46668));
    ClkMux I__11224 (
            .O(N__46845),
            .I(N__46668));
    ClkMux I__11223 (
            .O(N__46844),
            .I(N__46668));
    ClkMux I__11222 (
            .O(N__46843),
            .I(N__46668));
    ClkMux I__11221 (
            .O(N__46842),
            .I(N__46668));
    ClkMux I__11220 (
            .O(N__46841),
            .I(N__46668));
    ClkMux I__11219 (
            .O(N__46840),
            .I(N__46668));
    ClkMux I__11218 (
            .O(N__46839),
            .I(N__46668));
    GlobalMux I__11217 (
            .O(N__46668),
            .I(N__46665));
    gio2CtrlBuf I__11216 (
            .O(N__46665),
            .I(CLK_c));
    InMux I__11215 (
            .O(N__46662),
            .I(N__46659));
    LocalMux I__11214 (
            .O(N__46659),
            .I(pin_in_22));
    InMux I__11213 (
            .O(N__46656),
            .I(N__46653));
    LocalMux I__11212 (
            .O(N__46653),
            .I(N__46650));
    Span12Mux_h I__11211 (
            .O(N__46650),
            .I(N__46647));
    Odrv12 I__11210 (
            .O(N__46647),
            .I(n13352));
    InMux I__11209 (
            .O(N__46644),
            .I(N__46641));
    LocalMux I__11208 (
            .O(N__46641),
            .I(N__46638));
    Span12Mux_h I__11207 (
            .O(N__46638),
            .I(N__46635));
    Odrv12 I__11206 (
            .O(N__46635),
            .I(pin_in_17));
    CascadeMux I__11205 (
            .O(N__46632),
            .I(N__46629));
    InMux I__11204 (
            .O(N__46629),
            .I(N__46626));
    LocalMux I__11203 (
            .O(N__46626),
            .I(N__46623));
    Span4Mux_v I__11202 (
            .O(N__46623),
            .I(N__46620));
    Sp12to4 I__11201 (
            .O(N__46620),
            .I(N__46617));
    Span12Mux_s6_h I__11200 (
            .O(N__46617),
            .I(N__46614));
    Span12Mux_v I__11199 (
            .O(N__46614),
            .I(N__46611));
    Span12Mux_v I__11198 (
            .O(N__46611),
            .I(N__46608));
    Odrv12 I__11197 (
            .O(N__46608),
            .I(pin_in_16));
    InMux I__11196 (
            .O(N__46605),
            .I(N__46602));
    LocalMux I__11195 (
            .O(N__46602),
            .I(N__46599));
    Span12Mux_h I__11194 (
            .O(N__46599),
            .I(N__46596));
    Odrv12 I__11193 (
            .O(N__46596),
            .I(n13610));
    InMux I__11192 (
            .O(N__46593),
            .I(N__46590));
    LocalMux I__11191 (
            .O(N__46590),
            .I(pin_in_19));
    CascadeMux I__11190 (
            .O(N__46587),
            .I(N__46584));
    InMux I__11189 (
            .O(N__46584),
            .I(N__46581));
    LocalMux I__11188 (
            .O(N__46581),
            .I(N__46578));
    Span4Mux_h I__11187 (
            .O(N__46578),
            .I(N__46575));
    Odrv4 I__11186 (
            .O(N__46575),
            .I(pin_in_18));
    InMux I__11185 (
            .O(N__46572),
            .I(N__46568));
    InMux I__11184 (
            .O(N__46571),
            .I(N__46560));
    LocalMux I__11183 (
            .O(N__46568),
            .I(N__46556));
    InMux I__11182 (
            .O(N__46567),
            .I(N__46552));
    InMux I__11181 (
            .O(N__46566),
            .I(N__46549));
    InMux I__11180 (
            .O(N__46565),
            .I(N__46546));
    InMux I__11179 (
            .O(N__46564),
            .I(N__46542));
    InMux I__11178 (
            .O(N__46563),
            .I(N__46539));
    LocalMux I__11177 (
            .O(N__46560),
            .I(N__46536));
    InMux I__11176 (
            .O(N__46559),
            .I(N__46533));
    Span4Mux_s2_v I__11175 (
            .O(N__46556),
            .I(N__46530));
    InMux I__11174 (
            .O(N__46555),
            .I(N__46527));
    LocalMux I__11173 (
            .O(N__46552),
            .I(N__46524));
    LocalMux I__11172 (
            .O(N__46549),
            .I(N__46517));
    LocalMux I__11171 (
            .O(N__46546),
            .I(N__46517));
    InMux I__11170 (
            .O(N__46545),
            .I(N__46514));
    LocalMux I__11169 (
            .O(N__46542),
            .I(N__46505));
    LocalMux I__11168 (
            .O(N__46539),
            .I(N__46498));
    Span4Mux_v I__11167 (
            .O(N__46536),
            .I(N__46498));
    LocalMux I__11166 (
            .O(N__46533),
            .I(N__46498));
    Sp12to4 I__11165 (
            .O(N__46530),
            .I(N__46491));
    LocalMux I__11164 (
            .O(N__46527),
            .I(N__46491));
    Span12Mux_s3_v I__11163 (
            .O(N__46524),
            .I(N__46491));
    InMux I__11162 (
            .O(N__46523),
            .I(N__46486));
    InMux I__11161 (
            .O(N__46522),
            .I(N__46486));
    Span12Mux_v I__11160 (
            .O(N__46517),
            .I(N__46481));
    LocalMux I__11159 (
            .O(N__46514),
            .I(N__46481));
    InMux I__11158 (
            .O(N__46513),
            .I(N__46478));
    InMux I__11157 (
            .O(N__46512),
            .I(N__46473));
    InMux I__11156 (
            .O(N__46511),
            .I(N__46473));
    InMux I__11155 (
            .O(N__46510),
            .I(N__46470));
    InMux I__11154 (
            .O(N__46509),
            .I(N__46467));
    InMux I__11153 (
            .O(N__46508),
            .I(N__46464));
    Span4Mux_v I__11152 (
            .O(N__46505),
            .I(N__46459));
    Span4Mux_v I__11151 (
            .O(N__46498),
            .I(N__46459));
    Span12Mux_v I__11150 (
            .O(N__46491),
            .I(N__46454));
    LocalMux I__11149 (
            .O(N__46486),
            .I(N__46454));
    Span12Mux_h I__11148 (
            .O(N__46481),
            .I(N__46451));
    LocalMux I__11147 (
            .O(N__46478),
            .I(N__46448));
    LocalMux I__11146 (
            .O(N__46473),
            .I(N__46445));
    LocalMux I__11145 (
            .O(N__46470),
            .I(current_pin_1));
    LocalMux I__11144 (
            .O(N__46467),
            .I(current_pin_1));
    LocalMux I__11143 (
            .O(N__46464),
            .I(current_pin_1));
    Odrv4 I__11142 (
            .O(N__46459),
            .I(current_pin_1));
    Odrv12 I__11141 (
            .O(N__46454),
            .I(current_pin_1));
    Odrv12 I__11140 (
            .O(N__46451),
            .I(current_pin_1));
    Odrv4 I__11139 (
            .O(N__46448),
            .I(current_pin_1));
    Odrv4 I__11138 (
            .O(N__46445),
            .I(current_pin_1));
    InMux I__11137 (
            .O(N__46428),
            .I(N__46425));
    LocalMux I__11136 (
            .O(N__46425),
            .I(N__46422));
    Odrv12 I__11135 (
            .O(N__46422),
            .I(n13607));
    CascadeMux I__11134 (
            .O(N__46419),
            .I(N__46416));
    InMux I__11133 (
            .O(N__46416),
            .I(N__46413));
    LocalMux I__11132 (
            .O(N__46413),
            .I(N__46402));
    InMux I__11131 (
            .O(N__46412),
            .I(N__46397));
    InMux I__11130 (
            .O(N__46411),
            .I(N__46397));
    InMux I__11129 (
            .O(N__46410),
            .I(N__46393));
    InMux I__11128 (
            .O(N__46409),
            .I(N__46387));
    InMux I__11127 (
            .O(N__46408),
            .I(N__46387));
    InMux I__11126 (
            .O(N__46407),
            .I(N__46378));
    InMux I__11125 (
            .O(N__46406),
            .I(N__46378));
    InMux I__11124 (
            .O(N__46405),
            .I(N__46375));
    Span4Mux_s3_v I__11123 (
            .O(N__46402),
            .I(N__46372));
    LocalMux I__11122 (
            .O(N__46397),
            .I(N__46369));
    InMux I__11121 (
            .O(N__46396),
            .I(N__46366));
    LocalMux I__11120 (
            .O(N__46393),
            .I(N__46363));
    InMux I__11119 (
            .O(N__46392),
            .I(N__46360));
    LocalMux I__11118 (
            .O(N__46387),
            .I(N__46357));
    InMux I__11117 (
            .O(N__46386),
            .I(N__46352));
    InMux I__11116 (
            .O(N__46385),
            .I(N__46352));
    InMux I__11115 (
            .O(N__46384),
            .I(N__46349));
    InMux I__11114 (
            .O(N__46383),
            .I(N__46346));
    LocalMux I__11113 (
            .O(N__46378),
            .I(N__46338));
    LocalMux I__11112 (
            .O(N__46375),
            .I(N__46338));
    Sp12to4 I__11111 (
            .O(N__46372),
            .I(N__46332));
    Sp12to4 I__11110 (
            .O(N__46369),
            .I(N__46329));
    LocalMux I__11109 (
            .O(N__46366),
            .I(N__46324));
    Span4Mux_v I__11108 (
            .O(N__46363),
            .I(N__46324));
    LocalMux I__11107 (
            .O(N__46360),
            .I(N__46315));
    Span4Mux_v I__11106 (
            .O(N__46357),
            .I(N__46315));
    LocalMux I__11105 (
            .O(N__46352),
            .I(N__46308));
    LocalMux I__11104 (
            .O(N__46349),
            .I(N__46308));
    LocalMux I__11103 (
            .O(N__46346),
            .I(N__46308));
    InMux I__11102 (
            .O(N__46345),
            .I(N__46303));
    InMux I__11101 (
            .O(N__46344),
            .I(N__46303));
    InMux I__11100 (
            .O(N__46343),
            .I(N__46300));
    Span12Mux_v I__11099 (
            .O(N__46338),
            .I(N__46297));
    InMux I__11098 (
            .O(N__46337),
            .I(N__46294));
    InMux I__11097 (
            .O(N__46336),
            .I(N__46289));
    InMux I__11096 (
            .O(N__46335),
            .I(N__46289));
    Span12Mux_h I__11095 (
            .O(N__46332),
            .I(N__46284));
    Span12Mux_s3_v I__11094 (
            .O(N__46329),
            .I(N__46284));
    Sp12to4 I__11093 (
            .O(N__46324),
            .I(N__46281));
    InMux I__11092 (
            .O(N__46323),
            .I(N__46278));
    InMux I__11091 (
            .O(N__46322),
            .I(N__46275));
    InMux I__11090 (
            .O(N__46321),
            .I(N__46272));
    InMux I__11089 (
            .O(N__46320),
            .I(N__46269));
    Span4Mux_v I__11088 (
            .O(N__46315),
            .I(N__46264));
    Span4Mux_v I__11087 (
            .O(N__46308),
            .I(N__46264));
    LocalMux I__11086 (
            .O(N__46303),
            .I(N__46257));
    LocalMux I__11085 (
            .O(N__46300),
            .I(N__46257));
    Span12Mux_h I__11084 (
            .O(N__46297),
            .I(N__46257));
    LocalMux I__11083 (
            .O(N__46294),
            .I(N__46248));
    LocalMux I__11082 (
            .O(N__46289),
            .I(N__46248));
    Span12Mux_v I__11081 (
            .O(N__46284),
            .I(N__46248));
    Span12Mux_h I__11080 (
            .O(N__46281),
            .I(N__46248));
    LocalMux I__11079 (
            .O(N__46278),
            .I(current_pin_0));
    LocalMux I__11078 (
            .O(N__46275),
            .I(current_pin_0));
    LocalMux I__11077 (
            .O(N__46272),
            .I(current_pin_0));
    LocalMux I__11076 (
            .O(N__46269),
            .I(current_pin_0));
    Odrv4 I__11075 (
            .O(N__46264),
            .I(current_pin_0));
    Odrv12 I__11074 (
            .O(N__46257),
            .I(current_pin_0));
    Odrv12 I__11073 (
            .O(N__46248),
            .I(current_pin_0));
    InMux I__11072 (
            .O(N__46233),
            .I(N__46230));
    LocalMux I__11071 (
            .O(N__46230),
            .I(pin_in_21));
    InMux I__11070 (
            .O(N__46227),
            .I(N__46224));
    LocalMux I__11069 (
            .O(N__46224),
            .I(N__46221));
    Span4Mux_h I__11068 (
            .O(N__46221),
            .I(N__46218));
    Odrv4 I__11067 (
            .O(N__46218),
            .I(pin_in_20));
    InMux I__11066 (
            .O(N__46215),
            .I(N__46212));
    LocalMux I__11065 (
            .O(N__46212),
            .I(n19_adj_789));
    CascadeMux I__11064 (
            .O(N__46209),
            .I(n13375_cascade_));
    InMux I__11063 (
            .O(N__46206),
            .I(N__46203));
    LocalMux I__11062 (
            .O(N__46203),
            .I(N__46200));
    Span4Mux_h I__11061 (
            .O(N__46200),
            .I(N__46197));
    Odrv4 I__11060 (
            .O(N__46197),
            .I(n13637));
    InMux I__11059 (
            .O(N__46194),
            .I(N__46191));
    LocalMux I__11058 (
            .O(N__46191),
            .I(N__46188));
    Odrv4 I__11057 (
            .O(N__46188),
            .I(n8_adj_829));
    IoInMux I__11056 (
            .O(N__46185),
            .I(N__46182));
    LocalMux I__11055 (
            .O(N__46182),
            .I(N__46179));
    IoSpan4Mux I__11054 (
            .O(N__46179),
            .I(N__46176));
    Span4Mux_s2_v I__11053 (
            .O(N__46176),
            .I(N__46173));
    Sp12to4 I__11052 (
            .O(N__46173),
            .I(N__46170));
    Span12Mux_h I__11051 (
            .O(N__46170),
            .I(N__46167));
    Span12Mux_v I__11050 (
            .O(N__46167),
            .I(N__46162));
    InMux I__11049 (
            .O(N__46166),
            .I(N__46157));
    InMux I__11048 (
            .O(N__46165),
            .I(N__46157));
    Odrv12 I__11047 (
            .O(N__46162),
            .I(pin_out_12));
    LocalMux I__11046 (
            .O(N__46157),
            .I(pin_out_12));
    CascadeMux I__11045 (
            .O(N__46152),
            .I(N__46148));
    CascadeMux I__11044 (
            .O(N__46151),
            .I(N__46133));
    InMux I__11043 (
            .O(N__46148),
            .I(N__46129));
    InMux I__11042 (
            .O(N__46147),
            .I(N__46126));
    InMux I__11041 (
            .O(N__46146),
            .I(N__46121));
    InMux I__11040 (
            .O(N__46145),
            .I(N__46121));
    InMux I__11039 (
            .O(N__46144),
            .I(N__46118));
    InMux I__11038 (
            .O(N__46143),
            .I(N__46115));
    InMux I__11037 (
            .O(N__46142),
            .I(N__46112));
    InMux I__11036 (
            .O(N__46141),
            .I(N__46107));
    InMux I__11035 (
            .O(N__46140),
            .I(N__46104));
    InMux I__11034 (
            .O(N__46139),
            .I(N__46099));
    InMux I__11033 (
            .O(N__46138),
            .I(N__46099));
    InMux I__11032 (
            .O(N__46137),
            .I(N__46089));
    InMux I__11031 (
            .O(N__46136),
            .I(N__46089));
    InMux I__11030 (
            .O(N__46133),
            .I(N__46086));
    InMux I__11029 (
            .O(N__46132),
            .I(N__46083));
    LocalMux I__11028 (
            .O(N__46129),
            .I(N__46080));
    LocalMux I__11027 (
            .O(N__46126),
            .I(N__46077));
    LocalMux I__11026 (
            .O(N__46121),
            .I(N__46074));
    LocalMux I__11025 (
            .O(N__46118),
            .I(N__46067));
    LocalMux I__11024 (
            .O(N__46115),
            .I(N__46067));
    LocalMux I__11023 (
            .O(N__46112),
            .I(N__46067));
    InMux I__11022 (
            .O(N__46111),
            .I(N__46064));
    InMux I__11021 (
            .O(N__46110),
            .I(N__46061));
    LocalMux I__11020 (
            .O(N__46107),
            .I(N__46054));
    LocalMux I__11019 (
            .O(N__46104),
            .I(N__46054));
    LocalMux I__11018 (
            .O(N__46099),
            .I(N__46054));
    InMux I__11017 (
            .O(N__46098),
            .I(N__46049));
    InMux I__11016 (
            .O(N__46097),
            .I(N__46049));
    InMux I__11015 (
            .O(N__46096),
            .I(N__46046));
    InMux I__11014 (
            .O(N__46095),
            .I(N__46041));
    InMux I__11013 (
            .O(N__46094),
            .I(N__46041));
    LocalMux I__11012 (
            .O(N__46089),
            .I(N__46026));
    LocalMux I__11011 (
            .O(N__46086),
            .I(N__46026));
    LocalMux I__11010 (
            .O(N__46083),
            .I(N__46026));
    Span4Mux_v I__11009 (
            .O(N__46080),
            .I(N__46026));
    Span4Mux_h I__11008 (
            .O(N__46077),
            .I(N__46026));
    Span4Mux_h I__11007 (
            .O(N__46074),
            .I(N__46026));
    Span4Mux_v I__11006 (
            .O(N__46067),
            .I(N__46026));
    LocalMux I__11005 (
            .O(N__46064),
            .I(N__46019));
    LocalMux I__11004 (
            .O(N__46061),
            .I(N__46019));
    Span4Mux_v I__11003 (
            .O(N__46054),
            .I(N__46019));
    LocalMux I__11002 (
            .O(N__46049),
            .I(n9675));
    LocalMux I__11001 (
            .O(N__46046),
            .I(n9675));
    LocalMux I__11000 (
            .O(N__46041),
            .I(n9675));
    Odrv4 I__10999 (
            .O(N__46026),
            .I(n9675));
    Odrv4 I__10998 (
            .O(N__46019),
            .I(n9675));
    InMux I__10997 (
            .O(N__46008),
            .I(N__46005));
    LocalMux I__10996 (
            .O(N__46005),
            .I(N__46002));
    Span4Mux_h I__10995 (
            .O(N__46002),
            .I(N__45999));
    Odrv4 I__10994 (
            .O(N__45999),
            .I(n7_adj_830));
    InMux I__10993 (
            .O(N__45996),
            .I(N__45987));
    InMux I__10992 (
            .O(N__45995),
            .I(N__45987));
    InMux I__10991 (
            .O(N__45994),
            .I(N__45982));
    InMux I__10990 (
            .O(N__45993),
            .I(N__45982));
    CascadeMux I__10989 (
            .O(N__45992),
            .I(N__45975));
    LocalMux I__10988 (
            .O(N__45987),
            .I(N__45965));
    LocalMux I__10987 (
            .O(N__45982),
            .I(N__45965));
    CEMux I__10986 (
            .O(N__45981),
            .I(N__45962));
    InMux I__10985 (
            .O(N__45980),
            .I(N__45953));
    InMux I__10984 (
            .O(N__45979),
            .I(N__45949));
    InMux I__10983 (
            .O(N__45978),
            .I(N__45944));
    InMux I__10982 (
            .O(N__45975),
            .I(N__45944));
    InMux I__10981 (
            .O(N__45974),
            .I(N__45941));
    InMux I__10980 (
            .O(N__45973),
            .I(N__45936));
    InMux I__10979 (
            .O(N__45972),
            .I(N__45936));
    InMux I__10978 (
            .O(N__45971),
            .I(N__45931));
    InMux I__10977 (
            .O(N__45970),
            .I(N__45931));
    Span4Mux_v I__10976 (
            .O(N__45965),
            .I(N__45926));
    LocalMux I__10975 (
            .O(N__45962),
            .I(N__45926));
    CEMux I__10974 (
            .O(N__45961),
            .I(N__45923));
    InMux I__10973 (
            .O(N__45960),
            .I(N__45920));
    InMux I__10972 (
            .O(N__45959),
            .I(N__45917));
    InMux I__10971 (
            .O(N__45958),
            .I(N__45912));
    InMux I__10970 (
            .O(N__45957),
            .I(N__45912));
    InMux I__10969 (
            .O(N__45956),
            .I(N__45909));
    LocalMux I__10968 (
            .O(N__45953),
            .I(N__45906));
    InMux I__10967 (
            .O(N__45952),
            .I(N__45903));
    LocalMux I__10966 (
            .O(N__45949),
            .I(N__45893));
    LocalMux I__10965 (
            .O(N__45944),
            .I(N__45893));
    LocalMux I__10964 (
            .O(N__45941),
            .I(N__45886));
    LocalMux I__10963 (
            .O(N__45936),
            .I(N__45886));
    LocalMux I__10962 (
            .O(N__45931),
            .I(N__45886));
    Span4Mux_h I__10961 (
            .O(N__45926),
            .I(N__45883));
    LocalMux I__10960 (
            .O(N__45923),
            .I(N__45880));
    LocalMux I__10959 (
            .O(N__45920),
            .I(N__45867));
    LocalMux I__10958 (
            .O(N__45917),
            .I(N__45867));
    LocalMux I__10957 (
            .O(N__45912),
            .I(N__45867));
    LocalMux I__10956 (
            .O(N__45909),
            .I(N__45867));
    Sp12to4 I__10955 (
            .O(N__45906),
            .I(N__45867));
    LocalMux I__10954 (
            .O(N__45903),
            .I(N__45867));
    InMux I__10953 (
            .O(N__45902),
            .I(N__45864));
    InMux I__10952 (
            .O(N__45901),
            .I(N__45861));
    InMux I__10951 (
            .O(N__45900),
            .I(N__45856));
    InMux I__10950 (
            .O(N__45899),
            .I(N__45856));
    InMux I__10949 (
            .O(N__45898),
            .I(N__45853));
    Span4Mux_h I__10948 (
            .O(N__45893),
            .I(N__45848));
    Span4Mux_v I__10947 (
            .O(N__45886),
            .I(N__45848));
    Span4Mux_h I__10946 (
            .O(N__45883),
            .I(N__45845));
    Span4Mux_v I__10945 (
            .O(N__45880),
            .I(N__45842));
    Span12Mux_v I__10944 (
            .O(N__45867),
            .I(N__45839));
    LocalMux I__10943 (
            .O(N__45864),
            .I(N__45836));
    LocalMux I__10942 (
            .O(N__45861),
            .I(n11789));
    LocalMux I__10941 (
            .O(N__45856),
            .I(n11789));
    LocalMux I__10940 (
            .O(N__45853),
            .I(n11789));
    Odrv4 I__10939 (
            .O(N__45848),
            .I(n11789));
    Odrv4 I__10938 (
            .O(N__45845),
            .I(n11789));
    Odrv4 I__10937 (
            .O(N__45842),
            .I(n11789));
    Odrv12 I__10936 (
            .O(N__45839),
            .I(n11789));
    Odrv4 I__10935 (
            .O(N__45836),
            .I(n11789));
    IoInMux I__10934 (
            .O(N__45819),
            .I(N__45816));
    LocalMux I__10933 (
            .O(N__45816),
            .I(N__45813));
    Span12Mux_s7_h I__10932 (
            .O(N__45813),
            .I(N__45808));
    InMux I__10931 (
            .O(N__45812),
            .I(N__45803));
    InMux I__10930 (
            .O(N__45811),
            .I(N__45803));
    Odrv12 I__10929 (
            .O(N__45808),
            .I(pin_out_13));
    LocalMux I__10928 (
            .O(N__45803),
            .I(pin_out_13));
    IoInMux I__10927 (
            .O(N__45798),
            .I(N__45795));
    LocalMux I__10926 (
            .O(N__45795),
            .I(N__45792));
    IoSpan4Mux I__10925 (
            .O(N__45792),
            .I(N__45789));
    Sp12to4 I__10924 (
            .O(N__45789),
            .I(N__45784));
    InMux I__10923 (
            .O(N__45788),
            .I(N__45781));
    InMux I__10922 (
            .O(N__45787),
            .I(N__45778));
    Span12Mux_s9_h I__10921 (
            .O(N__45784),
            .I(N__45773));
    LocalMux I__10920 (
            .O(N__45781),
            .I(N__45773));
    LocalMux I__10919 (
            .O(N__45778),
            .I(pin_out_15));
    Odrv12 I__10918 (
            .O(N__45773),
            .I(pin_out_15));
    IoInMux I__10917 (
            .O(N__45768),
            .I(N__45765));
    LocalMux I__10916 (
            .O(N__45765),
            .I(N__45762));
    IoSpan4Mux I__10915 (
            .O(N__45762),
            .I(N__45759));
    Span4Mux_s0_h I__10914 (
            .O(N__45759),
            .I(N__45756));
    Sp12to4 I__10913 (
            .O(N__45756),
            .I(N__45753));
    Span12Mux_h I__10912 (
            .O(N__45753),
            .I(N__45748));
    InMux I__10911 (
            .O(N__45752),
            .I(N__45745));
    InMux I__10910 (
            .O(N__45751),
            .I(N__45742));
    Odrv12 I__10909 (
            .O(N__45748),
            .I(pin_out_14));
    LocalMux I__10908 (
            .O(N__45745),
            .I(pin_out_14));
    LocalMux I__10907 (
            .O(N__45742),
            .I(pin_out_14));
    InMux I__10906 (
            .O(N__45735),
            .I(N__45732));
    LocalMux I__10905 (
            .O(N__45732),
            .I(n13376));
    InMux I__10904 (
            .O(N__45729),
            .I(N__45726));
    LocalMux I__10903 (
            .O(N__45726),
            .I(n11956));
    IoInMux I__10902 (
            .O(N__45723),
            .I(N__45720));
    LocalMux I__10901 (
            .O(N__45720),
            .I(N__45717));
    IoSpan4Mux I__10900 (
            .O(N__45717),
            .I(N__45714));
    Span4Mux_s1_h I__10899 (
            .O(N__45714),
            .I(N__45711));
    Span4Mux_h I__10898 (
            .O(N__45711),
            .I(N__45708));
    Span4Mux_h I__10897 (
            .O(N__45708),
            .I(N__45704));
    InMux I__10896 (
            .O(N__45707),
            .I(N__45701));
    Odrv4 I__10895 (
            .O(N__45704),
            .I(pin_oe_13));
    LocalMux I__10894 (
            .O(N__45701),
            .I(pin_oe_13));
    CascadeMux I__10893 (
            .O(N__45696),
            .I(N__45692));
    CascadeMux I__10892 (
            .O(N__45695),
            .I(N__45689));
    InMux I__10891 (
            .O(N__45692),
            .I(N__45686));
    InMux I__10890 (
            .O(N__45689),
            .I(N__45683));
    LocalMux I__10889 (
            .O(N__45686),
            .I(N__45678));
    LocalMux I__10888 (
            .O(N__45683),
            .I(N__45675));
    CascadeMux I__10887 (
            .O(N__45682),
            .I(N__45672));
    CascadeMux I__10886 (
            .O(N__45681),
            .I(N__45665));
    Span4Mux_v I__10885 (
            .O(N__45678),
            .I(N__45661));
    Span4Mux_v I__10884 (
            .O(N__45675),
            .I(N__45658));
    InMux I__10883 (
            .O(N__45672),
            .I(N__45655));
    InMux I__10882 (
            .O(N__45671),
            .I(N__45646));
    CascadeMux I__10881 (
            .O(N__45670),
            .I(N__45638));
    CascadeMux I__10880 (
            .O(N__45669),
            .I(N__45635));
    InMux I__10879 (
            .O(N__45668),
            .I(N__45631));
    InMux I__10878 (
            .O(N__45665),
            .I(N__45628));
    CascadeMux I__10877 (
            .O(N__45664),
            .I(N__45624));
    Span4Mux_h I__10876 (
            .O(N__45661),
            .I(N__45619));
    Span4Mux_h I__10875 (
            .O(N__45658),
            .I(N__45619));
    LocalMux I__10874 (
            .O(N__45655),
            .I(N__45616));
    CascadeMux I__10873 (
            .O(N__45654),
            .I(N__45612));
    CascadeMux I__10872 (
            .O(N__45653),
            .I(N__45608));
    CascadeMux I__10871 (
            .O(N__45652),
            .I(N__45605));
    CascadeMux I__10870 (
            .O(N__45651),
            .I(N__45602));
    CascadeMux I__10869 (
            .O(N__45650),
            .I(N__45599));
    CascadeMux I__10868 (
            .O(N__45649),
            .I(N__45593));
    LocalMux I__10867 (
            .O(N__45646),
            .I(N__45589));
    InMux I__10866 (
            .O(N__45645),
            .I(N__45584));
    InMux I__10865 (
            .O(N__45644),
            .I(N__45581));
    CascadeMux I__10864 (
            .O(N__45643),
            .I(N__45578));
    CascadeMux I__10863 (
            .O(N__45642),
            .I(N__45575));
    CascadeMux I__10862 (
            .O(N__45641),
            .I(N__45571));
    InMux I__10861 (
            .O(N__45638),
            .I(N__45564));
    InMux I__10860 (
            .O(N__45635),
            .I(N__45561));
    CascadeMux I__10859 (
            .O(N__45634),
            .I(N__45557));
    LocalMux I__10858 (
            .O(N__45631),
            .I(N__45553));
    LocalMux I__10857 (
            .O(N__45628),
            .I(N__45550));
    InMux I__10856 (
            .O(N__45627),
            .I(N__45547));
    InMux I__10855 (
            .O(N__45624),
            .I(N__45544));
    Span4Mux_v I__10854 (
            .O(N__45619),
            .I(N__45539));
    Span4Mux_v I__10853 (
            .O(N__45616),
            .I(N__45539));
    CascadeMux I__10852 (
            .O(N__45615),
            .I(N__45535));
    InMux I__10851 (
            .O(N__45612),
            .I(N__45531));
    InMux I__10850 (
            .O(N__45611),
            .I(N__45526));
    InMux I__10849 (
            .O(N__45608),
            .I(N__45526));
    InMux I__10848 (
            .O(N__45605),
            .I(N__45523));
    InMux I__10847 (
            .O(N__45602),
            .I(N__45520));
    InMux I__10846 (
            .O(N__45599),
            .I(N__45515));
    InMux I__10845 (
            .O(N__45598),
            .I(N__45515));
    CascadeMux I__10844 (
            .O(N__45597),
            .I(N__45512));
    CascadeMux I__10843 (
            .O(N__45596),
            .I(N__45509));
    InMux I__10842 (
            .O(N__45593),
            .I(N__45502));
    InMux I__10841 (
            .O(N__45592),
            .I(N__45502));
    Span4Mux_h I__10840 (
            .O(N__45589),
            .I(N__45499));
    CascadeMux I__10839 (
            .O(N__45588),
            .I(N__45494));
    CascadeMux I__10838 (
            .O(N__45587),
            .I(N__45489));
    LocalMux I__10837 (
            .O(N__45584),
            .I(N__45482));
    LocalMux I__10836 (
            .O(N__45581),
            .I(N__45482));
    InMux I__10835 (
            .O(N__45578),
            .I(N__45478));
    InMux I__10834 (
            .O(N__45575),
            .I(N__45475));
    InMux I__10833 (
            .O(N__45574),
            .I(N__45472));
    InMux I__10832 (
            .O(N__45571),
            .I(N__45467));
    InMux I__10831 (
            .O(N__45570),
            .I(N__45467));
    CascadeMux I__10830 (
            .O(N__45569),
            .I(N__45463));
    CascadeMux I__10829 (
            .O(N__45568),
            .I(N__45458));
    CascadeMux I__10828 (
            .O(N__45567),
            .I(N__45455));
    LocalMux I__10827 (
            .O(N__45564),
            .I(N__45449));
    LocalMux I__10826 (
            .O(N__45561),
            .I(N__45446));
    InMux I__10825 (
            .O(N__45560),
            .I(N__45443));
    InMux I__10824 (
            .O(N__45557),
            .I(N__45438));
    InMux I__10823 (
            .O(N__45556),
            .I(N__45438));
    Span4Mux_h I__10822 (
            .O(N__45553),
            .I(N__45431));
    Span4Mux_v I__10821 (
            .O(N__45550),
            .I(N__45431));
    LocalMux I__10820 (
            .O(N__45547),
            .I(N__45431));
    LocalMux I__10819 (
            .O(N__45544),
            .I(N__45426));
    Span4Mux_h I__10818 (
            .O(N__45539),
            .I(N__45426));
    InMux I__10817 (
            .O(N__45538),
            .I(N__45419));
    InMux I__10816 (
            .O(N__45535),
            .I(N__45419));
    InMux I__10815 (
            .O(N__45534),
            .I(N__45419));
    LocalMux I__10814 (
            .O(N__45531),
            .I(N__45408));
    LocalMux I__10813 (
            .O(N__45526),
            .I(N__45408));
    LocalMux I__10812 (
            .O(N__45523),
            .I(N__45408));
    LocalMux I__10811 (
            .O(N__45520),
            .I(N__45408));
    LocalMux I__10810 (
            .O(N__45515),
            .I(N__45408));
    InMux I__10809 (
            .O(N__45512),
            .I(N__45403));
    InMux I__10808 (
            .O(N__45509),
            .I(N__45403));
    InMux I__10807 (
            .O(N__45508),
            .I(N__45398));
    InMux I__10806 (
            .O(N__45507),
            .I(N__45398));
    LocalMux I__10805 (
            .O(N__45502),
            .I(N__45393));
    Span4Mux_h I__10804 (
            .O(N__45499),
            .I(N__45393));
    InMux I__10803 (
            .O(N__45498),
            .I(N__45388));
    InMux I__10802 (
            .O(N__45497),
            .I(N__45388));
    InMux I__10801 (
            .O(N__45494),
            .I(N__45383));
    InMux I__10800 (
            .O(N__45493),
            .I(N__45383));
    InMux I__10799 (
            .O(N__45492),
            .I(N__45380));
    InMux I__10798 (
            .O(N__45489),
            .I(N__45377));
    InMux I__10797 (
            .O(N__45488),
            .I(N__45372));
    InMux I__10796 (
            .O(N__45487),
            .I(N__45372));
    Span12Mux_v I__10795 (
            .O(N__45482),
            .I(N__45369));
    InMux I__10794 (
            .O(N__45481),
            .I(N__45366));
    LocalMux I__10793 (
            .O(N__45478),
            .I(N__45361));
    LocalMux I__10792 (
            .O(N__45475),
            .I(N__45361));
    LocalMux I__10791 (
            .O(N__45472),
            .I(N__45356));
    LocalMux I__10790 (
            .O(N__45467),
            .I(N__45356));
    InMux I__10789 (
            .O(N__45466),
            .I(N__45351));
    InMux I__10788 (
            .O(N__45463),
            .I(N__45351));
    InMux I__10787 (
            .O(N__45462),
            .I(N__45348));
    InMux I__10786 (
            .O(N__45461),
            .I(N__45345));
    InMux I__10785 (
            .O(N__45458),
            .I(N__45338));
    InMux I__10784 (
            .O(N__45455),
            .I(N__45338));
    InMux I__10783 (
            .O(N__45454),
            .I(N__45338));
    InMux I__10782 (
            .O(N__45453),
            .I(N__45333));
    InMux I__10781 (
            .O(N__45452),
            .I(N__45333));
    Span4Mux_v I__10780 (
            .O(N__45449),
            .I(N__45316));
    Span4Mux_v I__10779 (
            .O(N__45446),
            .I(N__45316));
    LocalMux I__10778 (
            .O(N__45443),
            .I(N__45316));
    LocalMux I__10777 (
            .O(N__45438),
            .I(N__45316));
    Span4Mux_v I__10776 (
            .O(N__45431),
            .I(N__45316));
    Span4Mux_h I__10775 (
            .O(N__45426),
            .I(N__45316));
    LocalMux I__10774 (
            .O(N__45419),
            .I(N__45316));
    Span4Mux_v I__10773 (
            .O(N__45408),
            .I(N__45316));
    LocalMux I__10772 (
            .O(N__45403),
            .I(N__45305));
    LocalMux I__10771 (
            .O(N__45398),
            .I(N__45305));
    Span4Mux_h I__10770 (
            .O(N__45393),
            .I(N__45305));
    LocalMux I__10769 (
            .O(N__45388),
            .I(N__45305));
    LocalMux I__10768 (
            .O(N__45383),
            .I(N__45305));
    LocalMux I__10767 (
            .O(N__45380),
            .I(N__45302));
    LocalMux I__10766 (
            .O(N__45377),
            .I(N__45295));
    LocalMux I__10765 (
            .O(N__45372),
            .I(N__45295));
    Span12Mux_h I__10764 (
            .O(N__45369),
            .I(N__45295));
    LocalMux I__10763 (
            .O(N__45366),
            .I(current_pin_2));
    Odrv4 I__10762 (
            .O(N__45361),
            .I(current_pin_2));
    Odrv4 I__10761 (
            .O(N__45356),
            .I(current_pin_2));
    LocalMux I__10760 (
            .O(N__45351),
            .I(current_pin_2));
    LocalMux I__10759 (
            .O(N__45348),
            .I(current_pin_2));
    LocalMux I__10758 (
            .O(N__45345),
            .I(current_pin_2));
    LocalMux I__10757 (
            .O(N__45338),
            .I(current_pin_2));
    LocalMux I__10756 (
            .O(N__45333),
            .I(current_pin_2));
    Odrv4 I__10755 (
            .O(N__45316),
            .I(current_pin_2));
    Odrv4 I__10754 (
            .O(N__45305),
            .I(current_pin_2));
    Odrv4 I__10753 (
            .O(N__45302),
            .I(current_pin_2));
    Odrv12 I__10752 (
            .O(N__45295),
            .I(current_pin_2));
    CascadeMux I__10751 (
            .O(N__45270),
            .I(N__45264));
    InMux I__10750 (
            .O(N__45269),
            .I(N__45258));
    InMux I__10749 (
            .O(N__45268),
            .I(N__45255));
    InMux I__10748 (
            .O(N__45267),
            .I(N__45247));
    InMux I__10747 (
            .O(N__45264),
            .I(N__45240));
    InMux I__10746 (
            .O(N__45263),
            .I(N__45240));
    InMux I__10745 (
            .O(N__45262),
            .I(N__45240));
    InMux I__10744 (
            .O(N__45261),
            .I(N__45237));
    LocalMux I__10743 (
            .O(N__45258),
            .I(N__45234));
    LocalMux I__10742 (
            .O(N__45255),
            .I(N__45231));
    InMux I__10741 (
            .O(N__45254),
            .I(N__45226));
    InMux I__10740 (
            .O(N__45253),
            .I(N__45226));
    InMux I__10739 (
            .O(N__45252),
            .I(N__45219));
    InMux I__10738 (
            .O(N__45251),
            .I(N__45219));
    InMux I__10737 (
            .O(N__45250),
            .I(N__45219));
    LocalMux I__10736 (
            .O(N__45247),
            .I(N__45210));
    LocalMux I__10735 (
            .O(N__45240),
            .I(N__45210));
    LocalMux I__10734 (
            .O(N__45237),
            .I(N__45210));
    Span4Mux_v I__10733 (
            .O(N__45234),
            .I(N__45210));
    Odrv4 I__10732 (
            .O(N__45231),
            .I(current_pin_3));
    LocalMux I__10731 (
            .O(N__45226),
            .I(current_pin_3));
    LocalMux I__10730 (
            .O(N__45219),
            .I(current_pin_3));
    Odrv4 I__10729 (
            .O(N__45210),
            .I(current_pin_3));
    InMux I__10728 (
            .O(N__45201),
            .I(N__45198));
    LocalMux I__10727 (
            .O(N__45198),
            .I(N__45195));
    Span4Mux_h I__10726 (
            .O(N__45195),
            .I(N__45192));
    Odrv4 I__10725 (
            .O(N__45192),
            .I(n13465));
    InMux I__10724 (
            .O(N__45189),
            .I(N__45186));
    LocalMux I__10723 (
            .O(N__45186),
            .I(N__45183));
    Sp12to4 I__10722 (
            .O(N__45183),
            .I(N__45180));
    Span12Mux_v I__10721 (
            .O(N__45180),
            .I(N__45177));
    Odrv12 I__10720 (
            .O(N__45177),
            .I(pin_in_15));
    CascadeMux I__10719 (
            .O(N__45174),
            .I(N__45171));
    InMux I__10718 (
            .O(N__45171),
            .I(N__45168));
    LocalMux I__10717 (
            .O(N__45168),
            .I(N__45165));
    Span4Mux_v I__10716 (
            .O(N__45165),
            .I(N__45162));
    Sp12to4 I__10715 (
            .O(N__45162),
            .I(N__45159));
    Span12Mux_h I__10714 (
            .O(N__45159),
            .I(N__45156));
    Span12Mux_v I__10713 (
            .O(N__45156),
            .I(N__45153));
    Odrv12 I__10712 (
            .O(N__45153),
            .I(pin_in_14));
    InMux I__10711 (
            .O(N__45150),
            .I(N__45147));
    LocalMux I__10710 (
            .O(N__45147),
            .I(N__45144));
    Span12Mux_h I__10709 (
            .O(N__45144),
            .I(N__45141));
    Odrv12 I__10708 (
            .O(N__45141),
            .I(pin_in_13));
    CascadeMux I__10707 (
            .O(N__45138),
            .I(n13643_cascade_));
    InMux I__10706 (
            .O(N__45135),
            .I(N__45132));
    LocalMux I__10705 (
            .O(N__45132),
            .I(N__45129));
    Span4Mux_v I__10704 (
            .O(N__45129),
            .I(N__45126));
    Sp12to4 I__10703 (
            .O(N__45126),
            .I(N__45123));
    Span12Mux_v I__10702 (
            .O(N__45123),
            .I(N__45120));
    Odrv12 I__10701 (
            .O(N__45120),
            .I(pin_in_12));
    InMux I__10700 (
            .O(N__45117),
            .I(N__45114));
    LocalMux I__10699 (
            .O(N__45114),
            .I(N__45111));
    Odrv12 I__10698 (
            .O(N__45111),
            .I(n13646));
    InMux I__10697 (
            .O(N__45108),
            .I(N__45102));
    InMux I__10696 (
            .O(N__45107),
            .I(N__45095));
    InMux I__10695 (
            .O(N__45106),
            .I(N__45092));
    InMux I__10694 (
            .O(N__45105),
            .I(N__45086));
    LocalMux I__10693 (
            .O(N__45102),
            .I(N__45083));
    InMux I__10692 (
            .O(N__45101),
            .I(N__45080));
    InMux I__10691 (
            .O(N__45100),
            .I(N__45077));
    InMux I__10690 (
            .O(N__45099),
            .I(N__45072));
    InMux I__10689 (
            .O(N__45098),
            .I(N__45072));
    LocalMux I__10688 (
            .O(N__45095),
            .I(N__45069));
    LocalMux I__10687 (
            .O(N__45092),
            .I(N__45066));
    InMux I__10686 (
            .O(N__45091),
            .I(N__45063));
    InMux I__10685 (
            .O(N__45090),
            .I(N__45059));
    InMux I__10684 (
            .O(N__45089),
            .I(N__45056));
    LocalMux I__10683 (
            .O(N__45086),
            .I(N__45053));
    Span4Mux_h I__10682 (
            .O(N__45083),
            .I(N__45046));
    LocalMux I__10681 (
            .O(N__45080),
            .I(N__45046));
    LocalMux I__10680 (
            .O(N__45077),
            .I(N__45046));
    LocalMux I__10679 (
            .O(N__45072),
            .I(N__45037));
    Span4Mux_h I__10678 (
            .O(N__45069),
            .I(N__45037));
    Span4Mux_h I__10677 (
            .O(N__45066),
            .I(N__45037));
    LocalMux I__10676 (
            .O(N__45063),
            .I(N__45037));
    InMux I__10675 (
            .O(N__45062),
            .I(N__45034));
    LocalMux I__10674 (
            .O(N__45059),
            .I(n7_adj_797));
    LocalMux I__10673 (
            .O(N__45056),
            .I(n7_adj_797));
    Odrv4 I__10672 (
            .O(N__45053),
            .I(n7_adj_797));
    Odrv4 I__10671 (
            .O(N__45046),
            .I(n7_adj_797));
    Odrv4 I__10670 (
            .O(N__45037),
            .I(n7_adj_797));
    LocalMux I__10669 (
            .O(N__45034),
            .I(n7_adj_797));
    InMux I__10668 (
            .O(N__45021),
            .I(N__45014));
    InMux I__10667 (
            .O(N__45020),
            .I(N__45014));
    InMux I__10666 (
            .O(N__45019),
            .I(N__45011));
    LocalMux I__10665 (
            .O(N__45014),
            .I(N__45007));
    LocalMux I__10664 (
            .O(N__45011),
            .I(N__45003));
    InMux I__10663 (
            .O(N__45010),
            .I(N__45000));
    Span4Mux_v I__10662 (
            .O(N__45007),
            .I(N__44997));
    InMux I__10661 (
            .O(N__45006),
            .I(N__44992));
    Span4Mux_v I__10660 (
            .O(N__45003),
            .I(N__44985));
    LocalMux I__10659 (
            .O(N__45000),
            .I(N__44985));
    Span4Mux_h I__10658 (
            .O(N__44997),
            .I(N__44982));
    CascadeMux I__10657 (
            .O(N__44996),
            .I(N__44978));
    InMux I__10656 (
            .O(N__44995),
            .I(N__44975));
    LocalMux I__10655 (
            .O(N__44992),
            .I(N__44972));
    InMux I__10654 (
            .O(N__44991),
            .I(N__44969));
    InMux I__10653 (
            .O(N__44990),
            .I(N__44965));
    Span4Mux_h I__10652 (
            .O(N__44985),
            .I(N__44959));
    Span4Mux_h I__10651 (
            .O(N__44982),
            .I(N__44959));
    InMux I__10650 (
            .O(N__44981),
            .I(N__44956));
    InMux I__10649 (
            .O(N__44978),
            .I(N__44953));
    LocalMux I__10648 (
            .O(N__44975),
            .I(N__44946));
    Span4Mux_h I__10647 (
            .O(N__44972),
            .I(N__44946));
    LocalMux I__10646 (
            .O(N__44969),
            .I(N__44946));
    InMux I__10645 (
            .O(N__44968),
            .I(N__44943));
    LocalMux I__10644 (
            .O(N__44965),
            .I(N__44940));
    InMux I__10643 (
            .O(N__44964),
            .I(N__44937));
    Span4Mux_h I__10642 (
            .O(N__44959),
            .I(N__44934));
    LocalMux I__10641 (
            .O(N__44956),
            .I(N__44929));
    LocalMux I__10640 (
            .O(N__44953),
            .I(N__44929));
    Span4Mux_v I__10639 (
            .O(N__44946),
            .I(N__44926));
    LocalMux I__10638 (
            .O(N__44943),
            .I(n6));
    Odrv4 I__10637 (
            .O(N__44940),
            .I(n6));
    LocalMux I__10636 (
            .O(N__44937),
            .I(n6));
    Odrv4 I__10635 (
            .O(N__44934),
            .I(n6));
    Odrv12 I__10634 (
            .O(N__44929),
            .I(n6));
    Odrv4 I__10633 (
            .O(N__44926),
            .I(n6));
    CascadeMux I__10632 (
            .O(N__44913),
            .I(N__44904));
    CascadeMux I__10631 (
            .O(N__44912),
            .I(N__44899));
    InMux I__10630 (
            .O(N__44911),
            .I(N__44896));
    CascadeMux I__10629 (
            .O(N__44910),
            .I(N__44893));
    CascadeMux I__10628 (
            .O(N__44909),
            .I(N__44887));
    InMux I__10627 (
            .O(N__44908),
            .I(N__44883));
    InMux I__10626 (
            .O(N__44907),
            .I(N__44880));
    InMux I__10625 (
            .O(N__44904),
            .I(N__44875));
    InMux I__10624 (
            .O(N__44903),
            .I(N__44868));
    InMux I__10623 (
            .O(N__44902),
            .I(N__44863));
    InMux I__10622 (
            .O(N__44899),
            .I(N__44863));
    LocalMux I__10621 (
            .O(N__44896),
            .I(N__44860));
    InMux I__10620 (
            .O(N__44893),
            .I(N__44855));
    InMux I__10619 (
            .O(N__44892),
            .I(N__44855));
    InMux I__10618 (
            .O(N__44891),
            .I(N__44848));
    InMux I__10617 (
            .O(N__44890),
            .I(N__44848));
    InMux I__10616 (
            .O(N__44887),
            .I(N__44845));
    InMux I__10615 (
            .O(N__44886),
            .I(N__44842));
    LocalMux I__10614 (
            .O(N__44883),
            .I(N__44837));
    LocalMux I__10613 (
            .O(N__44880),
            .I(N__44837));
    InMux I__10612 (
            .O(N__44879),
            .I(N__44832));
    InMux I__10611 (
            .O(N__44878),
            .I(N__44832));
    LocalMux I__10610 (
            .O(N__44875),
            .I(N__44827));
    InMux I__10609 (
            .O(N__44874),
            .I(N__44824));
    InMux I__10608 (
            .O(N__44873),
            .I(N__44819));
    InMux I__10607 (
            .O(N__44872),
            .I(N__44819));
    InMux I__10606 (
            .O(N__44871),
            .I(N__44816));
    LocalMux I__10605 (
            .O(N__44868),
            .I(N__44807));
    LocalMux I__10604 (
            .O(N__44863),
            .I(N__44807));
    Span4Mux_v I__10603 (
            .O(N__44860),
            .I(N__44807));
    LocalMux I__10602 (
            .O(N__44855),
            .I(N__44807));
    InMux I__10601 (
            .O(N__44854),
            .I(N__44802));
    InMux I__10600 (
            .O(N__44853),
            .I(N__44802));
    LocalMux I__10599 (
            .O(N__44848),
            .I(N__44799));
    LocalMux I__10598 (
            .O(N__44845),
            .I(N__44790));
    LocalMux I__10597 (
            .O(N__44842),
            .I(N__44790));
    Span4Mux_v I__10596 (
            .O(N__44837),
            .I(N__44790));
    LocalMux I__10595 (
            .O(N__44832),
            .I(N__44790));
    InMux I__10594 (
            .O(N__44831),
            .I(N__44787));
    InMux I__10593 (
            .O(N__44830),
            .I(N__44784));
    Span4Mux_v I__10592 (
            .O(N__44827),
            .I(N__44777));
    LocalMux I__10591 (
            .O(N__44824),
            .I(N__44777));
    LocalMux I__10590 (
            .O(N__44819),
            .I(N__44777));
    LocalMux I__10589 (
            .O(N__44816),
            .I(N__44770));
    Span4Mux_v I__10588 (
            .O(N__44807),
            .I(N__44770));
    LocalMux I__10587 (
            .O(N__44802),
            .I(N__44770));
    Span4Mux_v I__10586 (
            .O(N__44799),
            .I(N__44765));
    Span4Mux_v I__10585 (
            .O(N__44790),
            .I(N__44765));
    LocalMux I__10584 (
            .O(N__44787),
            .I(n6_adj_819));
    LocalMux I__10583 (
            .O(N__44784),
            .I(n6_adj_819));
    Odrv4 I__10582 (
            .O(N__44777),
            .I(n6_adj_819));
    Odrv4 I__10581 (
            .O(N__44770),
            .I(n6_adj_819));
    Odrv4 I__10580 (
            .O(N__44765),
            .I(n6_adj_819));
    CascadeMux I__10579 (
            .O(N__44754),
            .I(n8_adj_834_cascade_));
    IoInMux I__10578 (
            .O(N__44751),
            .I(N__44748));
    LocalMux I__10577 (
            .O(N__44748),
            .I(N__44745));
    Span4Mux_s1_v I__10576 (
            .O(N__44745),
            .I(N__44742));
    Sp12to4 I__10575 (
            .O(N__44742),
            .I(N__44739));
    Span12Mux_h I__10574 (
            .O(N__44739),
            .I(N__44734));
    InMux I__10573 (
            .O(N__44738),
            .I(N__44729));
    InMux I__10572 (
            .O(N__44737),
            .I(N__44729));
    Odrv12 I__10571 (
            .O(N__44734),
            .I(pin_out_17));
    LocalMux I__10570 (
            .O(N__44729),
            .I(pin_out_17));
    InMux I__10569 (
            .O(N__44724),
            .I(N__44721));
    LocalMux I__10568 (
            .O(N__44721),
            .I(n13631));
    IoInMux I__10567 (
            .O(N__44718),
            .I(N__44715));
    LocalMux I__10566 (
            .O(N__44715),
            .I(N__44712));
    Span4Mux_s0_h I__10565 (
            .O(N__44712),
            .I(N__44709));
    Sp12to4 I__10564 (
            .O(N__44709),
            .I(N__44705));
    CascadeMux I__10563 (
            .O(N__44708),
            .I(N__44702));
    Span12Mux_v I__10562 (
            .O(N__44705),
            .I(N__44699));
    InMux I__10561 (
            .O(N__44702),
            .I(N__44695));
    Span12Mux_h I__10560 (
            .O(N__44699),
            .I(N__44692));
    InMux I__10559 (
            .O(N__44698),
            .I(N__44689));
    LocalMux I__10558 (
            .O(N__44695),
            .I(N__44686));
    Odrv12 I__10557 (
            .O(N__44692),
            .I(pin_out_16));
    LocalMux I__10556 (
            .O(N__44689),
            .I(pin_out_16));
    Odrv12 I__10555 (
            .O(N__44686),
            .I(pin_out_16));
    CascadeMux I__10554 (
            .O(N__44679),
            .I(n13634_cascade_));
    InMux I__10553 (
            .O(N__44676),
            .I(N__44673));
    LocalMux I__10552 (
            .O(N__44673),
            .I(N__44670));
    Odrv4 I__10551 (
            .O(N__44670),
            .I(n13389));
    InMux I__10550 (
            .O(N__44667),
            .I(N__44664));
    LocalMux I__10549 (
            .O(N__44664),
            .I(n7_adj_838));
    InMux I__10548 (
            .O(N__44661),
            .I(N__44658));
    LocalMux I__10547 (
            .O(N__44658),
            .I(n7_adj_837));
    IoInMux I__10546 (
            .O(N__44655),
            .I(N__44652));
    LocalMux I__10545 (
            .O(N__44652),
            .I(N__44649));
    IoSpan4Mux I__10544 (
            .O(N__44649),
            .I(N__44646));
    Span4Mux_s3_v I__10543 (
            .O(N__44646),
            .I(N__44643));
    Span4Mux_v I__10542 (
            .O(N__44643),
            .I(N__44639));
    CascadeMux I__10541 (
            .O(N__44642),
            .I(N__44636));
    Span4Mux_v I__10540 (
            .O(N__44639),
            .I(N__44632));
    InMux I__10539 (
            .O(N__44636),
            .I(N__44629));
    InMux I__10538 (
            .O(N__44635),
            .I(N__44626));
    Odrv4 I__10537 (
            .O(N__44632),
            .I(pin_out_21));
    LocalMux I__10536 (
            .O(N__44629),
            .I(pin_out_21));
    LocalMux I__10535 (
            .O(N__44626),
            .I(pin_out_21));
    IoInMux I__10534 (
            .O(N__44619),
            .I(N__44616));
    LocalMux I__10533 (
            .O(N__44616),
            .I(N__44612));
    CascadeMux I__10532 (
            .O(N__44615),
            .I(N__44609));
    Span12Mux_s10_v I__10531 (
            .O(N__44612),
            .I(N__44605));
    InMux I__10530 (
            .O(N__44609),
            .I(N__44600));
    InMux I__10529 (
            .O(N__44608),
            .I(N__44600));
    Odrv12 I__10528 (
            .O(N__44605),
            .I(pin_out_20));
    LocalMux I__10527 (
            .O(N__44600),
            .I(pin_out_20));
    IoInMux I__10526 (
            .O(N__44595),
            .I(N__44592));
    LocalMux I__10525 (
            .O(N__44592),
            .I(N__44589));
    Span4Mux_s2_v I__10524 (
            .O(N__44589),
            .I(N__44586));
    Span4Mux_h I__10523 (
            .O(N__44586),
            .I(N__44582));
    InMux I__10522 (
            .O(N__44585),
            .I(N__44578));
    Sp12to4 I__10521 (
            .O(N__44582),
            .I(N__44575));
    InMux I__10520 (
            .O(N__44581),
            .I(N__44572));
    LocalMux I__10519 (
            .O(N__44578),
            .I(N__44569));
    Odrv12 I__10518 (
            .O(N__44575),
            .I(pin_out_22));
    LocalMux I__10517 (
            .O(N__44572),
            .I(pin_out_22));
    Odrv4 I__10516 (
            .O(N__44569),
            .I(pin_out_22));
    CascadeMux I__10515 (
            .O(N__44562),
            .I(n19_adj_790_cascade_));
    InMux I__10514 (
            .O(N__44559),
            .I(N__44556));
    LocalMux I__10513 (
            .O(N__44556),
            .I(n13388));
    CascadeMux I__10512 (
            .O(N__44553),
            .I(n7_adj_833_cascade_));
    InMux I__10511 (
            .O(N__44550),
            .I(N__44547));
    LocalMux I__10510 (
            .O(N__44547),
            .I(n8_adj_836));
    CascadeMux I__10509 (
            .O(N__44544),
            .I(N__44541));
    InMux I__10508 (
            .O(N__44541),
            .I(N__44526));
    InMux I__10507 (
            .O(N__44540),
            .I(N__44523));
    InMux I__10506 (
            .O(N__44539),
            .I(N__44520));
    InMux I__10505 (
            .O(N__44538),
            .I(N__44517));
    InMux I__10504 (
            .O(N__44537),
            .I(N__44514));
    InMux I__10503 (
            .O(N__44536),
            .I(N__44509));
    InMux I__10502 (
            .O(N__44535),
            .I(N__44509));
    InMux I__10501 (
            .O(N__44534),
            .I(N__44504));
    InMux I__10500 (
            .O(N__44533),
            .I(N__44504));
    InMux I__10499 (
            .O(N__44532),
            .I(N__44500));
    InMux I__10498 (
            .O(N__44531),
            .I(N__44497));
    InMux I__10497 (
            .O(N__44530),
            .I(N__44494));
    InMux I__10496 (
            .O(N__44529),
            .I(N__44491));
    LocalMux I__10495 (
            .O(N__44526),
            .I(N__44488));
    LocalMux I__10494 (
            .O(N__44523),
            .I(N__44485));
    LocalMux I__10493 (
            .O(N__44520),
            .I(N__44474));
    LocalMux I__10492 (
            .O(N__44517),
            .I(N__44474));
    LocalMux I__10491 (
            .O(N__44514),
            .I(N__44474));
    LocalMux I__10490 (
            .O(N__44509),
            .I(N__44474));
    LocalMux I__10489 (
            .O(N__44504),
            .I(N__44474));
    InMux I__10488 (
            .O(N__44503),
            .I(N__44471));
    LocalMux I__10487 (
            .O(N__44500),
            .I(N__44468));
    LocalMux I__10486 (
            .O(N__44497),
            .I(N__44463));
    LocalMux I__10485 (
            .O(N__44494),
            .I(N__44463));
    LocalMux I__10484 (
            .O(N__44491),
            .I(N__44460));
    Span4Mux_v I__10483 (
            .O(N__44488),
            .I(N__44453));
    Span4Mux_h I__10482 (
            .O(N__44485),
            .I(N__44453));
    Span4Mux_v I__10481 (
            .O(N__44474),
            .I(N__44453));
    LocalMux I__10480 (
            .O(N__44471),
            .I(n7_adj_811));
    Odrv4 I__10479 (
            .O(N__44468),
            .I(n7_adj_811));
    Odrv4 I__10478 (
            .O(N__44463),
            .I(n7_adj_811));
    Odrv4 I__10477 (
            .O(N__44460),
            .I(n7_adj_811));
    Odrv4 I__10476 (
            .O(N__44453),
            .I(n7_adj_811));
    CascadeMux I__10475 (
            .O(N__44442),
            .I(n7_adj_835_cascade_));
    CascadeMux I__10474 (
            .O(N__44439),
            .I(N__44436));
    InMux I__10473 (
            .O(N__44436),
            .I(N__44432));
    InMux I__10472 (
            .O(N__44435),
            .I(N__44427));
    LocalMux I__10471 (
            .O(N__44432),
            .I(N__44423));
    InMux I__10470 (
            .O(N__44431),
            .I(N__44418));
    InMux I__10469 (
            .O(N__44430),
            .I(N__44415));
    LocalMux I__10468 (
            .O(N__44427),
            .I(N__44412));
    InMux I__10467 (
            .O(N__44426),
            .I(N__44409));
    Span4Mux_v I__10466 (
            .O(N__44423),
            .I(N__44406));
    InMux I__10465 (
            .O(N__44422),
            .I(N__44402));
    InMux I__10464 (
            .O(N__44421),
            .I(N__44399));
    LocalMux I__10463 (
            .O(N__44418),
            .I(N__44396));
    LocalMux I__10462 (
            .O(N__44415),
            .I(N__44393));
    Span4Mux_v I__10461 (
            .O(N__44412),
            .I(N__44390));
    LocalMux I__10460 (
            .O(N__44409),
            .I(N__44384));
    Span4Mux_h I__10459 (
            .O(N__44406),
            .I(N__44381));
    InMux I__10458 (
            .O(N__44405),
            .I(N__44378));
    LocalMux I__10457 (
            .O(N__44402),
            .I(N__44375));
    LocalMux I__10456 (
            .O(N__44399),
            .I(N__44372));
    Span4Mux_h I__10455 (
            .O(N__44396),
            .I(N__44367));
    Span4Mux_h I__10454 (
            .O(N__44393),
            .I(N__44367));
    Span4Mux_h I__10453 (
            .O(N__44390),
            .I(N__44364));
    InMux I__10452 (
            .O(N__44389),
            .I(N__44361));
    InMux I__10451 (
            .O(N__44388),
            .I(N__44358));
    InMux I__10450 (
            .O(N__44387),
            .I(N__44355));
    Span4Mux_v I__10449 (
            .O(N__44384),
            .I(N__44350));
    Span4Mux_h I__10448 (
            .O(N__44381),
            .I(N__44350));
    LocalMux I__10447 (
            .O(N__44378),
            .I(N__44339));
    Span4Mux_v I__10446 (
            .O(N__44375),
            .I(N__44339));
    Span4Mux_v I__10445 (
            .O(N__44372),
            .I(N__44339));
    Span4Mux_v I__10444 (
            .O(N__44367),
            .I(N__44339));
    Span4Mux_h I__10443 (
            .O(N__44364),
            .I(N__44339));
    LocalMux I__10442 (
            .O(N__44361),
            .I(n6_adj_810));
    LocalMux I__10441 (
            .O(N__44358),
            .I(n6_adj_810));
    LocalMux I__10440 (
            .O(N__44355),
            .I(n6_adj_810));
    Odrv4 I__10439 (
            .O(N__44350),
            .I(n6_adj_810));
    Odrv4 I__10438 (
            .O(N__44339),
            .I(n6_adj_810));
    CascadeMux I__10437 (
            .O(N__44328),
            .I(n7_adj_839_cascade_));
    IoInMux I__10436 (
            .O(N__44325),
            .I(N__44322));
    LocalMux I__10435 (
            .O(N__44322),
            .I(N__44319));
    IoSpan4Mux I__10434 (
            .O(N__44319),
            .I(N__44316));
    Sp12to4 I__10433 (
            .O(N__44316),
            .I(N__44313));
    Span12Mux_s6_v I__10432 (
            .O(N__44313),
            .I(N__44310));
    Span12Mux_h I__10431 (
            .O(N__44310),
            .I(N__44305));
    InMux I__10430 (
            .O(N__44309),
            .I(N__44302));
    InMux I__10429 (
            .O(N__44308),
            .I(N__44299));
    Odrv12 I__10428 (
            .O(N__44305),
            .I(pin_out_18));
    LocalMux I__10427 (
            .O(N__44302),
            .I(pin_out_18));
    LocalMux I__10426 (
            .O(N__44299),
            .I(pin_out_18));
    IoInMux I__10425 (
            .O(N__44292),
            .I(N__44289));
    LocalMux I__10424 (
            .O(N__44289),
            .I(N__44286));
    IoSpan4Mux I__10423 (
            .O(N__44286),
            .I(N__44283));
    Span4Mux_s1_v I__10422 (
            .O(N__44283),
            .I(N__44279));
    CascadeMux I__10421 (
            .O(N__44282),
            .I(N__44275));
    Sp12to4 I__10420 (
            .O(N__44279),
            .I(N__44272));
    CascadeMux I__10419 (
            .O(N__44278),
            .I(N__44269));
    InMux I__10418 (
            .O(N__44275),
            .I(N__44266));
    Span12Mux_v I__10417 (
            .O(N__44272),
            .I(N__44263));
    InMux I__10416 (
            .O(N__44269),
            .I(N__44260));
    LocalMux I__10415 (
            .O(N__44266),
            .I(N__44257));
    Odrv12 I__10414 (
            .O(N__44263),
            .I(pin_out_19));
    LocalMux I__10413 (
            .O(N__44260),
            .I(pin_out_19));
    Odrv4 I__10412 (
            .O(N__44257),
            .I(pin_out_19));
    CascadeMux I__10411 (
            .O(N__44250),
            .I(n11962_cascade_));
    IoInMux I__10410 (
            .O(N__44247),
            .I(N__44244));
    LocalMux I__10409 (
            .O(N__44244),
            .I(N__44241));
    Span4Mux_s3_h I__10408 (
            .O(N__44241),
            .I(N__44238));
    Span4Mux_v I__10407 (
            .O(N__44238),
            .I(N__44235));
    Sp12to4 I__10406 (
            .O(N__44235),
            .I(N__44232));
    Span12Mux_h I__10405 (
            .O(N__44232),
            .I(N__44228));
    InMux I__10404 (
            .O(N__44231),
            .I(N__44225));
    Odrv12 I__10403 (
            .O(N__44228),
            .I(pin_oe_14));
    LocalMux I__10402 (
            .O(N__44225),
            .I(pin_oe_14));
    InMux I__10401 (
            .O(N__44220),
            .I(N__44216));
    InMux I__10400 (
            .O(N__44219),
            .I(N__44213));
    LocalMux I__10399 (
            .O(N__44216),
            .I(N__44210));
    LocalMux I__10398 (
            .O(N__44213),
            .I(N__44207));
    Span4Mux_v I__10397 (
            .O(N__44210),
            .I(N__44204));
    Odrv4 I__10396 (
            .O(N__44207),
            .I(n9_adj_812));
    Odrv4 I__10395 (
            .O(N__44204),
            .I(n9_adj_812));
    CascadeMux I__10394 (
            .O(N__44199),
            .I(N__44196));
    InMux I__10393 (
            .O(N__44196),
            .I(N__44193));
    LocalMux I__10392 (
            .O(N__44193),
            .I(n8_adj_828));
    CascadeMux I__10391 (
            .O(N__44190),
            .I(n11958_cascade_));
    IoInMux I__10390 (
            .O(N__44187),
            .I(N__44184));
    LocalMux I__10389 (
            .O(N__44184),
            .I(N__44181));
    Span4Mux_s0_v I__10388 (
            .O(N__44181),
            .I(N__44178));
    Span4Mux_v I__10387 (
            .O(N__44178),
            .I(N__44175));
    Sp12to4 I__10386 (
            .O(N__44175),
            .I(N__44172));
    Span12Mux_h I__10385 (
            .O(N__44172),
            .I(N__44169));
    Span12Mux_v I__10384 (
            .O(N__44169),
            .I(N__44165));
    InMux I__10383 (
            .O(N__44168),
            .I(N__44162));
    Odrv12 I__10382 (
            .O(N__44165),
            .I(pin_oe_21));
    LocalMux I__10381 (
            .O(N__44162),
            .I(pin_oe_21));
    InMux I__10380 (
            .O(N__44157),
            .I(N__44154));
    LocalMux I__10379 (
            .O(N__44154),
            .I(N__44151));
    Span4Mux_v I__10378 (
            .O(N__44151),
            .I(N__44148));
    Sp12to4 I__10377 (
            .O(N__44148),
            .I(N__44145));
    Span12Mux_h I__10376 (
            .O(N__44145),
            .I(N__44142));
    Odrv12 I__10375 (
            .O(N__44142),
            .I(n13652));
    CascadeMux I__10374 (
            .O(N__44139),
            .I(n13536_cascade_));
    InMux I__10373 (
            .O(N__44136),
            .I(N__44133));
    LocalMux I__10372 (
            .O(N__44133),
            .I(N__44130));
    Span12Mux_h I__10371 (
            .O(N__44130),
            .I(N__44127));
    Odrv12 I__10370 (
            .O(N__44127),
            .I(n13616));
    InMux I__10369 (
            .O(N__44124),
            .I(N__44121));
    LocalMux I__10368 (
            .O(N__44121),
            .I(n13542));
    CascadeMux I__10367 (
            .O(N__44118),
            .I(n7_adj_831_cascade_));
    CascadeMux I__10366 (
            .O(N__44115),
            .I(N__44108));
    CascadeMux I__10365 (
            .O(N__44114),
            .I(N__44102));
    CascadeMux I__10364 (
            .O(N__44113),
            .I(N__44099));
    InMux I__10363 (
            .O(N__44112),
            .I(N__44096));
    CascadeMux I__10362 (
            .O(N__44111),
            .I(N__44092));
    InMux I__10361 (
            .O(N__44108),
            .I(N__44088));
    InMux I__10360 (
            .O(N__44107),
            .I(N__44085));
    InMux I__10359 (
            .O(N__44106),
            .I(N__44082));
    InMux I__10358 (
            .O(N__44105),
            .I(N__44079));
    InMux I__10357 (
            .O(N__44102),
            .I(N__44076));
    InMux I__10356 (
            .O(N__44099),
            .I(N__44073));
    LocalMux I__10355 (
            .O(N__44096),
            .I(N__44070));
    InMux I__10354 (
            .O(N__44095),
            .I(N__44067));
    InMux I__10353 (
            .O(N__44092),
            .I(N__44064));
    InMux I__10352 (
            .O(N__44091),
            .I(N__44060));
    LocalMux I__10351 (
            .O(N__44088),
            .I(N__44055));
    LocalMux I__10350 (
            .O(N__44085),
            .I(N__44055));
    LocalMux I__10349 (
            .O(N__44082),
            .I(N__44052));
    LocalMux I__10348 (
            .O(N__44079),
            .I(N__44047));
    LocalMux I__10347 (
            .O(N__44076),
            .I(N__44047));
    LocalMux I__10346 (
            .O(N__44073),
            .I(N__44044));
    Span4Mux_v I__10345 (
            .O(N__44070),
            .I(N__44041));
    LocalMux I__10344 (
            .O(N__44067),
            .I(N__44036));
    LocalMux I__10343 (
            .O(N__44064),
            .I(N__44036));
    InMux I__10342 (
            .O(N__44063),
            .I(N__44033));
    LocalMux I__10341 (
            .O(N__44060),
            .I(N__44028));
    Span4Mux_h I__10340 (
            .O(N__44055),
            .I(N__44028));
    Span4Mux_h I__10339 (
            .O(N__44052),
            .I(N__44021));
    Span4Mux_h I__10338 (
            .O(N__44047),
            .I(N__44021));
    Span4Mux_h I__10337 (
            .O(N__44044),
            .I(N__44021));
    Span4Mux_h I__10336 (
            .O(N__44041),
            .I(N__44016));
    Span4Mux_v I__10335 (
            .O(N__44036),
            .I(N__44016));
    LocalMux I__10334 (
            .O(N__44033),
            .I(n6_adj_813));
    Odrv4 I__10333 (
            .O(N__44028),
            .I(n6_adj_813));
    Odrv4 I__10332 (
            .O(N__44021),
            .I(n6_adj_813));
    Odrv4 I__10331 (
            .O(N__44016),
            .I(n6_adj_813));
    CascadeMux I__10330 (
            .O(N__44007),
            .I(n11825_cascade_));
    IoInMux I__10329 (
            .O(N__44004),
            .I(N__44001));
    LocalMux I__10328 (
            .O(N__44001),
            .I(N__43998));
    IoSpan4Mux I__10327 (
            .O(N__43998),
            .I(N__43995));
    Span4Mux_s3_h I__10326 (
            .O(N__43995),
            .I(N__43992));
    Span4Mux_h I__10325 (
            .O(N__43992),
            .I(N__43989));
    Span4Mux_h I__10324 (
            .O(N__43989),
            .I(N__43985));
    InMux I__10323 (
            .O(N__43988),
            .I(N__43982));
    Odrv4 I__10322 (
            .O(N__43985),
            .I(pin_oe_15));
    LocalMux I__10321 (
            .O(N__43982),
            .I(pin_oe_15));
    InMux I__10320 (
            .O(N__43977),
            .I(N__43971));
    InMux I__10319 (
            .O(N__43976),
            .I(N__43971));
    LocalMux I__10318 (
            .O(N__43971),
            .I(N__43968));
    Span4Mux_h I__10317 (
            .O(N__43968),
            .I(N__43965));
    Span4Mux_h I__10316 (
            .O(N__43965),
            .I(N__43962));
    Span4Mux_h I__10315 (
            .O(N__43962),
            .I(N__43959));
    Odrv4 I__10314 (
            .O(N__43959),
            .I(n1907));
    CascadeMux I__10313 (
            .O(N__43956),
            .I(N__43952));
    InMux I__10312 (
            .O(N__43955),
            .I(N__43948));
    InMux I__10311 (
            .O(N__43952),
            .I(N__43944));
    InMux I__10310 (
            .O(N__43951),
            .I(N__43941));
    LocalMux I__10309 (
            .O(N__43948),
            .I(N__43936));
    InMux I__10308 (
            .O(N__43947),
            .I(N__43933));
    LocalMux I__10307 (
            .O(N__43944),
            .I(N__43929));
    LocalMux I__10306 (
            .O(N__43941),
            .I(N__43926));
    CascadeMux I__10305 (
            .O(N__43940),
            .I(N__43922));
    InMux I__10304 (
            .O(N__43939),
            .I(N__43919));
    Span4Mux_v I__10303 (
            .O(N__43936),
            .I(N__43916));
    LocalMux I__10302 (
            .O(N__43933),
            .I(N__43913));
    InMux I__10301 (
            .O(N__43932),
            .I(N__43907));
    Span4Mux_v I__10300 (
            .O(N__43929),
            .I(N__43902));
    Span4Mux_h I__10299 (
            .O(N__43926),
            .I(N__43902));
    InMux I__10298 (
            .O(N__43925),
            .I(N__43899));
    InMux I__10297 (
            .O(N__43922),
            .I(N__43887));
    LocalMux I__10296 (
            .O(N__43919),
            .I(N__43884));
    Span4Mux_h I__10295 (
            .O(N__43916),
            .I(N__43879));
    Span4Mux_v I__10294 (
            .O(N__43913),
            .I(N__43879));
    CascadeMux I__10293 (
            .O(N__43912),
            .I(N__43876));
    InMux I__10292 (
            .O(N__43911),
            .I(N__43869));
    InMux I__10291 (
            .O(N__43910),
            .I(N__43869));
    LocalMux I__10290 (
            .O(N__43907),
            .I(N__43866));
    Span4Mux_v I__10289 (
            .O(N__43902),
            .I(N__43861));
    LocalMux I__10288 (
            .O(N__43899),
            .I(N__43861));
    InMux I__10287 (
            .O(N__43898),
            .I(N__43858));
    InMux I__10286 (
            .O(N__43897),
            .I(N__43853));
    InMux I__10285 (
            .O(N__43896),
            .I(N__43853));
    InMux I__10284 (
            .O(N__43895),
            .I(N__43846));
    InMux I__10283 (
            .O(N__43894),
            .I(N__43846));
    InMux I__10282 (
            .O(N__43893),
            .I(N__43846));
    InMux I__10281 (
            .O(N__43892),
            .I(N__43843));
    InMux I__10280 (
            .O(N__43891),
            .I(N__43840));
    CascadeMux I__10279 (
            .O(N__43890),
            .I(N__43837));
    LocalMux I__10278 (
            .O(N__43887),
            .I(N__43833));
    Span4Mux_v I__10277 (
            .O(N__43884),
            .I(N__43828));
    Span4Mux_v I__10276 (
            .O(N__43879),
            .I(N__43828));
    InMux I__10275 (
            .O(N__43876),
            .I(N__43825));
    CascadeMux I__10274 (
            .O(N__43875),
            .I(N__43819));
    InMux I__10273 (
            .O(N__43874),
            .I(N__43814));
    LocalMux I__10272 (
            .O(N__43869),
            .I(N__43811));
    Span4Mux_h I__10271 (
            .O(N__43866),
            .I(N__43806));
    Span4Mux_v I__10270 (
            .O(N__43861),
            .I(N__43806));
    LocalMux I__10269 (
            .O(N__43858),
            .I(N__43797));
    LocalMux I__10268 (
            .O(N__43853),
            .I(N__43797));
    LocalMux I__10267 (
            .O(N__43846),
            .I(N__43797));
    LocalMux I__10266 (
            .O(N__43843),
            .I(N__43797));
    LocalMux I__10265 (
            .O(N__43840),
            .I(N__43794));
    InMux I__10264 (
            .O(N__43837),
            .I(N__43791));
    InMux I__10263 (
            .O(N__43836),
            .I(N__43788));
    Span12Mux_v I__10262 (
            .O(N__43833),
            .I(N__43783));
    Sp12to4 I__10261 (
            .O(N__43828),
            .I(N__43783));
    LocalMux I__10260 (
            .O(N__43825),
            .I(N__43780));
    InMux I__10259 (
            .O(N__43824),
            .I(N__43777));
    InMux I__10258 (
            .O(N__43823),
            .I(N__43774));
    InMux I__10257 (
            .O(N__43822),
            .I(N__43771));
    InMux I__10256 (
            .O(N__43819),
            .I(N__43768));
    InMux I__10255 (
            .O(N__43818),
            .I(N__43765));
    InMux I__10254 (
            .O(N__43817),
            .I(N__43762));
    LocalMux I__10253 (
            .O(N__43814),
            .I(N__43755));
    Span4Mux_v I__10252 (
            .O(N__43811),
            .I(N__43755));
    Span4Mux_h I__10251 (
            .O(N__43806),
            .I(N__43755));
    Span12Mux_v I__10250 (
            .O(N__43797),
            .I(N__43752));
    Span4Mux_h I__10249 (
            .O(N__43794),
            .I(N__43745));
    LocalMux I__10248 (
            .O(N__43791),
            .I(N__43745));
    LocalMux I__10247 (
            .O(N__43788),
            .I(N__43745));
    Span12Mux_h I__10246 (
            .O(N__43783),
            .I(N__43740));
    Span12Mux_h I__10245 (
            .O(N__43780),
            .I(N__43740));
    LocalMux I__10244 (
            .O(N__43777),
            .I(N__43737));
    LocalMux I__10243 (
            .O(N__43774),
            .I(state_1));
    LocalMux I__10242 (
            .O(N__43771),
            .I(state_1));
    LocalMux I__10241 (
            .O(N__43768),
            .I(state_1));
    LocalMux I__10240 (
            .O(N__43765),
            .I(state_1));
    LocalMux I__10239 (
            .O(N__43762),
            .I(state_1));
    Odrv4 I__10238 (
            .O(N__43755),
            .I(state_1));
    Odrv12 I__10237 (
            .O(N__43752),
            .I(state_1));
    Odrv4 I__10236 (
            .O(N__43745),
            .I(state_1));
    Odrv12 I__10235 (
            .O(N__43740),
            .I(state_1));
    Odrv4 I__10234 (
            .O(N__43737),
            .I(state_1));
    InMux I__10233 (
            .O(N__43716),
            .I(N__43712));
    CascadeMux I__10232 (
            .O(N__43715),
            .I(N__43708));
    LocalMux I__10231 (
            .O(N__43712),
            .I(N__43705));
    InMux I__10230 (
            .O(N__43711),
            .I(N__43702));
    InMux I__10229 (
            .O(N__43708),
            .I(N__43698));
    Span4Mux_h I__10228 (
            .O(N__43705),
            .I(N__43693));
    LocalMux I__10227 (
            .O(N__43702),
            .I(N__43693));
    CascadeMux I__10226 (
            .O(N__43701),
            .I(N__43688));
    LocalMux I__10225 (
            .O(N__43698),
            .I(N__43685));
    Span4Mux_v I__10224 (
            .O(N__43693),
            .I(N__43682));
    CascadeMux I__10223 (
            .O(N__43692),
            .I(N__43677));
    CascadeMux I__10222 (
            .O(N__43691),
            .I(N__43672));
    InMux I__10221 (
            .O(N__43688),
            .I(N__43669));
    Span4Mux_v I__10220 (
            .O(N__43685),
            .I(N__43663));
    Span4Mux_v I__10219 (
            .O(N__43682),
            .I(N__43663));
    InMux I__10218 (
            .O(N__43681),
            .I(N__43660));
    InMux I__10217 (
            .O(N__43680),
            .I(N__43653));
    InMux I__10216 (
            .O(N__43677),
            .I(N__43653));
    InMux I__10215 (
            .O(N__43676),
            .I(N__43653));
    InMux I__10214 (
            .O(N__43675),
            .I(N__43648));
    InMux I__10213 (
            .O(N__43672),
            .I(N__43645));
    LocalMux I__10212 (
            .O(N__43669),
            .I(N__43642));
    CascadeMux I__10211 (
            .O(N__43668),
            .I(N__43637));
    Span4Mux_h I__10210 (
            .O(N__43663),
            .I(N__43632));
    LocalMux I__10209 (
            .O(N__43660),
            .I(N__43632));
    LocalMux I__10208 (
            .O(N__43653),
            .I(N__43629));
    InMux I__10207 (
            .O(N__43652),
            .I(N__43626));
    CascadeMux I__10206 (
            .O(N__43651),
            .I(N__43622));
    LocalMux I__10205 (
            .O(N__43648),
            .I(N__43619));
    LocalMux I__10204 (
            .O(N__43645),
            .I(N__43614));
    Span4Mux_h I__10203 (
            .O(N__43642),
            .I(N__43614));
    InMux I__10202 (
            .O(N__43641),
            .I(N__43611));
    InMux I__10201 (
            .O(N__43640),
            .I(N__43606));
    InMux I__10200 (
            .O(N__43637),
            .I(N__43606));
    Span4Mux_v I__10199 (
            .O(N__43632),
            .I(N__43601));
    Span4Mux_v I__10198 (
            .O(N__43629),
            .I(N__43601));
    LocalMux I__10197 (
            .O(N__43626),
            .I(N__43597));
    InMux I__10196 (
            .O(N__43625),
            .I(N__43593));
    InMux I__10195 (
            .O(N__43622),
            .I(N__43589));
    Span12Mux_v I__10194 (
            .O(N__43619),
            .I(N__43585));
    Span4Mux_v I__10193 (
            .O(N__43614),
            .I(N__43581));
    LocalMux I__10192 (
            .O(N__43611),
            .I(N__43576));
    LocalMux I__10191 (
            .O(N__43606),
            .I(N__43576));
    Span4Mux_h I__10190 (
            .O(N__43601),
            .I(N__43573));
    InMux I__10189 (
            .O(N__43600),
            .I(N__43570));
    Sp12to4 I__10188 (
            .O(N__43597),
            .I(N__43567));
    InMux I__10187 (
            .O(N__43596),
            .I(N__43564));
    LocalMux I__10186 (
            .O(N__43593),
            .I(N__43561));
    InMux I__10185 (
            .O(N__43592),
            .I(N__43558));
    LocalMux I__10184 (
            .O(N__43589),
            .I(N__43555));
    InMux I__10183 (
            .O(N__43588),
            .I(N__43552));
    Span12Mux_h I__10182 (
            .O(N__43585),
            .I(N__43549));
    InMux I__10181 (
            .O(N__43584),
            .I(N__43546));
    Span4Mux_h I__10180 (
            .O(N__43581),
            .I(N__43541));
    Span4Mux_v I__10179 (
            .O(N__43576),
            .I(N__43541));
    Span4Mux_h I__10178 (
            .O(N__43573),
            .I(N__43536));
    LocalMux I__10177 (
            .O(N__43570),
            .I(N__43536));
    Span12Mux_v I__10176 (
            .O(N__43567),
            .I(N__43533));
    LocalMux I__10175 (
            .O(N__43564),
            .I(N__43528));
    Span12Mux_h I__10174 (
            .O(N__43561),
            .I(N__43528));
    LocalMux I__10173 (
            .O(N__43558),
            .I(N__43521));
    Span4Mux_v I__10172 (
            .O(N__43555),
            .I(N__43521));
    LocalMux I__10171 (
            .O(N__43552),
            .I(N__43521));
    Odrv12 I__10170 (
            .O(N__43549),
            .I(state_2));
    LocalMux I__10169 (
            .O(N__43546),
            .I(state_2));
    Odrv4 I__10168 (
            .O(N__43541),
            .I(state_2));
    Odrv4 I__10167 (
            .O(N__43536),
            .I(state_2));
    Odrv12 I__10166 (
            .O(N__43533),
            .I(state_2));
    Odrv12 I__10165 (
            .O(N__43528),
            .I(state_2));
    Odrv4 I__10164 (
            .O(N__43521),
            .I(state_2));
    SRMux I__10163 (
            .O(N__43506),
            .I(N__43502));
    SRMux I__10162 (
            .O(N__43505),
            .I(N__43499));
    LocalMux I__10161 (
            .O(N__43502),
            .I(N__43496));
    LocalMux I__10160 (
            .O(N__43499),
            .I(N__43493));
    Span4Mux_s1_h I__10159 (
            .O(N__43496),
            .I(N__43486));
    Span4Mux_v I__10158 (
            .O(N__43493),
            .I(N__43486));
    SRMux I__10157 (
            .O(N__43492),
            .I(N__43483));
    SRMux I__10156 (
            .O(N__43491),
            .I(N__43480));
    Span4Mux_v I__10155 (
            .O(N__43486),
            .I(N__43473));
    LocalMux I__10154 (
            .O(N__43483),
            .I(N__43473));
    LocalMux I__10153 (
            .O(N__43480),
            .I(N__43473));
    Span4Mux_v I__10152 (
            .O(N__43473),
            .I(N__43470));
    Sp12to4 I__10151 (
            .O(N__43470),
            .I(N__43467));
    Span12Mux_s5_h I__10150 (
            .O(N__43467),
            .I(N__43464));
    Span12Mux_h I__10149 (
            .O(N__43464),
            .I(N__43461));
    Odrv12 I__10148 (
            .O(N__43461),
            .I(n8025));
    CascadeMux I__10147 (
            .O(N__43458),
            .I(n11954_cascade_));
    IoInMux I__10146 (
            .O(N__43455),
            .I(N__43452));
    LocalMux I__10145 (
            .O(N__43452),
            .I(N__43449));
    IoSpan4Mux I__10144 (
            .O(N__43449),
            .I(N__43446));
    Sp12to4 I__10143 (
            .O(N__43446),
            .I(N__43443));
    Span12Mux_v I__10142 (
            .O(N__43443),
            .I(N__43439));
    InMux I__10141 (
            .O(N__43442),
            .I(N__43436));
    Odrv12 I__10140 (
            .O(N__43439),
            .I(pin_oe_20));
    LocalMux I__10139 (
            .O(N__43436),
            .I(pin_oe_20));
    InMux I__10138 (
            .O(N__43431),
            .I(N__43425));
    InMux I__10137 (
            .O(N__43430),
            .I(N__43421));
    InMux I__10136 (
            .O(N__43429),
            .I(N__43418));
    InMux I__10135 (
            .O(N__43428),
            .I(N__43415));
    LocalMux I__10134 (
            .O(N__43425),
            .I(N__43411));
    InMux I__10133 (
            .O(N__43424),
            .I(N__43408));
    LocalMux I__10132 (
            .O(N__43421),
            .I(N__43405));
    LocalMux I__10131 (
            .O(N__43418),
            .I(N__43402));
    LocalMux I__10130 (
            .O(N__43415),
            .I(N__43399));
    InMux I__10129 (
            .O(N__43414),
            .I(N__43395));
    Span4Mux_v I__10128 (
            .O(N__43411),
            .I(N__43392));
    LocalMux I__10127 (
            .O(N__43408),
            .I(N__43389));
    Span4Mux_h I__10126 (
            .O(N__43405),
            .I(N__43386));
    Span4Mux_h I__10125 (
            .O(N__43402),
            .I(N__43381));
    Span4Mux_h I__10124 (
            .O(N__43399),
            .I(N__43381));
    InMux I__10123 (
            .O(N__43398),
            .I(N__43378));
    LocalMux I__10122 (
            .O(N__43395),
            .I(n9488));
    Odrv4 I__10121 (
            .O(N__43392),
            .I(n9488));
    Odrv12 I__10120 (
            .O(N__43389),
            .I(n9488));
    Odrv4 I__10119 (
            .O(N__43386),
            .I(n9488));
    Odrv4 I__10118 (
            .O(N__43381),
            .I(n9488));
    LocalMux I__10117 (
            .O(N__43378),
            .I(n9488));
    InMux I__10116 (
            .O(N__43365),
            .I(N__43362));
    LocalMux I__10115 (
            .O(N__43362),
            .I(n11821));
    InMux I__10114 (
            .O(N__43359),
            .I(N__43356));
    LocalMux I__10113 (
            .O(N__43356),
            .I(n8_adj_826));
    IoInMux I__10112 (
            .O(N__43353),
            .I(N__43350));
    LocalMux I__10111 (
            .O(N__43350),
            .I(N__43347));
    IoSpan4Mux I__10110 (
            .O(N__43347),
            .I(N__43344));
    IoSpan4Mux I__10109 (
            .O(N__43344),
            .I(N__43341));
    Span4Mux_s3_v I__10108 (
            .O(N__43341),
            .I(N__43337));
    InMux I__10107 (
            .O(N__43340),
            .I(N__43333));
    Sp12to4 I__10106 (
            .O(N__43337),
            .I(N__43330));
    CascadeMux I__10105 (
            .O(N__43336),
            .I(N__43327));
    LocalMux I__10104 (
            .O(N__43333),
            .I(N__43324));
    Span12Mux_s10_v I__10103 (
            .O(N__43330),
            .I(N__43321));
    InMux I__10102 (
            .O(N__43327),
            .I(N__43318));
    Span4Mux_h I__10101 (
            .O(N__43324),
            .I(N__43315));
    Odrv12 I__10100 (
            .O(N__43321),
            .I(pin_out_8));
    LocalMux I__10099 (
            .O(N__43318),
            .I(pin_out_8));
    Odrv4 I__10098 (
            .O(N__43315),
            .I(pin_out_8));
    InMux I__10097 (
            .O(N__43308),
            .I(N__43305));
    LocalMux I__10096 (
            .O(N__43305),
            .I(n8_adj_832));
    InMux I__10095 (
            .O(N__43302),
            .I(N__43299));
    LocalMux I__10094 (
            .O(N__43299),
            .I(pin_out_22__N_216));
    CascadeMux I__10093 (
            .O(N__43296),
            .I(pin_out_22__N_216_cascade_));
    InMux I__10092 (
            .O(N__43293),
            .I(N__43290));
    LocalMux I__10091 (
            .O(N__43290),
            .I(N__43287));
    Odrv4 I__10090 (
            .O(N__43287),
            .I(n13370));
    CascadeMux I__10089 (
            .O(N__43284),
            .I(N__43281));
    InMux I__10088 (
            .O(N__43281),
            .I(N__43278));
    LocalMux I__10087 (
            .O(N__43278),
            .I(N__43275));
    Odrv4 I__10086 (
            .O(N__43275),
            .I(n13369));
    CascadeMux I__10085 (
            .O(N__43272),
            .I(n13640_cascade_));
    InMux I__10084 (
            .O(N__43269),
            .I(N__43266));
    LocalMux I__10083 (
            .O(N__43266),
            .I(N__43263));
    Span4Mux_h I__10082 (
            .O(N__43263),
            .I(N__43260));
    Odrv4 I__10081 (
            .O(N__43260),
            .I(n13628));
    CascadeMux I__10080 (
            .O(N__43257),
            .I(N__43254));
    InMux I__10079 (
            .O(N__43254),
            .I(N__43251));
    LocalMux I__10078 (
            .O(N__43251),
            .I(n13540));
    InMux I__10077 (
            .O(N__43248),
            .I(N__43245));
    LocalMux I__10076 (
            .O(N__43245),
            .I(N__43233));
    InMux I__10075 (
            .O(N__43244),
            .I(N__43230));
    InMux I__10074 (
            .O(N__43243),
            .I(N__43225));
    InMux I__10073 (
            .O(N__43242),
            .I(N__43225));
    InMux I__10072 (
            .O(N__43241),
            .I(N__43218));
    InMux I__10071 (
            .O(N__43240),
            .I(N__43218));
    InMux I__10070 (
            .O(N__43239),
            .I(N__43218));
    InMux I__10069 (
            .O(N__43238),
            .I(N__43211));
    InMux I__10068 (
            .O(N__43237),
            .I(N__43211));
    InMux I__10067 (
            .O(N__43236),
            .I(N__43211));
    Odrv4 I__10066 (
            .O(N__43233),
            .I(current_pin_4));
    LocalMux I__10065 (
            .O(N__43230),
            .I(current_pin_4));
    LocalMux I__10064 (
            .O(N__43225),
            .I(current_pin_4));
    LocalMux I__10063 (
            .O(N__43218),
            .I(current_pin_4));
    LocalMux I__10062 (
            .O(N__43211),
            .I(current_pin_4));
    CascadeMux I__10061 (
            .O(N__43200),
            .I(n7_adj_797_cascade_));
    InMux I__10060 (
            .O(N__43197),
            .I(N__43194));
    LocalMux I__10059 (
            .O(N__43194),
            .I(n13551));
    CascadeMux I__10058 (
            .O(N__43191),
            .I(N__43187));
    InMux I__10057 (
            .O(N__43190),
            .I(N__43180));
    InMux I__10056 (
            .O(N__43187),
            .I(N__43175));
    InMux I__10055 (
            .O(N__43186),
            .I(N__43175));
    CascadeMux I__10054 (
            .O(N__43185),
            .I(N__43171));
    InMux I__10053 (
            .O(N__43184),
            .I(N__43168));
    CascadeMux I__10052 (
            .O(N__43183),
            .I(N__43165));
    LocalMux I__10051 (
            .O(N__43180),
            .I(N__43160));
    LocalMux I__10050 (
            .O(N__43175),
            .I(N__43160));
    InMux I__10049 (
            .O(N__43174),
            .I(N__43157));
    InMux I__10048 (
            .O(N__43171),
            .I(N__43154));
    LocalMux I__10047 (
            .O(N__43168),
            .I(N__43151));
    InMux I__10046 (
            .O(N__43165),
            .I(N__43148));
    Span4Mux_h I__10045 (
            .O(N__43160),
            .I(N__43143));
    LocalMux I__10044 (
            .O(N__43157),
            .I(N__43143));
    LocalMux I__10043 (
            .O(N__43154),
            .I(N__43140));
    Span4Mux_h I__10042 (
            .O(N__43151),
            .I(N__43137));
    LocalMux I__10041 (
            .O(N__43148),
            .I(state_7_N_167_2));
    Odrv4 I__10040 (
            .O(N__43143),
            .I(state_7_N_167_2));
    Odrv12 I__10039 (
            .O(N__43140),
            .I(state_7_N_167_2));
    Odrv4 I__10038 (
            .O(N__43137),
            .I(state_7_N_167_2));
    InMux I__10037 (
            .O(N__43128),
            .I(N__43125));
    LocalMux I__10036 (
            .O(N__43125),
            .I(N__43122));
    Odrv4 I__10035 (
            .O(N__43122),
            .I(n26));
    CascadeMux I__10034 (
            .O(N__43119),
            .I(N__43116));
    InMux I__10033 (
            .O(N__43116),
            .I(N__43112));
    InMux I__10032 (
            .O(N__43115),
            .I(N__43109));
    LocalMux I__10031 (
            .O(N__43112),
            .I(counter_4));
    LocalMux I__10030 (
            .O(N__43109),
            .I(counter_4));
    InMux I__10029 (
            .O(N__43104),
            .I(N__43100));
    InMux I__10028 (
            .O(N__43103),
            .I(N__43097));
    LocalMux I__10027 (
            .O(N__43100),
            .I(counter_5));
    LocalMux I__10026 (
            .O(N__43097),
            .I(counter_5));
    CascadeMux I__10025 (
            .O(N__43092),
            .I(N__43088));
    CascadeMux I__10024 (
            .O(N__43091),
            .I(N__43085));
    InMux I__10023 (
            .O(N__43088),
            .I(N__43082));
    InMux I__10022 (
            .O(N__43085),
            .I(N__43079));
    LocalMux I__10021 (
            .O(N__43082),
            .I(counter_2));
    LocalMux I__10020 (
            .O(N__43079),
            .I(counter_2));
    InMux I__10019 (
            .O(N__43074),
            .I(N__43070));
    InMux I__10018 (
            .O(N__43073),
            .I(N__43067));
    LocalMux I__10017 (
            .O(N__43070),
            .I(counter_3));
    LocalMux I__10016 (
            .O(N__43067),
            .I(counter_3));
    InMux I__10015 (
            .O(N__43062),
            .I(N__43059));
    LocalMux I__10014 (
            .O(N__43059),
            .I(n14));
    IoInMux I__10013 (
            .O(N__43056),
            .I(N__43053));
    LocalMux I__10012 (
            .O(N__43053),
            .I(N__43050));
    Span12Mux_s5_h I__10011 (
            .O(N__43050),
            .I(N__43047));
    Span12Mux_h I__10010 (
            .O(N__43047),
            .I(N__43044));
    Span12Mux_v I__10009 (
            .O(N__43044),
            .I(N__43039));
    InMux I__10008 (
            .O(N__43043),
            .I(N__43034));
    InMux I__10007 (
            .O(N__43042),
            .I(N__43034));
    Odrv12 I__10006 (
            .O(N__43039),
            .I(pin_out_11));
    LocalMux I__10005 (
            .O(N__43034),
            .I(pin_out_11));
    CascadeMux I__10004 (
            .O(N__43029),
            .I(n7_adj_827_cascade_));
    IoInMux I__10003 (
            .O(N__43026),
            .I(N__43023));
    LocalMux I__10002 (
            .O(N__43023),
            .I(N__43020));
    Span4Mux_s3_v I__10001 (
            .O(N__43020),
            .I(N__43017));
    Sp12to4 I__10000 (
            .O(N__43017),
            .I(N__43014));
    Span12Mux_h I__9999 (
            .O(N__43014),
            .I(N__43011));
    Span12Mux_v I__9998 (
            .O(N__43011),
            .I(N__43006));
    InMux I__9997 (
            .O(N__43010),
            .I(N__43001));
    InMux I__9996 (
            .O(N__43009),
            .I(N__43001));
    Odrv12 I__9995 (
            .O(N__43006),
            .I(pin_out_10));
    LocalMux I__9994 (
            .O(N__43001),
            .I(pin_out_10));
    CascadeMux I__9993 (
            .O(N__42996),
            .I(n9675_cascade_));
    CascadeMux I__9992 (
            .O(N__42993),
            .I(n7_adj_823_cascade_));
    IoInMux I__9991 (
            .O(N__42990),
            .I(N__42987));
    LocalMux I__9990 (
            .O(N__42987),
            .I(N__42984));
    IoSpan4Mux I__9989 (
            .O(N__42984),
            .I(N__42981));
    Sp12to4 I__9988 (
            .O(N__42981),
            .I(N__42978));
    Span12Mux_v I__9987 (
            .O(N__42978),
            .I(N__42974));
    InMux I__9986 (
            .O(N__42977),
            .I(N__42971));
    Odrv12 I__9985 (
            .O(N__42974),
            .I(pin_oe_19));
    LocalMux I__9984 (
            .O(N__42971),
            .I(pin_oe_19));
    IoInMux I__9983 (
            .O(N__42966),
            .I(N__42963));
    LocalMux I__9982 (
            .O(N__42963),
            .I(N__42960));
    IoSpan4Mux I__9981 (
            .O(N__42960),
            .I(N__42957));
    Span4Mux_s3_h I__9980 (
            .O(N__42957),
            .I(N__42954));
    Sp12to4 I__9979 (
            .O(N__42954),
            .I(N__42951));
    Span12Mux_v I__9978 (
            .O(N__42951),
            .I(N__42947));
    InMux I__9977 (
            .O(N__42950),
            .I(N__42943));
    Span12Mux_h I__9976 (
            .O(N__42947),
            .I(N__42940));
    InMux I__9975 (
            .O(N__42946),
            .I(N__42937));
    LocalMux I__9974 (
            .O(N__42943),
            .I(N__42934));
    Odrv12 I__9973 (
            .O(N__42940),
            .I(pin_out_7));
    LocalMux I__9972 (
            .O(N__42937),
            .I(pin_out_7));
    Odrv4 I__9971 (
            .O(N__42934),
            .I(pin_out_7));
    IoInMux I__9970 (
            .O(N__42927),
            .I(N__42924));
    LocalMux I__9969 (
            .O(N__42924),
            .I(N__42921));
    Span4Mux_s3_h I__9968 (
            .O(N__42921),
            .I(N__42918));
    Span4Mux_v I__9967 (
            .O(N__42918),
            .I(N__42915));
    Span4Mux_v I__9966 (
            .O(N__42915),
            .I(N__42912));
    Sp12to4 I__9965 (
            .O(N__42912),
            .I(N__42909));
    Span12Mux_h I__9964 (
            .O(N__42909),
            .I(N__42904));
    InMux I__9963 (
            .O(N__42908),
            .I(N__42899));
    InMux I__9962 (
            .O(N__42907),
            .I(N__42899));
    Odrv12 I__9961 (
            .O(N__42904),
            .I(pin_out_6));
    LocalMux I__9960 (
            .O(N__42899),
            .I(pin_out_6));
    InMux I__9959 (
            .O(N__42894),
            .I(N__42891));
    LocalMux I__9958 (
            .O(N__42891),
            .I(n13358));
    InMux I__9957 (
            .O(N__42888),
            .I(N__42884));
    InMux I__9956 (
            .O(N__42887),
            .I(N__42881));
    LocalMux I__9955 (
            .O(N__42884),
            .I(N__42869));
    LocalMux I__9954 (
            .O(N__42881),
            .I(N__42869));
    InMux I__9953 (
            .O(N__42880),
            .I(N__42862));
    InMux I__9952 (
            .O(N__42879),
            .I(N__42862));
    InMux I__9951 (
            .O(N__42878),
            .I(N__42862));
    InMux I__9950 (
            .O(N__42877),
            .I(N__42853));
    InMux I__9949 (
            .O(N__42876),
            .I(N__42853));
    InMux I__9948 (
            .O(N__42875),
            .I(N__42853));
    InMux I__9947 (
            .O(N__42874),
            .I(N__42853));
    Span4Mux_v I__9946 (
            .O(N__42869),
            .I(N__42850));
    LocalMux I__9945 (
            .O(N__42862),
            .I(n3762));
    LocalMux I__9944 (
            .O(N__42853),
            .I(n3762));
    Odrv4 I__9943 (
            .O(N__42850),
            .I(n3762));
    InMux I__9942 (
            .O(N__42843),
            .I(N__42840));
    LocalMux I__9941 (
            .O(N__42840),
            .I(N__42837));
    Odrv4 I__9940 (
            .O(N__42837),
            .I(n11964));
    IoInMux I__9939 (
            .O(N__42834),
            .I(N__42831));
    LocalMux I__9938 (
            .O(N__42831),
            .I(N__42828));
    IoSpan4Mux I__9937 (
            .O(N__42828),
            .I(N__42825));
    Span4Mux_s0_h I__9936 (
            .O(N__42825),
            .I(N__42822));
    Sp12to4 I__9935 (
            .O(N__42822),
            .I(N__42819));
    Span12Mux_h I__9934 (
            .O(N__42819),
            .I(N__42815));
    InMux I__9933 (
            .O(N__42818),
            .I(N__42812));
    Odrv12 I__9932 (
            .O(N__42815),
            .I(pin_oe_16));
    LocalMux I__9931 (
            .O(N__42812),
            .I(pin_oe_16));
    InMux I__9930 (
            .O(N__42807),
            .I(N__42804));
    LocalMux I__9929 (
            .O(N__42804),
            .I(n11820));
    CascadeMux I__9928 (
            .O(N__42801),
            .I(N__42798));
    InMux I__9927 (
            .O(N__42798),
            .I(N__42794));
    InMux I__9926 (
            .O(N__42797),
            .I(N__42791));
    LocalMux I__9925 (
            .O(N__42794),
            .I(counter_7));
    LocalMux I__9924 (
            .O(N__42791),
            .I(counter_7));
    InMux I__9923 (
            .O(N__42786),
            .I(N__42782));
    InMux I__9922 (
            .O(N__42785),
            .I(N__42779));
    LocalMux I__9921 (
            .O(N__42782),
            .I(N__42776));
    LocalMux I__9920 (
            .O(N__42779),
            .I(counter_0));
    Odrv4 I__9919 (
            .O(N__42776),
            .I(counter_0));
    CascadeMux I__9918 (
            .O(N__42771),
            .I(N__42768));
    InMux I__9917 (
            .O(N__42768),
            .I(N__42764));
    InMux I__9916 (
            .O(N__42767),
            .I(N__42761));
    LocalMux I__9915 (
            .O(N__42764),
            .I(counter_6));
    LocalMux I__9914 (
            .O(N__42761),
            .I(counter_6));
    InMux I__9913 (
            .O(N__42756),
            .I(N__42752));
    InMux I__9912 (
            .O(N__42755),
            .I(N__42749));
    LocalMux I__9911 (
            .O(N__42752),
            .I(counter_1));
    LocalMux I__9910 (
            .O(N__42749),
            .I(counter_1));
    CascadeMux I__9909 (
            .O(N__42744),
            .I(n10_cascade_));
    CascadeMux I__9908 (
            .O(N__42741),
            .I(n9_adj_824_cascade_));
    CascadeMux I__9907 (
            .O(N__42738),
            .I(n8_adj_822_cascade_));
    IoInMux I__9906 (
            .O(N__42735),
            .I(N__42732));
    LocalMux I__9905 (
            .O(N__42732),
            .I(N__42729));
    Span12Mux_s5_h I__9904 (
            .O(N__42729),
            .I(N__42725));
    InMux I__9903 (
            .O(N__42728),
            .I(N__42721));
    Span12Mux_v I__9902 (
            .O(N__42725),
            .I(N__42718));
    InMux I__9901 (
            .O(N__42724),
            .I(N__42715));
    LocalMux I__9900 (
            .O(N__42721),
            .I(N__42712));
    Odrv12 I__9899 (
            .O(N__42718),
            .I(pin_out_5));
    LocalMux I__9898 (
            .O(N__42715),
            .I(pin_out_5));
    Odrv4 I__9897 (
            .O(N__42712),
            .I(pin_out_5));
    IoInMux I__9896 (
            .O(N__42705),
            .I(N__42702));
    LocalMux I__9895 (
            .O(N__42702),
            .I(N__42699));
    Span12Mux_s4_h I__9894 (
            .O(N__42699),
            .I(N__42695));
    InMux I__9893 (
            .O(N__42698),
            .I(N__42691));
    Span12Mux_v I__9892 (
            .O(N__42695),
            .I(N__42688));
    InMux I__9891 (
            .O(N__42694),
            .I(N__42685));
    LocalMux I__9890 (
            .O(N__42691),
            .I(N__42682));
    Odrv12 I__9889 (
            .O(N__42688),
            .I(pin_out_4));
    LocalMux I__9888 (
            .O(N__42685),
            .I(pin_out_4));
    Odrv4 I__9887 (
            .O(N__42682),
            .I(pin_out_4));
    CascadeMux I__9886 (
            .O(N__42675),
            .I(n13357_cascade_));
    InMux I__9885 (
            .O(N__42672),
            .I(N__42669));
    LocalMux I__9884 (
            .O(N__42669),
            .I(n13625));
    CascadeMux I__9883 (
            .O(N__42666),
            .I(n6_adj_810_cascade_));
    InMux I__9882 (
            .O(N__42663),
            .I(N__42660));
    LocalMux I__9881 (
            .O(N__42660),
            .I(N__42657));
    Span4Mux_h I__9880 (
            .O(N__42657),
            .I(N__42654));
    Span4Mux_v I__9879 (
            .O(N__42654),
            .I(N__42651));
    Odrv4 I__9878 (
            .O(N__42651),
            .I(n11874));
    CascadeMux I__9877 (
            .O(N__42648),
            .I(N__42645));
    InMux I__9876 (
            .O(N__42645),
            .I(N__42642));
    LocalMux I__9875 (
            .O(N__42642),
            .I(n11823));
    InMux I__9874 (
            .O(N__42639),
            .I(N__42636));
    LocalMux I__9873 (
            .O(N__42636),
            .I(N__42632));
    InMux I__9872 (
            .O(N__42635),
            .I(N__42629));
    Span4Mux_s3_h I__9871 (
            .O(N__42632),
            .I(N__42622));
    LocalMux I__9870 (
            .O(N__42629),
            .I(N__42622));
    InMux I__9869 (
            .O(N__42628),
            .I(N__42619));
    InMux I__9868 (
            .O(N__42627),
            .I(N__42616));
    Span4Mux_v I__9867 (
            .O(N__42622),
            .I(N__42610));
    LocalMux I__9866 (
            .O(N__42619),
            .I(N__42605));
    LocalMux I__9865 (
            .O(N__42616),
            .I(N__42605));
    InMux I__9864 (
            .O(N__42615),
            .I(N__42600));
    InMux I__9863 (
            .O(N__42614),
            .I(N__42595));
    InMux I__9862 (
            .O(N__42613),
            .I(N__42595));
    Span4Mux_h I__9861 (
            .O(N__42610),
            .I(N__42592));
    Span4Mux_v I__9860 (
            .O(N__42605),
            .I(N__42589));
    InMux I__9859 (
            .O(N__42604),
            .I(N__42584));
    InMux I__9858 (
            .O(N__42603),
            .I(N__42579));
    LocalMux I__9857 (
            .O(N__42600),
            .I(N__42575));
    LocalMux I__9856 (
            .O(N__42595),
            .I(N__42572));
    Span4Mux_h I__9855 (
            .O(N__42592),
            .I(N__42569));
    Span4Mux_h I__9854 (
            .O(N__42589),
            .I(N__42566));
    InMux I__9853 (
            .O(N__42588),
            .I(N__42561));
    InMux I__9852 (
            .O(N__42587),
            .I(N__42561));
    LocalMux I__9851 (
            .O(N__42584),
            .I(N__42558));
    InMux I__9850 (
            .O(N__42583),
            .I(N__42553));
    InMux I__9849 (
            .O(N__42582),
            .I(N__42553));
    LocalMux I__9848 (
            .O(N__42579),
            .I(N__42550));
    InMux I__9847 (
            .O(N__42578),
            .I(N__42547));
    Span4Mux_v I__9846 (
            .O(N__42575),
            .I(N__42542));
    Span4Mux_v I__9845 (
            .O(N__42572),
            .I(N__42542));
    Span4Mux_h I__9844 (
            .O(N__42569),
            .I(N__42539));
    Span4Mux_h I__9843 (
            .O(N__42566),
            .I(N__42536));
    LocalMux I__9842 (
            .O(N__42561),
            .I(n7));
    Odrv12 I__9841 (
            .O(N__42558),
            .I(n7));
    LocalMux I__9840 (
            .O(N__42553),
            .I(n7));
    Odrv4 I__9839 (
            .O(N__42550),
            .I(n7));
    LocalMux I__9838 (
            .O(N__42547),
            .I(n7));
    Odrv4 I__9837 (
            .O(N__42542),
            .I(n7));
    Odrv4 I__9836 (
            .O(N__42539),
            .I(n7));
    Odrv4 I__9835 (
            .O(N__42536),
            .I(n7));
    InMux I__9834 (
            .O(N__42519),
            .I(n10576));
    InMux I__9833 (
            .O(N__42516),
            .I(n10577));
    InMux I__9832 (
            .O(N__42513),
            .I(n10578));
    InMux I__9831 (
            .O(N__42510),
            .I(N__42506));
    InMux I__9830 (
            .O(N__42509),
            .I(N__42503));
    LocalMux I__9829 (
            .O(N__42506),
            .I(current_pin_5));
    LocalMux I__9828 (
            .O(N__42503),
            .I(current_pin_5));
    InMux I__9827 (
            .O(N__42498),
            .I(n10579));
    InMux I__9826 (
            .O(N__42495),
            .I(N__42491));
    InMux I__9825 (
            .O(N__42494),
            .I(N__42488));
    LocalMux I__9824 (
            .O(N__42491),
            .I(current_pin_6));
    LocalMux I__9823 (
            .O(N__42488),
            .I(current_pin_6));
    InMux I__9822 (
            .O(N__42483),
            .I(n10580));
    InMux I__9821 (
            .O(N__42480),
            .I(n10581));
    InMux I__9820 (
            .O(N__42477),
            .I(N__42473));
    InMux I__9819 (
            .O(N__42476),
            .I(N__42470));
    LocalMux I__9818 (
            .O(N__42473),
            .I(current_pin_7));
    LocalMux I__9817 (
            .O(N__42470),
            .I(current_pin_7));
    SRMux I__9816 (
            .O(N__42465),
            .I(N__42462));
    LocalMux I__9815 (
            .O(N__42462),
            .I(N__42459));
    Odrv4 I__9814 (
            .O(N__42459),
            .I(n7985));
    CEMux I__9813 (
            .O(N__42456),
            .I(N__42452));
    InMux I__9812 (
            .O(N__42455),
            .I(N__42449));
    LocalMux I__9811 (
            .O(N__42452),
            .I(n7635));
    LocalMux I__9810 (
            .O(N__42449),
            .I(n7635));
    InMux I__9809 (
            .O(N__42444),
            .I(n10703));
    InMux I__9808 (
            .O(N__42441),
            .I(n10704));
    InMux I__9807 (
            .O(N__42438),
            .I(n10705));
    CascadeMux I__9806 (
            .O(N__42435),
            .I(N__42428));
    CascadeMux I__9805 (
            .O(N__42434),
            .I(N__42424));
    CascadeMux I__9804 (
            .O(N__42433),
            .I(N__42420));
    InMux I__9803 (
            .O(N__42432),
            .I(N__42405));
    InMux I__9802 (
            .O(N__42431),
            .I(N__42405));
    InMux I__9801 (
            .O(N__42428),
            .I(N__42405));
    InMux I__9800 (
            .O(N__42427),
            .I(N__42405));
    InMux I__9799 (
            .O(N__42424),
            .I(N__42405));
    InMux I__9798 (
            .O(N__42423),
            .I(N__42405));
    InMux I__9797 (
            .O(N__42420),
            .I(N__42405));
    LocalMux I__9796 (
            .O(N__42405),
            .I(n13603));
    InMux I__9795 (
            .O(N__42402),
            .I(n10706));
    CEMux I__9794 (
            .O(N__42399),
            .I(N__42395));
    CEMux I__9793 (
            .O(N__42398),
            .I(N__42392));
    LocalMux I__9792 (
            .O(N__42395),
            .I(N__42387));
    LocalMux I__9791 (
            .O(N__42392),
            .I(N__42387));
    Span4Mux_v I__9790 (
            .O(N__42387),
            .I(N__42384));
    Odrv4 I__9789 (
            .O(N__42384),
            .I(n7681));
    InMux I__9788 (
            .O(N__42381),
            .I(N__42378));
    LocalMux I__9787 (
            .O(N__42378),
            .I(N__42375));
    Span4Mux_h I__9786 (
            .O(N__42375),
            .I(N__42372));
    Odrv4 I__9785 (
            .O(N__42372),
            .I(n11824));
    InMux I__9784 (
            .O(N__42369),
            .I(bfn_17_17_0_));
    InMux I__9783 (
            .O(N__42366),
            .I(n10575));
    CascadeMux I__9782 (
            .O(N__42363),
            .I(N__42359));
    CascadeMux I__9781 (
            .O(N__42362),
            .I(N__42356));
    InMux I__9780 (
            .O(N__42359),
            .I(N__42353));
    InMux I__9779 (
            .O(N__42356),
            .I(N__42350));
    LocalMux I__9778 (
            .O(N__42353),
            .I(\nx.n2491 ));
    LocalMux I__9777 (
            .O(N__42350),
            .I(\nx.n2491 ));
    InMux I__9776 (
            .O(N__42345),
            .I(N__42342));
    LocalMux I__9775 (
            .O(N__42342),
            .I(\nx.n2558 ));
    InMux I__9774 (
            .O(N__42339),
            .I(\nx.n10956 ));
    CascadeMux I__9773 (
            .O(N__42336),
            .I(N__42333));
    InMux I__9772 (
            .O(N__42333),
            .I(N__42329));
    CascadeMux I__9771 (
            .O(N__42332),
            .I(N__42326));
    LocalMux I__9770 (
            .O(N__42329),
            .I(N__42323));
    InMux I__9769 (
            .O(N__42326),
            .I(N__42320));
    Span4Mux_v I__9768 (
            .O(N__42323),
            .I(N__42317));
    LocalMux I__9767 (
            .O(N__42320),
            .I(\nx.n2490 ));
    Odrv4 I__9766 (
            .O(N__42317),
            .I(\nx.n2490 ));
    InMux I__9765 (
            .O(N__42312),
            .I(N__42309));
    LocalMux I__9764 (
            .O(N__42309),
            .I(N__42306));
    Odrv4 I__9763 (
            .O(N__42306),
            .I(\nx.n2557 ));
    InMux I__9762 (
            .O(N__42303),
            .I(\nx.n10957 ));
    CascadeMux I__9761 (
            .O(N__42300),
            .I(N__42290));
    CascadeMux I__9760 (
            .O(N__42299),
            .I(N__42284));
    CascadeMux I__9759 (
            .O(N__42298),
            .I(N__42276));
    CascadeMux I__9758 (
            .O(N__42297),
            .I(N__42271));
    CascadeMux I__9757 (
            .O(N__42296),
            .I(N__42264));
    CascadeMux I__9756 (
            .O(N__42295),
            .I(N__42259));
    InMux I__9755 (
            .O(N__42294),
            .I(N__42244));
    InMux I__9754 (
            .O(N__42293),
            .I(N__42244));
    InMux I__9753 (
            .O(N__42290),
            .I(N__42244));
    InMux I__9752 (
            .O(N__42289),
            .I(N__42239));
    InMux I__9751 (
            .O(N__42288),
            .I(N__42239));
    InMux I__9750 (
            .O(N__42287),
            .I(N__42230));
    InMux I__9749 (
            .O(N__42284),
            .I(N__42230));
    InMux I__9748 (
            .O(N__42283),
            .I(N__42230));
    InMux I__9747 (
            .O(N__42282),
            .I(N__42230));
    CascadeMux I__9746 (
            .O(N__42281),
            .I(N__42226));
    InMux I__9745 (
            .O(N__42280),
            .I(N__42188));
    InMux I__9744 (
            .O(N__42279),
            .I(N__42188));
    InMux I__9743 (
            .O(N__42276),
            .I(N__42176));
    InMux I__9742 (
            .O(N__42275),
            .I(N__42176));
    InMux I__9741 (
            .O(N__42274),
            .I(N__42176));
    InMux I__9740 (
            .O(N__42271),
            .I(N__42176));
    InMux I__9739 (
            .O(N__42270),
            .I(N__42176));
    InMux I__9738 (
            .O(N__42269),
            .I(N__42163));
    InMux I__9737 (
            .O(N__42268),
            .I(N__42163));
    InMux I__9736 (
            .O(N__42267),
            .I(N__42154));
    InMux I__9735 (
            .O(N__42264),
            .I(N__42154));
    InMux I__9734 (
            .O(N__42263),
            .I(N__42154));
    InMux I__9733 (
            .O(N__42262),
            .I(N__42154));
    InMux I__9732 (
            .O(N__42259),
            .I(N__42145));
    InMux I__9731 (
            .O(N__42258),
            .I(N__42145));
    InMux I__9730 (
            .O(N__42257),
            .I(N__42145));
    InMux I__9729 (
            .O(N__42256),
            .I(N__42145));
    InMux I__9728 (
            .O(N__42255),
            .I(N__42142));
    InMux I__9727 (
            .O(N__42254),
            .I(N__42129));
    InMux I__9726 (
            .O(N__42253),
            .I(N__42129));
    InMux I__9725 (
            .O(N__42252),
            .I(N__42129));
    InMux I__9724 (
            .O(N__42251),
            .I(N__42129));
    LocalMux I__9723 (
            .O(N__42244),
            .I(N__42113));
    LocalMux I__9722 (
            .O(N__42239),
            .I(N__42113));
    LocalMux I__9721 (
            .O(N__42230),
            .I(N__42113));
    InMux I__9720 (
            .O(N__42229),
            .I(N__42110));
    InMux I__9719 (
            .O(N__42226),
            .I(N__42105));
    InMux I__9718 (
            .O(N__42225),
            .I(N__42105));
    InMux I__9717 (
            .O(N__42224),
            .I(N__42102));
    InMux I__9716 (
            .O(N__42223),
            .I(N__42099));
    InMux I__9715 (
            .O(N__42222),
            .I(N__42077));
    InMux I__9714 (
            .O(N__42221),
            .I(N__42077));
    InMux I__9713 (
            .O(N__42220),
            .I(N__42077));
    InMux I__9712 (
            .O(N__42219),
            .I(N__42077));
    InMux I__9711 (
            .O(N__42218),
            .I(N__42072));
    InMux I__9710 (
            .O(N__42217),
            .I(N__42072));
    InMux I__9709 (
            .O(N__42216),
            .I(N__42068));
    InMux I__9708 (
            .O(N__42215),
            .I(N__42044));
    InMux I__9707 (
            .O(N__42214),
            .I(N__42034));
    InMux I__9706 (
            .O(N__42213),
            .I(N__42034));
    InMux I__9705 (
            .O(N__42212),
            .I(N__42034));
    CascadeMux I__9704 (
            .O(N__42211),
            .I(N__42027));
    CascadeMux I__9703 (
            .O(N__42210),
            .I(N__42016));
    CascadeMux I__9702 (
            .O(N__42209),
            .I(N__42006));
    InMux I__9701 (
            .O(N__42208),
            .I(N__41988));
    InMux I__9700 (
            .O(N__42207),
            .I(N__41988));
    InMux I__9699 (
            .O(N__42206),
            .I(N__41988));
    InMux I__9698 (
            .O(N__42205),
            .I(N__41988));
    InMux I__9697 (
            .O(N__42204),
            .I(N__41979));
    InMux I__9696 (
            .O(N__42203),
            .I(N__41979));
    InMux I__9695 (
            .O(N__42202),
            .I(N__41979));
    InMux I__9694 (
            .O(N__42201),
            .I(N__41979));
    InMux I__9693 (
            .O(N__42200),
            .I(N__41969));
    InMux I__9692 (
            .O(N__42199),
            .I(N__41969));
    InMux I__9691 (
            .O(N__42198),
            .I(N__41960));
    InMux I__9690 (
            .O(N__42197),
            .I(N__41953));
    InMux I__9689 (
            .O(N__42196),
            .I(N__41953));
    InMux I__9688 (
            .O(N__42195),
            .I(N__41953));
    InMux I__9687 (
            .O(N__42194),
            .I(N__41948));
    InMux I__9686 (
            .O(N__42193),
            .I(N__41948));
    LocalMux I__9685 (
            .O(N__42188),
            .I(N__41945));
    CascadeMux I__9684 (
            .O(N__42187),
            .I(N__41940));
    LocalMux I__9683 (
            .O(N__42176),
            .I(N__41932));
    InMux I__9682 (
            .O(N__42175),
            .I(N__41923));
    InMux I__9681 (
            .O(N__42174),
            .I(N__41923));
    InMux I__9680 (
            .O(N__42173),
            .I(N__41923));
    InMux I__9679 (
            .O(N__42172),
            .I(N__41923));
    InMux I__9678 (
            .O(N__42171),
            .I(N__41914));
    InMux I__9677 (
            .O(N__42170),
            .I(N__41914));
    InMux I__9676 (
            .O(N__42169),
            .I(N__41914));
    InMux I__9675 (
            .O(N__42168),
            .I(N__41914));
    LocalMux I__9674 (
            .O(N__42163),
            .I(N__41905));
    LocalMux I__9673 (
            .O(N__42154),
            .I(N__41905));
    LocalMux I__9672 (
            .O(N__42145),
            .I(N__41905));
    LocalMux I__9671 (
            .O(N__42142),
            .I(N__41905));
    InMux I__9670 (
            .O(N__42141),
            .I(N__41896));
    InMux I__9669 (
            .O(N__42140),
            .I(N__41896));
    InMux I__9668 (
            .O(N__42139),
            .I(N__41896));
    InMux I__9667 (
            .O(N__42138),
            .I(N__41896));
    LocalMux I__9666 (
            .O(N__42129),
            .I(N__41893));
    InMux I__9665 (
            .O(N__42128),
            .I(N__41886));
    InMux I__9664 (
            .O(N__42127),
            .I(N__41886));
    InMux I__9663 (
            .O(N__42126),
            .I(N__41886));
    InMux I__9662 (
            .O(N__42125),
            .I(N__41879));
    InMux I__9661 (
            .O(N__42124),
            .I(N__41879));
    InMux I__9660 (
            .O(N__42123),
            .I(N__41879));
    CascadeMux I__9659 (
            .O(N__42122),
            .I(N__41876));
    CascadeMux I__9658 (
            .O(N__42121),
            .I(N__41872));
    CascadeMux I__9657 (
            .O(N__42120),
            .I(N__41869));
    Span4Mux_v I__9656 (
            .O(N__42113),
            .I(N__41855));
    LocalMux I__9655 (
            .O(N__42110),
            .I(N__41855));
    LocalMux I__9654 (
            .O(N__42105),
            .I(N__41855));
    LocalMux I__9653 (
            .O(N__42102),
            .I(N__41850));
    LocalMux I__9652 (
            .O(N__42099),
            .I(N__41850));
    InMux I__9651 (
            .O(N__42098),
            .I(N__41843));
    InMux I__9650 (
            .O(N__42097),
            .I(N__41843));
    InMux I__9649 (
            .O(N__42096),
            .I(N__41843));
    InMux I__9648 (
            .O(N__42095),
            .I(N__41836));
    InMux I__9647 (
            .O(N__42094),
            .I(N__41836));
    InMux I__9646 (
            .O(N__42093),
            .I(N__41836));
    InMux I__9645 (
            .O(N__42092),
            .I(N__41827));
    InMux I__9644 (
            .O(N__42091),
            .I(N__41827));
    InMux I__9643 (
            .O(N__42090),
            .I(N__41827));
    InMux I__9642 (
            .O(N__42089),
            .I(N__41827));
    InMux I__9641 (
            .O(N__42088),
            .I(N__41820));
    InMux I__9640 (
            .O(N__42087),
            .I(N__41820));
    InMux I__9639 (
            .O(N__42086),
            .I(N__41820));
    LocalMux I__9638 (
            .O(N__42077),
            .I(N__41815));
    LocalMux I__9637 (
            .O(N__42072),
            .I(N__41815));
    CascadeMux I__9636 (
            .O(N__42071),
            .I(N__41807));
    LocalMux I__9635 (
            .O(N__42068),
            .I(N__41802));
    InMux I__9634 (
            .O(N__42067),
            .I(N__41793));
    InMux I__9633 (
            .O(N__42066),
            .I(N__41793));
    InMux I__9632 (
            .O(N__42065),
            .I(N__41793));
    InMux I__9631 (
            .O(N__42064),
            .I(N__41793));
    InMux I__9630 (
            .O(N__42063),
            .I(N__41786));
    InMux I__9629 (
            .O(N__42062),
            .I(N__41786));
    InMux I__9628 (
            .O(N__42061),
            .I(N__41786));
    InMux I__9627 (
            .O(N__42060),
            .I(N__41783));
    InMux I__9626 (
            .O(N__42059),
            .I(N__41772));
    InMux I__9625 (
            .O(N__42058),
            .I(N__41772));
    InMux I__9624 (
            .O(N__42057),
            .I(N__41772));
    InMux I__9623 (
            .O(N__42056),
            .I(N__41772));
    InMux I__9622 (
            .O(N__42055),
            .I(N__41772));
    InMux I__9621 (
            .O(N__42054),
            .I(N__41763));
    InMux I__9620 (
            .O(N__42053),
            .I(N__41763));
    InMux I__9619 (
            .O(N__42052),
            .I(N__41763));
    InMux I__9618 (
            .O(N__42051),
            .I(N__41763));
    InMux I__9617 (
            .O(N__42050),
            .I(N__41754));
    InMux I__9616 (
            .O(N__42049),
            .I(N__41754));
    InMux I__9615 (
            .O(N__42048),
            .I(N__41754));
    InMux I__9614 (
            .O(N__42047),
            .I(N__41754));
    LocalMux I__9613 (
            .O(N__42044),
            .I(N__41739));
    InMux I__9612 (
            .O(N__42043),
            .I(N__41732));
    InMux I__9611 (
            .O(N__42042),
            .I(N__41732));
    InMux I__9610 (
            .O(N__42041),
            .I(N__41732));
    LocalMux I__9609 (
            .O(N__42034),
            .I(N__41729));
    InMux I__9608 (
            .O(N__42033),
            .I(N__41724));
    InMux I__9607 (
            .O(N__42032),
            .I(N__41724));
    InMux I__9606 (
            .O(N__42031),
            .I(N__41713));
    InMux I__9605 (
            .O(N__42030),
            .I(N__41713));
    InMux I__9604 (
            .O(N__42027),
            .I(N__41713));
    InMux I__9603 (
            .O(N__42026),
            .I(N__41713));
    InMux I__9602 (
            .O(N__42025),
            .I(N__41713));
    InMux I__9601 (
            .O(N__42024),
            .I(N__41704));
    InMux I__9600 (
            .O(N__42023),
            .I(N__41704));
    InMux I__9599 (
            .O(N__42022),
            .I(N__41704));
    InMux I__9598 (
            .O(N__42021),
            .I(N__41704));
    InMux I__9597 (
            .O(N__42020),
            .I(N__41695));
    InMux I__9596 (
            .O(N__42019),
            .I(N__41695));
    InMux I__9595 (
            .O(N__42016),
            .I(N__41695));
    InMux I__9594 (
            .O(N__42015),
            .I(N__41695));
    InMux I__9593 (
            .O(N__42014),
            .I(N__41688));
    InMux I__9592 (
            .O(N__42013),
            .I(N__41688));
    InMux I__9591 (
            .O(N__42012),
            .I(N__41688));
    InMux I__9590 (
            .O(N__42011),
            .I(N__41681));
    InMux I__9589 (
            .O(N__42010),
            .I(N__41681));
    InMux I__9588 (
            .O(N__42009),
            .I(N__41681));
    InMux I__9587 (
            .O(N__42006),
            .I(N__41672));
    InMux I__9586 (
            .O(N__42005),
            .I(N__41672));
    InMux I__9585 (
            .O(N__42004),
            .I(N__41672));
    InMux I__9584 (
            .O(N__42003),
            .I(N__41663));
    InMux I__9583 (
            .O(N__42002),
            .I(N__41663));
    InMux I__9582 (
            .O(N__42001),
            .I(N__41663));
    InMux I__9581 (
            .O(N__42000),
            .I(N__41663));
    InMux I__9580 (
            .O(N__41999),
            .I(N__41658));
    InMux I__9579 (
            .O(N__41998),
            .I(N__41658));
    CascadeMux I__9578 (
            .O(N__41997),
            .I(N__41649));
    LocalMux I__9577 (
            .O(N__41988),
            .I(N__41633));
    LocalMux I__9576 (
            .O(N__41979),
            .I(N__41633));
    InMux I__9575 (
            .O(N__41978),
            .I(N__41620));
    InMux I__9574 (
            .O(N__41977),
            .I(N__41620));
    InMux I__9573 (
            .O(N__41976),
            .I(N__41620));
    CascadeMux I__9572 (
            .O(N__41975),
            .I(N__41601));
    CascadeMux I__9571 (
            .O(N__41974),
            .I(N__41593));
    LocalMux I__9570 (
            .O(N__41969),
            .I(N__41586));
    InMux I__9569 (
            .O(N__41968),
            .I(N__41579));
    InMux I__9568 (
            .O(N__41967),
            .I(N__41579));
    InMux I__9567 (
            .O(N__41966),
            .I(N__41579));
    CascadeMux I__9566 (
            .O(N__41965),
            .I(N__41574));
    CascadeMux I__9565 (
            .O(N__41964),
            .I(N__41569));
    CascadeMux I__9564 (
            .O(N__41963),
            .I(N__41562));
    LocalMux I__9563 (
            .O(N__41960),
            .I(N__41552));
    LocalMux I__9562 (
            .O(N__41953),
            .I(N__41552));
    LocalMux I__9561 (
            .O(N__41948),
            .I(N__41552));
    Span4Mux_v I__9560 (
            .O(N__41945),
            .I(N__41549));
    InMux I__9559 (
            .O(N__41944),
            .I(N__41540));
    InMux I__9558 (
            .O(N__41943),
            .I(N__41540));
    InMux I__9557 (
            .O(N__41940),
            .I(N__41540));
    InMux I__9556 (
            .O(N__41939),
            .I(N__41540));
    InMux I__9555 (
            .O(N__41938),
            .I(N__41531));
    InMux I__9554 (
            .O(N__41937),
            .I(N__41531));
    InMux I__9553 (
            .O(N__41936),
            .I(N__41531));
    InMux I__9552 (
            .O(N__41935),
            .I(N__41531));
    Span4Mux_v I__9551 (
            .O(N__41932),
            .I(N__41524));
    LocalMux I__9550 (
            .O(N__41923),
            .I(N__41524));
    LocalMux I__9549 (
            .O(N__41914),
            .I(N__41524));
    Span4Mux_v I__9548 (
            .O(N__41905),
            .I(N__41519));
    LocalMux I__9547 (
            .O(N__41896),
            .I(N__41519));
    Span4Mux_v I__9546 (
            .O(N__41893),
            .I(N__41512));
    LocalMux I__9545 (
            .O(N__41886),
            .I(N__41512));
    LocalMux I__9544 (
            .O(N__41879),
            .I(N__41512));
    InMux I__9543 (
            .O(N__41876),
            .I(N__41509));
    InMux I__9542 (
            .O(N__41875),
            .I(N__41502));
    InMux I__9541 (
            .O(N__41872),
            .I(N__41502));
    InMux I__9540 (
            .O(N__41869),
            .I(N__41502));
    CascadeMux I__9539 (
            .O(N__41868),
            .I(N__41499));
    CascadeMux I__9538 (
            .O(N__41867),
            .I(N__41496));
    CascadeMux I__9537 (
            .O(N__41866),
            .I(N__41493));
    CascadeMux I__9536 (
            .O(N__41865),
            .I(N__41490));
    CascadeMux I__9535 (
            .O(N__41864),
            .I(N__41487));
    CascadeMux I__9534 (
            .O(N__41863),
            .I(N__41484));
    CascadeMux I__9533 (
            .O(N__41862),
            .I(N__41480));
    Span4Mux_v I__9532 (
            .O(N__41855),
            .I(N__41467));
    Span4Mux_v I__9531 (
            .O(N__41850),
            .I(N__41467));
    LocalMux I__9530 (
            .O(N__41843),
            .I(N__41462));
    LocalMux I__9529 (
            .O(N__41836),
            .I(N__41462));
    LocalMux I__9528 (
            .O(N__41827),
            .I(N__41457));
    LocalMux I__9527 (
            .O(N__41820),
            .I(N__41457));
    Span4Mux_v I__9526 (
            .O(N__41815),
            .I(N__41454));
    InMux I__9525 (
            .O(N__41814),
            .I(N__41445));
    InMux I__9524 (
            .O(N__41813),
            .I(N__41445));
    InMux I__9523 (
            .O(N__41812),
            .I(N__41445));
    InMux I__9522 (
            .O(N__41811),
            .I(N__41445));
    InMux I__9521 (
            .O(N__41810),
            .I(N__41436));
    InMux I__9520 (
            .O(N__41807),
            .I(N__41436));
    InMux I__9519 (
            .O(N__41806),
            .I(N__41436));
    InMux I__9518 (
            .O(N__41805),
            .I(N__41436));
    Span4Mux_v I__9517 (
            .O(N__41802),
            .I(N__41421));
    LocalMux I__9516 (
            .O(N__41793),
            .I(N__41421));
    LocalMux I__9515 (
            .O(N__41786),
            .I(N__41421));
    LocalMux I__9514 (
            .O(N__41783),
            .I(N__41421));
    LocalMux I__9513 (
            .O(N__41772),
            .I(N__41421));
    LocalMux I__9512 (
            .O(N__41763),
            .I(N__41421));
    LocalMux I__9511 (
            .O(N__41754),
            .I(N__41421));
    InMux I__9510 (
            .O(N__41753),
            .I(N__41414));
    InMux I__9509 (
            .O(N__41752),
            .I(N__41414));
    InMux I__9508 (
            .O(N__41751),
            .I(N__41414));
    InMux I__9507 (
            .O(N__41750),
            .I(N__41407));
    InMux I__9506 (
            .O(N__41749),
            .I(N__41407));
    InMux I__9505 (
            .O(N__41748),
            .I(N__41407));
    InMux I__9504 (
            .O(N__41747),
            .I(N__41400));
    InMux I__9503 (
            .O(N__41746),
            .I(N__41400));
    InMux I__9502 (
            .O(N__41745),
            .I(N__41400));
    InMux I__9501 (
            .O(N__41744),
            .I(N__41393));
    InMux I__9500 (
            .O(N__41743),
            .I(N__41393));
    InMux I__9499 (
            .O(N__41742),
            .I(N__41393));
    Span4Mux_v I__9498 (
            .O(N__41739),
            .I(N__41390));
    LocalMux I__9497 (
            .O(N__41732),
            .I(N__41387));
    Span4Mux_v I__9496 (
            .O(N__41729),
            .I(N__41372));
    LocalMux I__9495 (
            .O(N__41724),
            .I(N__41372));
    LocalMux I__9494 (
            .O(N__41713),
            .I(N__41372));
    LocalMux I__9493 (
            .O(N__41704),
            .I(N__41372));
    LocalMux I__9492 (
            .O(N__41695),
            .I(N__41372));
    LocalMux I__9491 (
            .O(N__41688),
            .I(N__41372));
    LocalMux I__9490 (
            .O(N__41681),
            .I(N__41372));
    InMux I__9489 (
            .O(N__41680),
            .I(N__41367));
    InMux I__9488 (
            .O(N__41679),
            .I(N__41367));
    LocalMux I__9487 (
            .O(N__41672),
            .I(N__41360));
    LocalMux I__9486 (
            .O(N__41663),
            .I(N__41360));
    LocalMux I__9485 (
            .O(N__41658),
            .I(N__41360));
    InMux I__9484 (
            .O(N__41657),
            .I(N__41353));
    InMux I__9483 (
            .O(N__41656),
            .I(N__41353));
    InMux I__9482 (
            .O(N__41655),
            .I(N__41353));
    InMux I__9481 (
            .O(N__41654),
            .I(N__41342));
    InMux I__9480 (
            .O(N__41653),
            .I(N__41342));
    InMux I__9479 (
            .O(N__41652),
            .I(N__41342));
    InMux I__9478 (
            .O(N__41649),
            .I(N__41342));
    InMux I__9477 (
            .O(N__41648),
            .I(N__41342));
    InMux I__9476 (
            .O(N__41647),
            .I(N__41333));
    InMux I__9475 (
            .O(N__41646),
            .I(N__41333));
    InMux I__9474 (
            .O(N__41645),
            .I(N__41333));
    InMux I__9473 (
            .O(N__41644),
            .I(N__41333));
    InMux I__9472 (
            .O(N__41643),
            .I(N__41324));
    InMux I__9471 (
            .O(N__41642),
            .I(N__41324));
    InMux I__9470 (
            .O(N__41641),
            .I(N__41324));
    InMux I__9469 (
            .O(N__41640),
            .I(N__41324));
    CascadeMux I__9468 (
            .O(N__41639),
            .I(N__41318));
    CascadeMux I__9467 (
            .O(N__41638),
            .I(N__41311));
    Span4Mux_v I__9466 (
            .O(N__41633),
            .I(N__41305));
    InMux I__9465 (
            .O(N__41632),
            .I(N__41298));
    InMux I__9464 (
            .O(N__41631),
            .I(N__41298));
    InMux I__9463 (
            .O(N__41630),
            .I(N__41298));
    InMux I__9462 (
            .O(N__41629),
            .I(N__41291));
    InMux I__9461 (
            .O(N__41628),
            .I(N__41291));
    InMux I__9460 (
            .O(N__41627),
            .I(N__41291));
    LocalMux I__9459 (
            .O(N__41620),
            .I(N__41288));
    InMux I__9458 (
            .O(N__41619),
            .I(N__41285));
    InMux I__9457 (
            .O(N__41618),
            .I(N__41278));
    InMux I__9456 (
            .O(N__41617),
            .I(N__41278));
    InMux I__9455 (
            .O(N__41616),
            .I(N__41278));
    InMux I__9454 (
            .O(N__41615),
            .I(N__41271));
    InMux I__9453 (
            .O(N__41614),
            .I(N__41271));
    InMux I__9452 (
            .O(N__41613),
            .I(N__41271));
    InMux I__9451 (
            .O(N__41612),
            .I(N__41264));
    InMux I__9450 (
            .O(N__41611),
            .I(N__41264));
    InMux I__9449 (
            .O(N__41610),
            .I(N__41264));
    InMux I__9448 (
            .O(N__41609),
            .I(N__41259));
    InMux I__9447 (
            .O(N__41608),
            .I(N__41259));
    InMux I__9446 (
            .O(N__41607),
            .I(N__41252));
    InMux I__9445 (
            .O(N__41606),
            .I(N__41252));
    InMux I__9444 (
            .O(N__41605),
            .I(N__41252));
    InMux I__9443 (
            .O(N__41604),
            .I(N__41241));
    InMux I__9442 (
            .O(N__41601),
            .I(N__41241));
    InMux I__9441 (
            .O(N__41600),
            .I(N__41241));
    InMux I__9440 (
            .O(N__41599),
            .I(N__41241));
    InMux I__9439 (
            .O(N__41598),
            .I(N__41241));
    InMux I__9438 (
            .O(N__41597),
            .I(N__41232));
    InMux I__9437 (
            .O(N__41596),
            .I(N__41232));
    InMux I__9436 (
            .O(N__41593),
            .I(N__41232));
    InMux I__9435 (
            .O(N__41592),
            .I(N__41232));
    InMux I__9434 (
            .O(N__41591),
            .I(N__41227));
    InMux I__9433 (
            .O(N__41590),
            .I(N__41227));
    InMux I__9432 (
            .O(N__41589),
            .I(N__41224));
    Span4Mux_v I__9431 (
            .O(N__41586),
            .I(N__41219));
    LocalMux I__9430 (
            .O(N__41579),
            .I(N__41219));
    InMux I__9429 (
            .O(N__41578),
            .I(N__41210));
    InMux I__9428 (
            .O(N__41577),
            .I(N__41210));
    InMux I__9427 (
            .O(N__41574),
            .I(N__41210));
    InMux I__9426 (
            .O(N__41573),
            .I(N__41210));
    InMux I__9425 (
            .O(N__41572),
            .I(N__41201));
    InMux I__9424 (
            .O(N__41569),
            .I(N__41201));
    InMux I__9423 (
            .O(N__41568),
            .I(N__41201));
    InMux I__9422 (
            .O(N__41567),
            .I(N__41201));
    InMux I__9421 (
            .O(N__41566),
            .I(N__41192));
    InMux I__9420 (
            .O(N__41565),
            .I(N__41192));
    InMux I__9419 (
            .O(N__41562),
            .I(N__41192));
    InMux I__9418 (
            .O(N__41561),
            .I(N__41192));
    InMux I__9417 (
            .O(N__41560),
            .I(N__41187));
    InMux I__9416 (
            .O(N__41559),
            .I(N__41187));
    Span4Mux_v I__9415 (
            .O(N__41552),
            .I(N__41184));
    Span4Mux_h I__9414 (
            .O(N__41549),
            .I(N__41177));
    LocalMux I__9413 (
            .O(N__41540),
            .I(N__41177));
    LocalMux I__9412 (
            .O(N__41531),
            .I(N__41177));
    Span4Mux_v I__9411 (
            .O(N__41524),
            .I(N__41174));
    Span4Mux_v I__9410 (
            .O(N__41519),
            .I(N__41169));
    Span4Mux_v I__9409 (
            .O(N__41512),
            .I(N__41169));
    LocalMux I__9408 (
            .O(N__41509),
            .I(N__41164));
    LocalMux I__9407 (
            .O(N__41502),
            .I(N__41164));
    InMux I__9406 (
            .O(N__41499),
            .I(N__41157));
    InMux I__9405 (
            .O(N__41496),
            .I(N__41157));
    InMux I__9404 (
            .O(N__41493),
            .I(N__41157));
    InMux I__9403 (
            .O(N__41490),
            .I(N__41146));
    InMux I__9402 (
            .O(N__41487),
            .I(N__41146));
    InMux I__9401 (
            .O(N__41484),
            .I(N__41146));
    InMux I__9400 (
            .O(N__41483),
            .I(N__41146));
    InMux I__9399 (
            .O(N__41480),
            .I(N__41146));
    InMux I__9398 (
            .O(N__41479),
            .I(N__41137));
    InMux I__9397 (
            .O(N__41478),
            .I(N__41137));
    InMux I__9396 (
            .O(N__41477),
            .I(N__41137));
    InMux I__9395 (
            .O(N__41476),
            .I(N__41137));
    InMux I__9394 (
            .O(N__41475),
            .I(N__41128));
    InMux I__9393 (
            .O(N__41474),
            .I(N__41128));
    InMux I__9392 (
            .O(N__41473),
            .I(N__41128));
    InMux I__9391 (
            .O(N__41472),
            .I(N__41128));
    Span4Mux_h I__9390 (
            .O(N__41467),
            .I(N__41123));
    Span4Mux_v I__9389 (
            .O(N__41462),
            .I(N__41123));
    Span4Mux_v I__9388 (
            .O(N__41457),
            .I(N__41116));
    Span4Mux_h I__9387 (
            .O(N__41454),
            .I(N__41116));
    LocalMux I__9386 (
            .O(N__41445),
            .I(N__41116));
    LocalMux I__9385 (
            .O(N__41436),
            .I(N__41103));
    Span4Mux_v I__9384 (
            .O(N__41421),
            .I(N__41103));
    LocalMux I__9383 (
            .O(N__41414),
            .I(N__41103));
    LocalMux I__9382 (
            .O(N__41407),
            .I(N__41103));
    LocalMux I__9381 (
            .O(N__41400),
            .I(N__41103));
    LocalMux I__9380 (
            .O(N__41393),
            .I(N__41103));
    Span4Mux_v I__9379 (
            .O(N__41390),
            .I(N__41094));
    Span4Mux_h I__9378 (
            .O(N__41387),
            .I(N__41094));
    Span4Mux_v I__9377 (
            .O(N__41372),
            .I(N__41094));
    LocalMux I__9376 (
            .O(N__41367),
            .I(N__41094));
    Span4Mux_v I__9375 (
            .O(N__41360),
            .I(N__41083));
    LocalMux I__9374 (
            .O(N__41353),
            .I(N__41083));
    LocalMux I__9373 (
            .O(N__41342),
            .I(N__41083));
    LocalMux I__9372 (
            .O(N__41333),
            .I(N__41083));
    LocalMux I__9371 (
            .O(N__41324),
            .I(N__41083));
    InMux I__9370 (
            .O(N__41323),
            .I(N__41078));
    InMux I__9369 (
            .O(N__41322),
            .I(N__41078));
    InMux I__9368 (
            .O(N__41321),
            .I(N__41069));
    InMux I__9367 (
            .O(N__41318),
            .I(N__41069));
    InMux I__9366 (
            .O(N__41317),
            .I(N__41069));
    InMux I__9365 (
            .O(N__41316),
            .I(N__41069));
    InMux I__9364 (
            .O(N__41315),
            .I(N__41064));
    InMux I__9363 (
            .O(N__41314),
            .I(N__41064));
    InMux I__9362 (
            .O(N__41311),
            .I(N__41055));
    InMux I__9361 (
            .O(N__41310),
            .I(N__41055));
    InMux I__9360 (
            .O(N__41309),
            .I(N__41055));
    InMux I__9359 (
            .O(N__41308),
            .I(N__41055));
    Sp12to4 I__9358 (
            .O(N__41305),
            .I(N__41042));
    LocalMux I__9357 (
            .O(N__41298),
            .I(N__41042));
    LocalMux I__9356 (
            .O(N__41291),
            .I(N__41042));
    Span12Mux_h I__9355 (
            .O(N__41288),
            .I(N__41042));
    LocalMux I__9354 (
            .O(N__41285),
            .I(N__41042));
    LocalMux I__9353 (
            .O(N__41278),
            .I(N__41042));
    LocalMux I__9352 (
            .O(N__41271),
            .I(N__41037));
    LocalMux I__9351 (
            .O(N__41264),
            .I(N__41037));
    LocalMux I__9350 (
            .O(N__41259),
            .I(N__41014));
    LocalMux I__9349 (
            .O(N__41252),
            .I(N__41014));
    LocalMux I__9348 (
            .O(N__41241),
            .I(N__41014));
    LocalMux I__9347 (
            .O(N__41232),
            .I(N__41014));
    LocalMux I__9346 (
            .O(N__41227),
            .I(N__41014));
    LocalMux I__9345 (
            .O(N__41224),
            .I(N__41014));
    Sp12to4 I__9344 (
            .O(N__41219),
            .I(N__41014));
    LocalMux I__9343 (
            .O(N__41210),
            .I(N__41014));
    LocalMux I__9342 (
            .O(N__41201),
            .I(N__41014));
    LocalMux I__9341 (
            .O(N__41192),
            .I(N__41014));
    LocalMux I__9340 (
            .O(N__41187),
            .I(N__41014));
    Span4Mux_h I__9339 (
            .O(N__41184),
            .I(N__41009));
    Span4Mux_v I__9338 (
            .O(N__41177),
            .I(N__41009));
    Span4Mux_h I__9337 (
            .O(N__41174),
            .I(N__40994));
    Span4Mux_h I__9336 (
            .O(N__41169),
            .I(N__40994));
    Span4Mux_v I__9335 (
            .O(N__41164),
            .I(N__40994));
    LocalMux I__9334 (
            .O(N__41157),
            .I(N__40994));
    LocalMux I__9333 (
            .O(N__41146),
            .I(N__40994));
    LocalMux I__9332 (
            .O(N__41137),
            .I(N__40994));
    LocalMux I__9331 (
            .O(N__41128),
            .I(N__40994));
    Span4Mux_h I__9330 (
            .O(N__41123),
            .I(N__40987));
    Span4Mux_v I__9329 (
            .O(N__41116),
            .I(N__40987));
    Span4Mux_v I__9328 (
            .O(N__41103),
            .I(N__40987));
    Span4Mux_v I__9327 (
            .O(N__41094),
            .I(N__40974));
    Span4Mux_v I__9326 (
            .O(N__41083),
            .I(N__40974));
    LocalMux I__9325 (
            .O(N__41078),
            .I(N__40974));
    LocalMux I__9324 (
            .O(N__41069),
            .I(N__40974));
    LocalMux I__9323 (
            .O(N__41064),
            .I(N__40974));
    LocalMux I__9322 (
            .O(N__41055),
            .I(N__40974));
    Span12Mux_v I__9321 (
            .O(N__41042),
            .I(N__40971));
    Span12Mux_s10_h I__9320 (
            .O(N__41037),
            .I(N__40966));
    Span12Mux_s9_v I__9319 (
            .O(N__41014),
            .I(N__40966));
    Span4Mux_v I__9318 (
            .O(N__41009),
            .I(N__40961));
    Span4Mux_v I__9317 (
            .O(N__40994),
            .I(N__40961));
    Span4Mux_v I__9316 (
            .O(N__40987),
            .I(N__40956));
    Span4Mux_v I__9315 (
            .O(N__40974),
            .I(N__40956));
    Odrv12 I__9314 (
            .O(N__40971),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__9313 (
            .O(N__40966),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__9312 (
            .O(N__40961),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__9311 (
            .O(N__40956),
            .I(CONSTANT_ONE_NET));
    InMux I__9310 (
            .O(N__40947),
            .I(N__40943));
    InMux I__9309 (
            .O(N__40946),
            .I(N__40940));
    LocalMux I__9308 (
            .O(N__40943),
            .I(N__40937));
    LocalMux I__9307 (
            .O(N__40940),
            .I(N__40934));
    Odrv4 I__9306 (
            .O(N__40937),
            .I(\nx.n2489 ));
    Odrv4 I__9305 (
            .O(N__40934),
            .I(\nx.n2489 ));
    CascadeMux I__9304 (
            .O(N__40929),
            .I(N__40923));
    InMux I__9303 (
            .O(N__40928),
            .I(N__40918));
    CascadeMux I__9302 (
            .O(N__40927),
            .I(N__40915));
    InMux I__9301 (
            .O(N__40926),
            .I(N__40911));
    InMux I__9300 (
            .O(N__40923),
            .I(N__40908));
    CascadeMux I__9299 (
            .O(N__40922),
            .I(N__40904));
    CascadeMux I__9298 (
            .O(N__40921),
            .I(N__40895));
    LocalMux I__9297 (
            .O(N__40918),
            .I(N__40891));
    InMux I__9296 (
            .O(N__40915),
            .I(N__40886));
    InMux I__9295 (
            .O(N__40914),
            .I(N__40886));
    LocalMux I__9294 (
            .O(N__40911),
            .I(N__40881));
    LocalMux I__9293 (
            .O(N__40908),
            .I(N__40881));
    InMux I__9292 (
            .O(N__40907),
            .I(N__40874));
    InMux I__9291 (
            .O(N__40904),
            .I(N__40874));
    InMux I__9290 (
            .O(N__40903),
            .I(N__40874));
    InMux I__9289 (
            .O(N__40902),
            .I(N__40871));
    InMux I__9288 (
            .O(N__40901),
            .I(N__40868));
    CascadeMux I__9287 (
            .O(N__40900),
            .I(N__40865));
    InMux I__9286 (
            .O(N__40899),
            .I(N__40856));
    InMux I__9285 (
            .O(N__40898),
            .I(N__40849));
    InMux I__9284 (
            .O(N__40895),
            .I(N__40849));
    InMux I__9283 (
            .O(N__40894),
            .I(N__40849));
    Span4Mux_v I__9282 (
            .O(N__40891),
            .I(N__40840));
    LocalMux I__9281 (
            .O(N__40886),
            .I(N__40840));
    Span4Mux_v I__9280 (
            .O(N__40881),
            .I(N__40840));
    LocalMux I__9279 (
            .O(N__40874),
            .I(N__40840));
    LocalMux I__9278 (
            .O(N__40871),
            .I(N__40835));
    LocalMux I__9277 (
            .O(N__40868),
            .I(N__40835));
    InMux I__9276 (
            .O(N__40865),
            .I(N__40828));
    InMux I__9275 (
            .O(N__40864),
            .I(N__40828));
    InMux I__9274 (
            .O(N__40863),
            .I(N__40828));
    InMux I__9273 (
            .O(N__40862),
            .I(N__40819));
    InMux I__9272 (
            .O(N__40861),
            .I(N__40819));
    InMux I__9271 (
            .O(N__40860),
            .I(N__40819));
    InMux I__9270 (
            .O(N__40859),
            .I(N__40819));
    LocalMux I__9269 (
            .O(N__40856),
            .I(\nx.n2522 ));
    LocalMux I__9268 (
            .O(N__40849),
            .I(\nx.n2522 ));
    Odrv4 I__9267 (
            .O(N__40840),
            .I(\nx.n2522 ));
    Odrv4 I__9266 (
            .O(N__40835),
            .I(\nx.n2522 ));
    LocalMux I__9265 (
            .O(N__40828),
            .I(\nx.n2522 ));
    LocalMux I__9264 (
            .O(N__40819),
            .I(\nx.n2522 ));
    InMux I__9263 (
            .O(N__40806),
            .I(\nx.n10958 ));
    CascadeMux I__9262 (
            .O(N__40803),
            .I(N__40799));
    InMux I__9261 (
            .O(N__40802),
            .I(N__40796));
    InMux I__9260 (
            .O(N__40799),
            .I(N__40793));
    LocalMux I__9259 (
            .O(N__40796),
            .I(N__40790));
    LocalMux I__9258 (
            .O(N__40793),
            .I(N__40787));
    Span4Mux_v I__9257 (
            .O(N__40790),
            .I(N__40784));
    Odrv4 I__9256 (
            .O(N__40787),
            .I(\nx.n2588 ));
    Odrv4 I__9255 (
            .O(N__40784),
            .I(\nx.n2588 ));
    IoInMux I__9254 (
            .O(N__40779),
            .I(N__40776));
    LocalMux I__9253 (
            .O(N__40776),
            .I(N__40773));
    Span12Mux_s11_h I__9252 (
            .O(N__40773),
            .I(N__40770));
    Span12Mux_v I__9251 (
            .O(N__40770),
            .I(N__40766));
    InMux I__9250 (
            .O(N__40769),
            .I(N__40763));
    Odrv12 I__9249 (
            .O(N__40766),
            .I(pin_oe_12));
    LocalMux I__9248 (
            .O(N__40763),
            .I(pin_oe_12));
    InMux I__9247 (
            .O(N__40758),
            .I(N__40755));
    LocalMux I__9246 (
            .O(N__40755),
            .I(n45));
    InMux I__9245 (
            .O(N__40752),
            .I(bfn_17_15_0_));
    InMux I__9244 (
            .O(N__40749),
            .I(n10700));
    InMux I__9243 (
            .O(N__40746),
            .I(n10701));
    InMux I__9242 (
            .O(N__40743),
            .I(n10702));
    CascadeMux I__9241 (
            .O(N__40740),
            .I(N__40737));
    InMux I__9240 (
            .O(N__40737),
            .I(N__40733));
    InMux I__9239 (
            .O(N__40736),
            .I(N__40730));
    LocalMux I__9238 (
            .O(N__40733),
            .I(N__40726));
    LocalMux I__9237 (
            .O(N__40730),
            .I(N__40723));
    InMux I__9236 (
            .O(N__40729),
            .I(N__40720));
    Span4Mux_h I__9235 (
            .O(N__40726),
            .I(N__40717));
    Span4Mux_h I__9234 (
            .O(N__40723),
            .I(N__40714));
    LocalMux I__9233 (
            .O(N__40720),
            .I(\nx.n2498 ));
    Odrv4 I__9232 (
            .O(N__40717),
            .I(\nx.n2498 ));
    Odrv4 I__9231 (
            .O(N__40714),
            .I(\nx.n2498 ));
    InMux I__9230 (
            .O(N__40707),
            .I(N__40704));
    LocalMux I__9229 (
            .O(N__40704),
            .I(N__40701));
    Span4Mux_v I__9228 (
            .O(N__40701),
            .I(N__40698));
    Odrv4 I__9227 (
            .O(N__40698),
            .I(\nx.n2565 ));
    InMux I__9226 (
            .O(N__40695),
            .I(\nx.n10949 ));
    InMux I__9225 (
            .O(N__40692),
            .I(N__40687));
    InMux I__9224 (
            .O(N__40691),
            .I(N__40684));
    InMux I__9223 (
            .O(N__40690),
            .I(N__40681));
    LocalMux I__9222 (
            .O(N__40687),
            .I(\nx.n2497 ));
    LocalMux I__9221 (
            .O(N__40684),
            .I(\nx.n2497 ));
    LocalMux I__9220 (
            .O(N__40681),
            .I(\nx.n2497 ));
    CascadeMux I__9219 (
            .O(N__40674),
            .I(N__40671));
    InMux I__9218 (
            .O(N__40671),
            .I(N__40668));
    LocalMux I__9217 (
            .O(N__40668),
            .I(N__40665));
    Odrv4 I__9216 (
            .O(N__40665),
            .I(\nx.n2564 ));
    InMux I__9215 (
            .O(N__40662),
            .I(\nx.n10950 ));
    InMux I__9214 (
            .O(N__40659),
            .I(N__40655));
    InMux I__9213 (
            .O(N__40658),
            .I(N__40652));
    LocalMux I__9212 (
            .O(N__40655),
            .I(\nx.n2496 ));
    LocalMux I__9211 (
            .O(N__40652),
            .I(\nx.n2496 ));
    InMux I__9210 (
            .O(N__40647),
            .I(N__40644));
    LocalMux I__9209 (
            .O(N__40644),
            .I(\nx.n2563 ));
    InMux I__9208 (
            .O(N__40641),
            .I(\nx.n10951 ));
    CascadeMux I__9207 (
            .O(N__40638),
            .I(N__40634));
    InMux I__9206 (
            .O(N__40637),
            .I(N__40631));
    InMux I__9205 (
            .O(N__40634),
            .I(N__40628));
    LocalMux I__9204 (
            .O(N__40631),
            .I(\nx.n2495 ));
    LocalMux I__9203 (
            .O(N__40628),
            .I(\nx.n2495 ));
    CascadeMux I__9202 (
            .O(N__40623),
            .I(N__40620));
    InMux I__9201 (
            .O(N__40620),
            .I(N__40617));
    LocalMux I__9200 (
            .O(N__40617),
            .I(N__40614));
    Odrv4 I__9199 (
            .O(N__40614),
            .I(\nx.n2562 ));
    InMux I__9198 (
            .O(N__40611),
            .I(\nx.n10952 ));
    CascadeMux I__9197 (
            .O(N__40608),
            .I(N__40605));
    InMux I__9196 (
            .O(N__40605),
            .I(N__40601));
    InMux I__9195 (
            .O(N__40604),
            .I(N__40597));
    LocalMux I__9194 (
            .O(N__40601),
            .I(N__40594));
    InMux I__9193 (
            .O(N__40600),
            .I(N__40591));
    LocalMux I__9192 (
            .O(N__40597),
            .I(\nx.n2494 ));
    Odrv4 I__9191 (
            .O(N__40594),
            .I(\nx.n2494 ));
    LocalMux I__9190 (
            .O(N__40591),
            .I(\nx.n2494 ));
    CascadeMux I__9189 (
            .O(N__40584),
            .I(N__40581));
    InMux I__9188 (
            .O(N__40581),
            .I(N__40578));
    LocalMux I__9187 (
            .O(N__40578),
            .I(N__40575));
    Odrv4 I__9186 (
            .O(N__40575),
            .I(\nx.n2561 ));
    InMux I__9185 (
            .O(N__40572),
            .I(bfn_16_26_0_));
    CascadeMux I__9184 (
            .O(N__40569),
            .I(N__40566));
    InMux I__9183 (
            .O(N__40566),
            .I(N__40562));
    CascadeMux I__9182 (
            .O(N__40565),
            .I(N__40559));
    LocalMux I__9181 (
            .O(N__40562),
            .I(N__40555));
    InMux I__9180 (
            .O(N__40559),
            .I(N__40552));
    InMux I__9179 (
            .O(N__40558),
            .I(N__40549));
    Odrv4 I__9178 (
            .O(N__40555),
            .I(\nx.n2493 ));
    LocalMux I__9177 (
            .O(N__40552),
            .I(\nx.n2493 ));
    LocalMux I__9176 (
            .O(N__40549),
            .I(\nx.n2493 ));
    InMux I__9175 (
            .O(N__40542),
            .I(N__40539));
    LocalMux I__9174 (
            .O(N__40539),
            .I(N__40536));
    Span4Mux_h I__9173 (
            .O(N__40536),
            .I(N__40533));
    Odrv4 I__9172 (
            .O(N__40533),
            .I(\nx.n2560 ));
    InMux I__9171 (
            .O(N__40530),
            .I(\nx.n10954 ));
    InMux I__9170 (
            .O(N__40527),
            .I(N__40524));
    LocalMux I__9169 (
            .O(N__40524),
            .I(N__40520));
    CascadeMux I__9168 (
            .O(N__40523),
            .I(N__40517));
    Span4Mux_v I__9167 (
            .O(N__40520),
            .I(N__40513));
    InMux I__9166 (
            .O(N__40517),
            .I(N__40510));
    InMux I__9165 (
            .O(N__40516),
            .I(N__40507));
    Odrv4 I__9164 (
            .O(N__40513),
            .I(\nx.n2492 ));
    LocalMux I__9163 (
            .O(N__40510),
            .I(\nx.n2492 ));
    LocalMux I__9162 (
            .O(N__40507),
            .I(\nx.n2492 ));
    CascadeMux I__9161 (
            .O(N__40500),
            .I(N__40497));
    InMux I__9160 (
            .O(N__40497),
            .I(N__40494));
    LocalMux I__9159 (
            .O(N__40494),
            .I(N__40491));
    Span4Mux_v I__9158 (
            .O(N__40491),
            .I(N__40488));
    Odrv4 I__9157 (
            .O(N__40488),
            .I(\nx.n2559 ));
    InMux I__9156 (
            .O(N__40485),
            .I(\nx.n10955 ));
    CascadeMux I__9155 (
            .O(N__40482),
            .I(N__40479));
    InMux I__9154 (
            .O(N__40479),
            .I(N__40476));
    LocalMux I__9153 (
            .O(N__40476),
            .I(N__40471));
    InMux I__9152 (
            .O(N__40475),
            .I(N__40466));
    InMux I__9151 (
            .O(N__40474),
            .I(N__40466));
    Span4Mux_h I__9150 (
            .O(N__40471),
            .I(N__40463));
    LocalMux I__9149 (
            .O(N__40466),
            .I(\nx.n2506 ));
    Odrv4 I__9148 (
            .O(N__40463),
            .I(\nx.n2506 ));
    InMux I__9147 (
            .O(N__40458),
            .I(N__40455));
    LocalMux I__9146 (
            .O(N__40455),
            .I(N__40452));
    Odrv4 I__9145 (
            .O(N__40452),
            .I(\nx.n2573 ));
    InMux I__9144 (
            .O(N__40449),
            .I(\nx.n10941 ));
    CascadeMux I__9143 (
            .O(N__40446),
            .I(N__40442));
    CascadeMux I__9142 (
            .O(N__40445),
            .I(N__40439));
    InMux I__9141 (
            .O(N__40442),
            .I(N__40436));
    InMux I__9140 (
            .O(N__40439),
            .I(N__40433));
    LocalMux I__9139 (
            .O(N__40436),
            .I(\nx.n2505 ));
    LocalMux I__9138 (
            .O(N__40433),
            .I(\nx.n2505 ));
    InMux I__9137 (
            .O(N__40428),
            .I(N__40425));
    LocalMux I__9136 (
            .O(N__40425),
            .I(\nx.n2572 ));
    InMux I__9135 (
            .O(N__40422),
            .I(\nx.n10942 ));
    CascadeMux I__9134 (
            .O(N__40419),
            .I(N__40416));
    InMux I__9133 (
            .O(N__40416),
            .I(N__40412));
    CascadeMux I__9132 (
            .O(N__40415),
            .I(N__40409));
    LocalMux I__9131 (
            .O(N__40412),
            .I(N__40405));
    InMux I__9130 (
            .O(N__40409),
            .I(N__40402));
    InMux I__9129 (
            .O(N__40408),
            .I(N__40399));
    Span4Mux_h I__9128 (
            .O(N__40405),
            .I(N__40396));
    LocalMux I__9127 (
            .O(N__40402),
            .I(\nx.n2504 ));
    LocalMux I__9126 (
            .O(N__40399),
            .I(\nx.n2504 ));
    Odrv4 I__9125 (
            .O(N__40396),
            .I(\nx.n2504 ));
    InMux I__9124 (
            .O(N__40389),
            .I(N__40386));
    LocalMux I__9123 (
            .O(N__40386),
            .I(N__40383));
    Span4Mux_h I__9122 (
            .O(N__40383),
            .I(N__40380));
    Odrv4 I__9121 (
            .O(N__40380),
            .I(\nx.n2571 ));
    InMux I__9120 (
            .O(N__40377),
            .I(\nx.n10943 ));
    InMux I__9119 (
            .O(N__40374),
            .I(N__40369));
    InMux I__9118 (
            .O(N__40373),
            .I(N__40366));
    InMux I__9117 (
            .O(N__40372),
            .I(N__40363));
    LocalMux I__9116 (
            .O(N__40369),
            .I(N__40360));
    LocalMux I__9115 (
            .O(N__40366),
            .I(N__40357));
    LocalMux I__9114 (
            .O(N__40363),
            .I(N__40354));
    Odrv4 I__9113 (
            .O(N__40360),
            .I(\nx.n2503 ));
    Odrv4 I__9112 (
            .O(N__40357),
            .I(\nx.n2503 ));
    Odrv4 I__9111 (
            .O(N__40354),
            .I(\nx.n2503 ));
    CascadeMux I__9110 (
            .O(N__40347),
            .I(N__40344));
    InMux I__9109 (
            .O(N__40344),
            .I(N__40341));
    LocalMux I__9108 (
            .O(N__40341),
            .I(N__40338));
    Span4Mux_h I__9107 (
            .O(N__40338),
            .I(N__40335));
    Odrv4 I__9106 (
            .O(N__40335),
            .I(\nx.n2570 ));
    InMux I__9105 (
            .O(N__40332),
            .I(\nx.n10944 ));
    CascadeMux I__9104 (
            .O(N__40329),
            .I(N__40326));
    InMux I__9103 (
            .O(N__40326),
            .I(N__40323));
    LocalMux I__9102 (
            .O(N__40323),
            .I(N__40318));
    InMux I__9101 (
            .O(N__40322),
            .I(N__40315));
    InMux I__9100 (
            .O(N__40321),
            .I(N__40312));
    Span4Mux_h I__9099 (
            .O(N__40318),
            .I(N__40309));
    LocalMux I__9098 (
            .O(N__40315),
            .I(\nx.n2502 ));
    LocalMux I__9097 (
            .O(N__40312),
            .I(\nx.n2502 ));
    Odrv4 I__9096 (
            .O(N__40309),
            .I(\nx.n2502 ));
    InMux I__9095 (
            .O(N__40302),
            .I(N__40299));
    LocalMux I__9094 (
            .O(N__40299),
            .I(N__40296));
    Span4Mux_h I__9093 (
            .O(N__40296),
            .I(N__40293));
    Odrv4 I__9092 (
            .O(N__40293),
            .I(\nx.n2569 ));
    InMux I__9091 (
            .O(N__40290),
            .I(bfn_16_25_0_));
    CascadeMux I__9090 (
            .O(N__40287),
            .I(N__40284));
    InMux I__9089 (
            .O(N__40284),
            .I(N__40280));
    CascadeMux I__9088 (
            .O(N__40283),
            .I(N__40277));
    LocalMux I__9087 (
            .O(N__40280),
            .I(N__40274));
    InMux I__9086 (
            .O(N__40277),
            .I(N__40271));
    Span4Mux_h I__9085 (
            .O(N__40274),
            .I(N__40268));
    LocalMux I__9084 (
            .O(N__40271),
            .I(\nx.n2501 ));
    Odrv4 I__9083 (
            .O(N__40268),
            .I(\nx.n2501 ));
    InMux I__9082 (
            .O(N__40263),
            .I(N__40260));
    LocalMux I__9081 (
            .O(N__40260),
            .I(N__40257));
    Span4Mux_h I__9080 (
            .O(N__40257),
            .I(N__40254));
    Odrv4 I__9079 (
            .O(N__40254),
            .I(\nx.n2568 ));
    InMux I__9078 (
            .O(N__40251),
            .I(\nx.n10946 ));
    CascadeMux I__9077 (
            .O(N__40248),
            .I(N__40245));
    InMux I__9076 (
            .O(N__40245),
            .I(N__40242));
    LocalMux I__9075 (
            .O(N__40242),
            .I(N__40238));
    InMux I__9074 (
            .O(N__40241),
            .I(N__40234));
    Span4Mux_h I__9073 (
            .O(N__40238),
            .I(N__40231));
    InMux I__9072 (
            .O(N__40237),
            .I(N__40228));
    LocalMux I__9071 (
            .O(N__40234),
            .I(\nx.n2500 ));
    Odrv4 I__9070 (
            .O(N__40231),
            .I(\nx.n2500 ));
    LocalMux I__9069 (
            .O(N__40228),
            .I(\nx.n2500 ));
    CascadeMux I__9068 (
            .O(N__40221),
            .I(N__40218));
    InMux I__9067 (
            .O(N__40218),
            .I(N__40215));
    LocalMux I__9066 (
            .O(N__40215),
            .I(N__40212));
    Span4Mux_v I__9065 (
            .O(N__40212),
            .I(N__40209));
    Odrv4 I__9064 (
            .O(N__40209),
            .I(\nx.n2567 ));
    InMux I__9063 (
            .O(N__40206),
            .I(\nx.n10947 ));
    CascadeMux I__9062 (
            .O(N__40203),
            .I(N__40198));
    CascadeMux I__9061 (
            .O(N__40202),
            .I(N__40195));
    InMux I__9060 (
            .O(N__40201),
            .I(N__40192));
    InMux I__9059 (
            .O(N__40198),
            .I(N__40189));
    InMux I__9058 (
            .O(N__40195),
            .I(N__40186));
    LocalMux I__9057 (
            .O(N__40192),
            .I(N__40181));
    LocalMux I__9056 (
            .O(N__40189),
            .I(N__40181));
    LocalMux I__9055 (
            .O(N__40186),
            .I(\nx.n2499 ));
    Odrv4 I__9054 (
            .O(N__40181),
            .I(\nx.n2499 ));
    InMux I__9053 (
            .O(N__40176),
            .I(N__40173));
    LocalMux I__9052 (
            .O(N__40173),
            .I(N__40170));
    Odrv4 I__9051 (
            .O(N__40170),
            .I(\nx.n2566 ));
    InMux I__9050 (
            .O(N__40167),
            .I(\nx.n10948 ));
    CascadeMux I__9049 (
            .O(N__40164),
            .I(N__40160));
    CascadeMux I__9048 (
            .O(N__40163),
            .I(N__40156));
    InMux I__9047 (
            .O(N__40160),
            .I(N__40153));
    InMux I__9046 (
            .O(N__40159),
            .I(N__40148));
    InMux I__9045 (
            .O(N__40156),
            .I(N__40148));
    LocalMux I__9044 (
            .O(N__40153),
            .I(N__40145));
    LocalMux I__9043 (
            .O(N__40148),
            .I(N__40142));
    Span4Mux_h I__9042 (
            .O(N__40145),
            .I(N__40137));
    Span4Mux_h I__9041 (
            .O(N__40142),
            .I(N__40137));
    Odrv4 I__9040 (
            .O(N__40137),
            .I(\nx.n2590 ));
    CascadeMux I__9039 (
            .O(N__40134),
            .I(N__40131));
    InMux I__9038 (
            .O(N__40131),
            .I(N__40128));
    LocalMux I__9037 (
            .O(N__40128),
            .I(N__40125));
    Odrv12 I__9036 (
            .O(N__40125),
            .I(\nx.n2657 ));
    InMux I__9035 (
            .O(N__40122),
            .I(\nx.n10978 ));
    InMux I__9034 (
            .O(N__40119),
            .I(N__40116));
    LocalMux I__9033 (
            .O(N__40116),
            .I(N__40113));
    Odrv12 I__9032 (
            .O(N__40113),
            .I(\nx.n2656 ));
    InMux I__9031 (
            .O(N__40110),
            .I(\nx.n10979 ));
    CascadeMux I__9030 (
            .O(N__40107),
            .I(N__40102));
    InMux I__9029 (
            .O(N__40106),
            .I(N__40088));
    InMux I__9028 (
            .O(N__40105),
            .I(N__40085));
    InMux I__9027 (
            .O(N__40102),
            .I(N__40080));
    InMux I__9026 (
            .O(N__40101),
            .I(N__40080));
    InMux I__9025 (
            .O(N__40100),
            .I(N__40065));
    InMux I__9024 (
            .O(N__40099),
            .I(N__40065));
    InMux I__9023 (
            .O(N__40098),
            .I(N__40065));
    InMux I__9022 (
            .O(N__40097),
            .I(N__40065));
    InMux I__9021 (
            .O(N__40096),
            .I(N__40065));
    InMux I__9020 (
            .O(N__40095),
            .I(N__40062));
    CascadeMux I__9019 (
            .O(N__40094),
            .I(N__40059));
    CascadeMux I__9018 (
            .O(N__40093),
            .I(N__40055));
    CascadeMux I__9017 (
            .O(N__40092),
            .I(N__40052));
    CascadeMux I__9016 (
            .O(N__40091),
            .I(N__40048));
    LocalMux I__9015 (
            .O(N__40088),
            .I(N__40039));
    LocalMux I__9014 (
            .O(N__40085),
            .I(N__40039));
    LocalMux I__9013 (
            .O(N__40080),
            .I(N__40039));
    InMux I__9012 (
            .O(N__40079),
            .I(N__40034));
    InMux I__9011 (
            .O(N__40078),
            .I(N__40034));
    InMux I__9010 (
            .O(N__40077),
            .I(N__40031));
    InMux I__9009 (
            .O(N__40076),
            .I(N__40028));
    LocalMux I__9008 (
            .O(N__40065),
            .I(N__40023));
    LocalMux I__9007 (
            .O(N__40062),
            .I(N__40023));
    InMux I__9006 (
            .O(N__40059),
            .I(N__40012));
    InMux I__9005 (
            .O(N__40058),
            .I(N__40012));
    InMux I__9004 (
            .O(N__40055),
            .I(N__40012));
    InMux I__9003 (
            .O(N__40052),
            .I(N__40012));
    InMux I__9002 (
            .O(N__40051),
            .I(N__40012));
    InMux I__9001 (
            .O(N__40048),
            .I(N__40005));
    InMux I__9000 (
            .O(N__40047),
            .I(N__40005));
    InMux I__8999 (
            .O(N__40046),
            .I(N__40005));
    Span4Mux_h I__8998 (
            .O(N__40039),
            .I(N__40002));
    LocalMux I__8997 (
            .O(N__40034),
            .I(\nx.n2621 ));
    LocalMux I__8996 (
            .O(N__40031),
            .I(\nx.n2621 ));
    LocalMux I__8995 (
            .O(N__40028),
            .I(\nx.n2621 ));
    Odrv12 I__8994 (
            .O(N__40023),
            .I(\nx.n2621 ));
    LocalMux I__8993 (
            .O(N__40012),
            .I(\nx.n2621 ));
    LocalMux I__8992 (
            .O(N__40005),
            .I(\nx.n2621 ));
    Odrv4 I__8991 (
            .O(N__40002),
            .I(\nx.n2621 ));
    InMux I__8990 (
            .O(N__39987),
            .I(\nx.n10980 ));
    CascadeMux I__8989 (
            .O(N__39984),
            .I(N__39980));
    InMux I__8988 (
            .O(N__39983),
            .I(N__39977));
    InMux I__8987 (
            .O(N__39980),
            .I(N__39974));
    LocalMux I__8986 (
            .O(N__39977),
            .I(N__39971));
    LocalMux I__8985 (
            .O(N__39974),
            .I(N__39968));
    Span4Mux_h I__8984 (
            .O(N__39971),
            .I(N__39965));
    Span4Mux_h I__8983 (
            .O(N__39968),
            .I(N__39962));
    Span4Mux_h I__8982 (
            .O(N__39965),
            .I(N__39959));
    Span4Mux_h I__8981 (
            .O(N__39962),
            .I(N__39956));
    Odrv4 I__8980 (
            .O(N__39959),
            .I(\nx.n2687 ));
    Odrv4 I__8979 (
            .O(N__39956),
            .I(\nx.n2687 ));
    InMux I__8978 (
            .O(N__39951),
            .I(N__39944));
    InMux I__8977 (
            .O(N__39950),
            .I(N__39944));
    CascadeMux I__8976 (
            .O(N__39949),
            .I(N__39941));
    LocalMux I__8975 (
            .O(N__39944),
            .I(N__39938));
    InMux I__8974 (
            .O(N__39941),
            .I(N__39935));
    Span4Mux_h I__8973 (
            .O(N__39938),
            .I(N__39932));
    LocalMux I__8972 (
            .O(N__39935),
            .I(\nx.n2589 ));
    Odrv4 I__8971 (
            .O(N__39932),
            .I(\nx.n2589 ));
    InMux I__8970 (
            .O(N__39927),
            .I(N__39924));
    LocalMux I__8969 (
            .O(N__39924),
            .I(N__39918));
    InMux I__8968 (
            .O(N__39923),
            .I(N__39915));
    InMux I__8967 (
            .O(N__39922),
            .I(N__39912));
    InMux I__8966 (
            .O(N__39921),
            .I(N__39909));
    Span4Mux_h I__8965 (
            .O(N__39918),
            .I(N__39906));
    LocalMux I__8964 (
            .O(N__39915),
            .I(N__39903));
    LocalMux I__8963 (
            .O(N__39912),
            .I(N__39900));
    LocalMux I__8962 (
            .O(N__39909),
            .I(N__39896));
    Span4Mux_h I__8961 (
            .O(N__39906),
            .I(N__39893));
    Span4Mux_v I__8960 (
            .O(N__39903),
            .I(N__39890));
    Span4Mux_h I__8959 (
            .O(N__39900),
            .I(N__39887));
    InMux I__8958 (
            .O(N__39899),
            .I(N__39884));
    Sp12to4 I__8957 (
            .O(N__39896),
            .I(N__39881));
    Span4Mux_h I__8956 (
            .O(N__39893),
            .I(N__39878));
    Span4Mux_h I__8955 (
            .O(N__39890),
            .I(N__39873));
    Span4Mux_h I__8954 (
            .O(N__39887),
            .I(N__39873));
    LocalMux I__8953 (
            .O(N__39884),
            .I(\nx.bit_ctr_10 ));
    Odrv12 I__8952 (
            .O(N__39881),
            .I(\nx.bit_ctr_10 ));
    Odrv4 I__8951 (
            .O(N__39878),
            .I(\nx.bit_ctr_10 ));
    Odrv4 I__8950 (
            .O(N__39873),
            .I(\nx.bit_ctr_10 ));
    InMux I__8949 (
            .O(N__39864),
            .I(N__39861));
    LocalMux I__8948 (
            .O(N__39861),
            .I(N__39858));
    Span4Mux_v I__8947 (
            .O(N__39858),
            .I(N__39855));
    Odrv4 I__8946 (
            .O(N__39855),
            .I(\nx.n2577 ));
    InMux I__8945 (
            .O(N__39852),
            .I(bfn_16_24_0_));
    CascadeMux I__8944 (
            .O(N__39849),
            .I(N__39845));
    InMux I__8943 (
            .O(N__39848),
            .I(N__39842));
    InMux I__8942 (
            .O(N__39845),
            .I(N__39839));
    LocalMux I__8941 (
            .O(N__39842),
            .I(N__39835));
    LocalMux I__8940 (
            .O(N__39839),
            .I(N__39832));
    InMux I__8939 (
            .O(N__39838),
            .I(N__39829));
    Span4Mux_v I__8938 (
            .O(N__39835),
            .I(N__39824));
    Span4Mux_v I__8937 (
            .O(N__39832),
            .I(N__39824));
    LocalMux I__8936 (
            .O(N__39829),
            .I(\nx.n2509 ));
    Odrv4 I__8935 (
            .O(N__39824),
            .I(\nx.n2509 ));
    InMux I__8934 (
            .O(N__39819),
            .I(N__39816));
    LocalMux I__8933 (
            .O(N__39816),
            .I(N__39813));
    Odrv4 I__8932 (
            .O(N__39813),
            .I(\nx.n2576 ));
    InMux I__8931 (
            .O(N__39810),
            .I(\nx.n10938 ));
    CascadeMux I__8930 (
            .O(N__39807),
            .I(N__39802));
    InMux I__8929 (
            .O(N__39806),
            .I(N__39797));
    InMux I__8928 (
            .O(N__39805),
            .I(N__39797));
    InMux I__8927 (
            .O(N__39802),
            .I(N__39794));
    LocalMux I__8926 (
            .O(N__39797),
            .I(\nx.n2508 ));
    LocalMux I__8925 (
            .O(N__39794),
            .I(\nx.n2508 ));
    CascadeMux I__8924 (
            .O(N__39789),
            .I(N__39786));
    InMux I__8923 (
            .O(N__39786),
            .I(N__39783));
    LocalMux I__8922 (
            .O(N__39783),
            .I(N__39780));
    Odrv4 I__8921 (
            .O(N__39780),
            .I(\nx.n2575 ));
    InMux I__8920 (
            .O(N__39777),
            .I(\nx.n10939 ));
    CascadeMux I__8919 (
            .O(N__39774),
            .I(N__39771));
    InMux I__8918 (
            .O(N__39771),
            .I(N__39767));
    InMux I__8917 (
            .O(N__39770),
            .I(N__39764));
    LocalMux I__8916 (
            .O(N__39767),
            .I(N__39761));
    LocalMux I__8915 (
            .O(N__39764),
            .I(N__39758));
    Span4Mux_h I__8914 (
            .O(N__39761),
            .I(N__39755));
    Span4Mux_v I__8913 (
            .O(N__39758),
            .I(N__39752));
    Odrv4 I__8912 (
            .O(N__39755),
            .I(\nx.n2507 ));
    Odrv4 I__8911 (
            .O(N__39752),
            .I(\nx.n2507 ));
    InMux I__8910 (
            .O(N__39747),
            .I(N__39744));
    LocalMux I__8909 (
            .O(N__39744),
            .I(N__39741));
    Odrv4 I__8908 (
            .O(N__39741),
            .I(\nx.n2574 ));
    InMux I__8907 (
            .O(N__39738),
            .I(\nx.n10940 ));
    CascadeMux I__8906 (
            .O(N__39735),
            .I(N__39732));
    InMux I__8905 (
            .O(N__39732),
            .I(N__39728));
    CascadeMux I__8904 (
            .O(N__39731),
            .I(N__39724));
    LocalMux I__8903 (
            .O(N__39728),
            .I(N__39721));
    InMux I__8902 (
            .O(N__39727),
            .I(N__39718));
    InMux I__8901 (
            .O(N__39724),
            .I(N__39715));
    Span4Mux_v I__8900 (
            .O(N__39721),
            .I(N__39710));
    LocalMux I__8899 (
            .O(N__39718),
            .I(N__39710));
    LocalMux I__8898 (
            .O(N__39715),
            .I(\nx.n2598 ));
    Odrv4 I__8897 (
            .O(N__39710),
            .I(\nx.n2598 ));
    InMux I__8896 (
            .O(N__39705),
            .I(N__39702));
    LocalMux I__8895 (
            .O(N__39702),
            .I(N__39699));
    Span4Mux_v I__8894 (
            .O(N__39699),
            .I(N__39696));
    Span4Mux_h I__8893 (
            .O(N__39696),
            .I(N__39693));
    Odrv4 I__8892 (
            .O(N__39693),
            .I(\nx.n2665 ));
    InMux I__8891 (
            .O(N__39690),
            .I(\nx.n10970 ));
    CascadeMux I__8890 (
            .O(N__39687),
            .I(N__39684));
    InMux I__8889 (
            .O(N__39684),
            .I(N__39680));
    InMux I__8888 (
            .O(N__39683),
            .I(N__39677));
    LocalMux I__8887 (
            .O(N__39680),
            .I(N__39674));
    LocalMux I__8886 (
            .O(N__39677),
            .I(\nx.n2597 ));
    Odrv12 I__8885 (
            .O(N__39674),
            .I(\nx.n2597 ));
    CascadeMux I__8884 (
            .O(N__39669),
            .I(N__39666));
    InMux I__8883 (
            .O(N__39666),
            .I(N__39663));
    LocalMux I__8882 (
            .O(N__39663),
            .I(N__39660));
    Span4Mux_v I__8881 (
            .O(N__39660),
            .I(N__39657));
    Span4Mux_h I__8880 (
            .O(N__39657),
            .I(N__39654));
    Odrv4 I__8879 (
            .O(N__39654),
            .I(\nx.n2664 ));
    InMux I__8878 (
            .O(N__39651),
            .I(\nx.n10971 ));
    InMux I__8877 (
            .O(N__39648),
            .I(N__39645));
    LocalMux I__8876 (
            .O(N__39645),
            .I(N__39640));
    CascadeMux I__8875 (
            .O(N__39644),
            .I(N__39637));
    InMux I__8874 (
            .O(N__39643),
            .I(N__39634));
    Span4Mux_v I__8873 (
            .O(N__39640),
            .I(N__39631));
    InMux I__8872 (
            .O(N__39637),
            .I(N__39628));
    LocalMux I__8871 (
            .O(N__39634),
            .I(N__39625));
    Odrv4 I__8870 (
            .O(N__39631),
            .I(\nx.n2596 ));
    LocalMux I__8869 (
            .O(N__39628),
            .I(\nx.n2596 ));
    Odrv4 I__8868 (
            .O(N__39625),
            .I(\nx.n2596 ));
    CascadeMux I__8867 (
            .O(N__39618),
            .I(N__39615));
    InMux I__8866 (
            .O(N__39615),
            .I(N__39612));
    LocalMux I__8865 (
            .O(N__39612),
            .I(N__39609));
    Span4Mux_v I__8864 (
            .O(N__39609),
            .I(N__39606));
    Odrv4 I__8863 (
            .O(N__39606),
            .I(\nx.n2663 ));
    InMux I__8862 (
            .O(N__39603),
            .I(\nx.n10972 ));
    InMux I__8861 (
            .O(N__39600),
            .I(N__39596));
    CascadeMux I__8860 (
            .O(N__39599),
            .I(N__39593));
    LocalMux I__8859 (
            .O(N__39596),
            .I(N__39589));
    InMux I__8858 (
            .O(N__39593),
            .I(N__39586));
    InMux I__8857 (
            .O(N__39592),
            .I(N__39583));
    Span4Mux_h I__8856 (
            .O(N__39589),
            .I(N__39580));
    LocalMux I__8855 (
            .O(N__39586),
            .I(N__39577));
    LocalMux I__8854 (
            .O(N__39583),
            .I(N__39574));
    Odrv4 I__8853 (
            .O(N__39580),
            .I(\nx.n2595 ));
    Odrv4 I__8852 (
            .O(N__39577),
            .I(\nx.n2595 ));
    Odrv12 I__8851 (
            .O(N__39574),
            .I(\nx.n2595 ));
    InMux I__8850 (
            .O(N__39567),
            .I(N__39564));
    LocalMux I__8849 (
            .O(N__39564),
            .I(N__39561));
    Span4Mux_h I__8848 (
            .O(N__39561),
            .I(N__39558));
    Span4Mux_h I__8847 (
            .O(N__39558),
            .I(N__39555));
    Odrv4 I__8846 (
            .O(N__39555),
            .I(\nx.n2662 ));
    InMux I__8845 (
            .O(N__39552),
            .I(\nx.n10973 ));
    InMux I__8844 (
            .O(N__39549),
            .I(N__39546));
    LocalMux I__8843 (
            .O(N__39546),
            .I(N__39542));
    CascadeMux I__8842 (
            .O(N__39545),
            .I(N__39539));
    Span4Mux_h I__8841 (
            .O(N__39542),
            .I(N__39535));
    InMux I__8840 (
            .O(N__39539),
            .I(N__39532));
    InMux I__8839 (
            .O(N__39538),
            .I(N__39529));
    Odrv4 I__8838 (
            .O(N__39535),
            .I(\nx.n2594 ));
    LocalMux I__8837 (
            .O(N__39532),
            .I(\nx.n2594 ));
    LocalMux I__8836 (
            .O(N__39529),
            .I(\nx.n2594 ));
    CascadeMux I__8835 (
            .O(N__39522),
            .I(N__39519));
    InMux I__8834 (
            .O(N__39519),
            .I(N__39516));
    LocalMux I__8833 (
            .O(N__39516),
            .I(N__39513));
    Span4Mux_h I__8832 (
            .O(N__39513),
            .I(N__39510));
    Span4Mux_h I__8831 (
            .O(N__39510),
            .I(N__39507));
    Odrv4 I__8830 (
            .O(N__39507),
            .I(\nx.n2661 ));
    InMux I__8829 (
            .O(N__39504),
            .I(bfn_16_23_0_));
    CascadeMux I__8828 (
            .O(N__39501),
            .I(N__39498));
    InMux I__8827 (
            .O(N__39498),
            .I(N__39495));
    LocalMux I__8826 (
            .O(N__39495),
            .I(N__39491));
    CascadeMux I__8825 (
            .O(N__39494),
            .I(N__39488));
    Span4Mux_v I__8824 (
            .O(N__39491),
            .I(N__39484));
    InMux I__8823 (
            .O(N__39488),
            .I(N__39481));
    InMux I__8822 (
            .O(N__39487),
            .I(N__39478));
    Odrv4 I__8821 (
            .O(N__39484),
            .I(\nx.n2593 ));
    LocalMux I__8820 (
            .O(N__39481),
            .I(\nx.n2593 ));
    LocalMux I__8819 (
            .O(N__39478),
            .I(\nx.n2593 ));
    InMux I__8818 (
            .O(N__39471),
            .I(N__39468));
    LocalMux I__8817 (
            .O(N__39468),
            .I(N__39465));
    Span4Mux_h I__8816 (
            .O(N__39465),
            .I(N__39462));
    Span4Mux_h I__8815 (
            .O(N__39462),
            .I(N__39459));
    Odrv4 I__8814 (
            .O(N__39459),
            .I(\nx.n2660 ));
    InMux I__8813 (
            .O(N__39456),
            .I(\nx.n10975 ));
    InMux I__8812 (
            .O(N__39453),
            .I(N__39449));
    CascadeMux I__8811 (
            .O(N__39452),
            .I(N__39446));
    LocalMux I__8810 (
            .O(N__39449),
            .I(N__39443));
    InMux I__8809 (
            .O(N__39446),
            .I(N__39440));
    Odrv12 I__8808 (
            .O(N__39443),
            .I(\nx.n2592 ));
    LocalMux I__8807 (
            .O(N__39440),
            .I(\nx.n2592 ));
    CascadeMux I__8806 (
            .O(N__39435),
            .I(N__39432));
    InMux I__8805 (
            .O(N__39432),
            .I(N__39429));
    LocalMux I__8804 (
            .O(N__39429),
            .I(N__39426));
    Span4Mux_v I__8803 (
            .O(N__39426),
            .I(N__39423));
    Span4Mux_h I__8802 (
            .O(N__39423),
            .I(N__39420));
    Odrv4 I__8801 (
            .O(N__39420),
            .I(\nx.n2659 ));
    InMux I__8800 (
            .O(N__39417),
            .I(\nx.n10976 ));
    CascadeMux I__8799 (
            .O(N__39414),
            .I(N__39411));
    InMux I__8798 (
            .O(N__39411),
            .I(N__39407));
    CascadeMux I__8797 (
            .O(N__39410),
            .I(N__39404));
    LocalMux I__8796 (
            .O(N__39407),
            .I(N__39401));
    InMux I__8795 (
            .O(N__39404),
            .I(N__39397));
    Span4Mux_h I__8794 (
            .O(N__39401),
            .I(N__39394));
    InMux I__8793 (
            .O(N__39400),
            .I(N__39391));
    LocalMux I__8792 (
            .O(N__39397),
            .I(\nx.n2591 ));
    Odrv4 I__8791 (
            .O(N__39394),
            .I(\nx.n2591 ));
    LocalMux I__8790 (
            .O(N__39391),
            .I(\nx.n2591 ));
    InMux I__8789 (
            .O(N__39384),
            .I(N__39381));
    LocalMux I__8788 (
            .O(N__39381),
            .I(N__39378));
    Odrv12 I__8787 (
            .O(N__39378),
            .I(\nx.n2658 ));
    InMux I__8786 (
            .O(N__39375),
            .I(\nx.n10977 ));
    InMux I__8785 (
            .O(N__39372),
            .I(N__39369));
    LocalMux I__8784 (
            .O(N__39369),
            .I(N__39365));
    CascadeMux I__8783 (
            .O(N__39368),
            .I(N__39362));
    Span4Mux_v I__8782 (
            .O(N__39365),
            .I(N__39359));
    InMux I__8781 (
            .O(N__39362),
            .I(N__39356));
    Odrv4 I__8780 (
            .O(N__39359),
            .I(\nx.n2606 ));
    LocalMux I__8779 (
            .O(N__39356),
            .I(\nx.n2606 ));
    InMux I__8778 (
            .O(N__39351),
            .I(N__39348));
    LocalMux I__8777 (
            .O(N__39348),
            .I(\nx.n2673 ));
    InMux I__8776 (
            .O(N__39345),
            .I(\nx.n10962 ));
    InMux I__8775 (
            .O(N__39342),
            .I(N__39339));
    LocalMux I__8774 (
            .O(N__39339),
            .I(N__39334));
    CascadeMux I__8773 (
            .O(N__39338),
            .I(N__39331));
    InMux I__8772 (
            .O(N__39337),
            .I(N__39328));
    Span4Mux_v I__8771 (
            .O(N__39334),
            .I(N__39325));
    InMux I__8770 (
            .O(N__39331),
            .I(N__39322));
    LocalMux I__8769 (
            .O(N__39328),
            .I(\nx.n2605 ));
    Odrv4 I__8768 (
            .O(N__39325),
            .I(\nx.n2605 ));
    LocalMux I__8767 (
            .O(N__39322),
            .I(\nx.n2605 ));
    InMux I__8766 (
            .O(N__39315),
            .I(N__39312));
    LocalMux I__8765 (
            .O(N__39312),
            .I(\nx.n2672 ));
    InMux I__8764 (
            .O(N__39309),
            .I(\nx.n10963 ));
    CascadeMux I__8763 (
            .O(N__39306),
            .I(N__39301));
    CascadeMux I__8762 (
            .O(N__39305),
            .I(N__39298));
    InMux I__8761 (
            .O(N__39304),
            .I(N__39295));
    InMux I__8760 (
            .O(N__39301),
            .I(N__39292));
    InMux I__8759 (
            .O(N__39298),
            .I(N__39289));
    LocalMux I__8758 (
            .O(N__39295),
            .I(N__39284));
    LocalMux I__8757 (
            .O(N__39292),
            .I(N__39284));
    LocalMux I__8756 (
            .O(N__39289),
            .I(N__39281));
    Span4Mux_h I__8755 (
            .O(N__39284),
            .I(N__39278));
    Odrv4 I__8754 (
            .O(N__39281),
            .I(\nx.n2604 ));
    Odrv4 I__8753 (
            .O(N__39278),
            .I(\nx.n2604 ));
    CascadeMux I__8752 (
            .O(N__39273),
            .I(N__39270));
    InMux I__8751 (
            .O(N__39270),
            .I(N__39267));
    LocalMux I__8750 (
            .O(N__39267),
            .I(N__39264));
    Odrv4 I__8749 (
            .O(N__39264),
            .I(\nx.n2671 ));
    InMux I__8748 (
            .O(N__39261),
            .I(\nx.n10964 ));
    CascadeMux I__8747 (
            .O(N__39258),
            .I(N__39255));
    InMux I__8746 (
            .O(N__39255),
            .I(N__39252));
    LocalMux I__8745 (
            .O(N__39252),
            .I(N__39248));
    InMux I__8744 (
            .O(N__39251),
            .I(N__39245));
    Span4Mux_v I__8743 (
            .O(N__39248),
            .I(N__39242));
    LocalMux I__8742 (
            .O(N__39245),
            .I(\nx.n2603 ));
    Odrv4 I__8741 (
            .O(N__39242),
            .I(\nx.n2603 ));
    InMux I__8740 (
            .O(N__39237),
            .I(N__39234));
    LocalMux I__8739 (
            .O(N__39234),
            .I(N__39231));
    Span4Mux_h I__8738 (
            .O(N__39231),
            .I(N__39228));
    Odrv4 I__8737 (
            .O(N__39228),
            .I(\nx.n2670 ));
    InMux I__8736 (
            .O(N__39225),
            .I(\nx.n10965 ));
    CascadeMux I__8735 (
            .O(N__39222),
            .I(N__39218));
    InMux I__8734 (
            .O(N__39221),
            .I(N__39215));
    InMux I__8733 (
            .O(N__39218),
            .I(N__39211));
    LocalMux I__8732 (
            .O(N__39215),
            .I(N__39208));
    InMux I__8731 (
            .O(N__39214),
            .I(N__39205));
    LocalMux I__8730 (
            .O(N__39211),
            .I(N__39202));
    Odrv4 I__8729 (
            .O(N__39208),
            .I(\nx.n2602 ));
    LocalMux I__8728 (
            .O(N__39205),
            .I(\nx.n2602 ));
    Odrv12 I__8727 (
            .O(N__39202),
            .I(\nx.n2602 ));
    InMux I__8726 (
            .O(N__39195),
            .I(N__39192));
    LocalMux I__8725 (
            .O(N__39192),
            .I(N__39189));
    Span4Mux_v I__8724 (
            .O(N__39189),
            .I(N__39186));
    Span4Mux_h I__8723 (
            .O(N__39186),
            .I(N__39183));
    Odrv4 I__8722 (
            .O(N__39183),
            .I(\nx.n2669 ));
    InMux I__8721 (
            .O(N__39180),
            .I(bfn_16_22_0_));
    CascadeMux I__8720 (
            .O(N__39177),
            .I(N__39174));
    InMux I__8719 (
            .O(N__39174),
            .I(N__39170));
    InMux I__8718 (
            .O(N__39173),
            .I(N__39166));
    LocalMux I__8717 (
            .O(N__39170),
            .I(N__39163));
    InMux I__8716 (
            .O(N__39169),
            .I(N__39160));
    LocalMux I__8715 (
            .O(N__39166),
            .I(\nx.n2601 ));
    Odrv4 I__8714 (
            .O(N__39163),
            .I(\nx.n2601 ));
    LocalMux I__8713 (
            .O(N__39160),
            .I(\nx.n2601 ));
    CascadeMux I__8712 (
            .O(N__39153),
            .I(N__39150));
    InMux I__8711 (
            .O(N__39150),
            .I(N__39147));
    LocalMux I__8710 (
            .O(N__39147),
            .I(N__39144));
    Odrv12 I__8709 (
            .O(N__39144),
            .I(\nx.n2668 ));
    InMux I__8708 (
            .O(N__39141),
            .I(\nx.n10967 ));
    InMux I__8707 (
            .O(N__39138),
            .I(N__39134));
    CascadeMux I__8706 (
            .O(N__39137),
            .I(N__39131));
    LocalMux I__8705 (
            .O(N__39134),
            .I(N__39128));
    InMux I__8704 (
            .O(N__39131),
            .I(N__39125));
    Span4Mux_h I__8703 (
            .O(N__39128),
            .I(N__39121));
    LocalMux I__8702 (
            .O(N__39125),
            .I(N__39118));
    InMux I__8701 (
            .O(N__39124),
            .I(N__39115));
    Odrv4 I__8700 (
            .O(N__39121),
            .I(\nx.n2600 ));
    Odrv4 I__8699 (
            .O(N__39118),
            .I(\nx.n2600 ));
    LocalMux I__8698 (
            .O(N__39115),
            .I(\nx.n2600 ));
    CascadeMux I__8697 (
            .O(N__39108),
            .I(N__39105));
    InMux I__8696 (
            .O(N__39105),
            .I(N__39102));
    LocalMux I__8695 (
            .O(N__39102),
            .I(N__39099));
    Span4Mux_v I__8694 (
            .O(N__39099),
            .I(N__39096));
    Span4Mux_h I__8693 (
            .O(N__39096),
            .I(N__39093));
    Odrv4 I__8692 (
            .O(N__39093),
            .I(\nx.n2667 ));
    InMux I__8691 (
            .O(N__39090),
            .I(\nx.n10968 ));
    CascadeMux I__8690 (
            .O(N__39087),
            .I(N__39083));
    InMux I__8689 (
            .O(N__39086),
            .I(N__39080));
    InMux I__8688 (
            .O(N__39083),
            .I(N__39076));
    LocalMux I__8687 (
            .O(N__39080),
            .I(N__39073));
    InMux I__8686 (
            .O(N__39079),
            .I(N__39070));
    LocalMux I__8685 (
            .O(N__39076),
            .I(N__39067));
    Span4Mux_v I__8684 (
            .O(N__39073),
            .I(N__39062));
    LocalMux I__8683 (
            .O(N__39070),
            .I(N__39062));
    Odrv4 I__8682 (
            .O(N__39067),
            .I(\nx.n2599 ));
    Odrv4 I__8681 (
            .O(N__39062),
            .I(\nx.n2599 ));
    InMux I__8680 (
            .O(N__39057),
            .I(N__39054));
    LocalMux I__8679 (
            .O(N__39054),
            .I(N__39051));
    Span4Mux_v I__8678 (
            .O(N__39051),
            .I(N__39048));
    Span4Mux_h I__8677 (
            .O(N__39048),
            .I(N__39045));
    Odrv4 I__8676 (
            .O(N__39045),
            .I(\nx.n2666 ));
    InMux I__8675 (
            .O(N__39042),
            .I(\nx.n10969 ));
    CascadeMux I__8674 (
            .O(N__39039),
            .I(n7_adj_840_cascade_));
    IoInMux I__8673 (
            .O(N__39036),
            .I(N__39033));
    LocalMux I__8672 (
            .O(N__39033),
            .I(N__39030));
    IoSpan4Mux I__8671 (
            .O(N__39030),
            .I(N__39027));
    Span4Mux_s2_v I__8670 (
            .O(N__39027),
            .I(N__39024));
    Sp12to4 I__8669 (
            .O(N__39024),
            .I(N__39021));
    Span12Mux_h I__8668 (
            .O(N__39021),
            .I(N__39016));
    InMux I__8667 (
            .O(N__39020),
            .I(N__39013));
    InMux I__8666 (
            .O(N__39019),
            .I(N__39010));
    Odrv12 I__8665 (
            .O(N__39016),
            .I(pin_out_0));
    LocalMux I__8664 (
            .O(N__39013),
            .I(pin_out_0));
    LocalMux I__8663 (
            .O(N__39010),
            .I(pin_out_0));
    InMux I__8662 (
            .O(N__39003),
            .I(N__39000));
    LocalMux I__8661 (
            .O(N__39000),
            .I(n8_adj_817));
    IoInMux I__8660 (
            .O(N__38997),
            .I(N__38994));
    LocalMux I__8659 (
            .O(N__38994),
            .I(N__38991));
    IoSpan4Mux I__8658 (
            .O(N__38991),
            .I(N__38988));
    Span4Mux_s2_v I__8657 (
            .O(N__38988),
            .I(N__38985));
    Sp12to4 I__8656 (
            .O(N__38985),
            .I(N__38982));
    Span12Mux_s8_v I__8655 (
            .O(N__38982),
            .I(N__38979));
    Span12Mux_h I__8654 (
            .O(N__38979),
            .I(N__38974));
    InMux I__8653 (
            .O(N__38978),
            .I(N__38969));
    InMux I__8652 (
            .O(N__38977),
            .I(N__38969));
    Odrv12 I__8651 (
            .O(N__38974),
            .I(pin_out_1));
    LocalMux I__8650 (
            .O(N__38969),
            .I(pin_out_1));
    InMux I__8649 (
            .O(N__38964),
            .I(N__38961));
    LocalMux I__8648 (
            .O(N__38961),
            .I(N__38958));
    Span12Mux_v I__8647 (
            .O(N__38958),
            .I(N__38955));
    Odrv12 I__8646 (
            .O(N__38955),
            .I(n11952));
    IoInMux I__8645 (
            .O(N__38952),
            .I(N__38949));
    LocalMux I__8644 (
            .O(N__38949),
            .I(N__38946));
    Span12Mux_s5_v I__8643 (
            .O(N__38946),
            .I(N__38943));
    Span12Mux_h I__8642 (
            .O(N__38943),
            .I(N__38939));
    InMux I__8641 (
            .O(N__38942),
            .I(N__38936));
    Odrv12 I__8640 (
            .O(N__38939),
            .I(pin_oe_8));
    LocalMux I__8639 (
            .O(N__38936),
            .I(pin_oe_8));
    InMux I__8638 (
            .O(N__38931),
            .I(N__38928));
    LocalMux I__8637 (
            .O(N__38928),
            .I(N__38924));
    InMux I__8636 (
            .O(N__38927),
            .I(N__38921));
    Span4Mux_v I__8635 (
            .O(N__38924),
            .I(N__38917));
    LocalMux I__8634 (
            .O(N__38921),
            .I(N__38914));
    InMux I__8633 (
            .O(N__38920),
            .I(N__38909));
    Span4Mux_h I__8632 (
            .O(N__38917),
            .I(N__38906));
    Span4Mux_v I__8631 (
            .O(N__38914),
            .I(N__38903));
    InMux I__8630 (
            .O(N__38913),
            .I(N__38900));
    InMux I__8629 (
            .O(N__38912),
            .I(N__38897));
    LocalMux I__8628 (
            .O(N__38909),
            .I(N__38890));
    Sp12to4 I__8627 (
            .O(N__38906),
            .I(N__38890));
    Sp12to4 I__8626 (
            .O(N__38903),
            .I(N__38890));
    LocalMux I__8625 (
            .O(N__38900),
            .I(\nx.bit_ctr_9 ));
    LocalMux I__8624 (
            .O(N__38897),
            .I(\nx.bit_ctr_9 ));
    Odrv12 I__8623 (
            .O(N__38890),
            .I(\nx.bit_ctr_9 ));
    InMux I__8622 (
            .O(N__38883),
            .I(N__38880));
    LocalMux I__8621 (
            .O(N__38880),
            .I(N__38877));
    Span4Mux_v I__8620 (
            .O(N__38877),
            .I(N__38874));
    Span4Mux_h I__8619 (
            .O(N__38874),
            .I(N__38871));
    Odrv4 I__8618 (
            .O(N__38871),
            .I(\nx.n2677 ));
    InMux I__8617 (
            .O(N__38868),
            .I(bfn_16_21_0_));
    InMux I__8616 (
            .O(N__38865),
            .I(N__38862));
    LocalMux I__8615 (
            .O(N__38862),
            .I(N__38858));
    CascadeMux I__8614 (
            .O(N__38861),
            .I(N__38855));
    Span4Mux_h I__8613 (
            .O(N__38858),
            .I(N__38852));
    InMux I__8612 (
            .O(N__38855),
            .I(N__38849));
    Odrv4 I__8611 (
            .O(N__38852),
            .I(\nx.n2609 ));
    LocalMux I__8610 (
            .O(N__38849),
            .I(\nx.n2609 ));
    InMux I__8609 (
            .O(N__38844),
            .I(N__38841));
    LocalMux I__8608 (
            .O(N__38841),
            .I(N__38838));
    Span4Mux_h I__8607 (
            .O(N__38838),
            .I(N__38835));
    Odrv4 I__8606 (
            .O(N__38835),
            .I(\nx.n2676 ));
    InMux I__8605 (
            .O(N__38832),
            .I(\nx.n10959 ));
    InMux I__8604 (
            .O(N__38829),
            .I(N__38826));
    LocalMux I__8603 (
            .O(N__38826),
            .I(N__38822));
    CascadeMux I__8602 (
            .O(N__38825),
            .I(N__38818));
    Span4Mux_h I__8601 (
            .O(N__38822),
            .I(N__38815));
    InMux I__8600 (
            .O(N__38821),
            .I(N__38812));
    InMux I__8599 (
            .O(N__38818),
            .I(N__38809));
    Odrv4 I__8598 (
            .O(N__38815),
            .I(\nx.n2608 ));
    LocalMux I__8597 (
            .O(N__38812),
            .I(\nx.n2608 ));
    LocalMux I__8596 (
            .O(N__38809),
            .I(\nx.n2608 ));
    CascadeMux I__8595 (
            .O(N__38802),
            .I(N__38799));
    InMux I__8594 (
            .O(N__38799),
            .I(N__38796));
    LocalMux I__8593 (
            .O(N__38796),
            .I(N__38793));
    Span4Mux_v I__8592 (
            .O(N__38793),
            .I(N__38790));
    Odrv4 I__8591 (
            .O(N__38790),
            .I(\nx.n2675 ));
    InMux I__8590 (
            .O(N__38787),
            .I(\nx.n10960 ));
    InMux I__8589 (
            .O(N__38784),
            .I(N__38781));
    LocalMux I__8588 (
            .O(N__38781),
            .I(N__38777));
    CascadeMux I__8587 (
            .O(N__38780),
            .I(N__38774));
    Span4Mux_h I__8586 (
            .O(N__38777),
            .I(N__38770));
    InMux I__8585 (
            .O(N__38774),
            .I(N__38767));
    InMux I__8584 (
            .O(N__38773),
            .I(N__38764));
    Odrv4 I__8583 (
            .O(N__38770),
            .I(\nx.n2607 ));
    LocalMux I__8582 (
            .O(N__38767),
            .I(\nx.n2607 ));
    LocalMux I__8581 (
            .O(N__38764),
            .I(\nx.n2607 ));
    CascadeMux I__8580 (
            .O(N__38757),
            .I(N__38754));
    InMux I__8579 (
            .O(N__38754),
            .I(N__38751));
    LocalMux I__8578 (
            .O(N__38751),
            .I(N__38748));
    Span4Mux_v I__8577 (
            .O(N__38748),
            .I(N__38745));
    Span4Mux_h I__8576 (
            .O(N__38745),
            .I(N__38742));
    Odrv4 I__8575 (
            .O(N__38742),
            .I(\nx.n2674 ));
    InMux I__8574 (
            .O(N__38739),
            .I(\nx.n10961 ));
    CascadeMux I__8573 (
            .O(N__38736),
            .I(n9488_cascade_));
    CascadeMux I__8572 (
            .O(N__38733),
            .I(n7_adj_818_cascade_));
    CascadeMux I__8571 (
            .O(N__38730),
            .I(N__38727));
    InMux I__8570 (
            .O(N__38727),
            .I(N__38724));
    LocalMux I__8569 (
            .O(N__38724),
            .I(n7_adj_821));
    IoInMux I__8568 (
            .O(N__38721),
            .I(N__38718));
    LocalMux I__8567 (
            .O(N__38718),
            .I(N__38715));
    Span12Mux_s3_h I__8566 (
            .O(N__38715),
            .I(N__38712));
    Span12Mux_v I__8565 (
            .O(N__38712),
            .I(N__38708));
    InMux I__8564 (
            .O(N__38711),
            .I(N__38704));
    Span12Mux_h I__8563 (
            .O(N__38708),
            .I(N__38701));
    InMux I__8562 (
            .O(N__38707),
            .I(N__38698));
    LocalMux I__8561 (
            .O(N__38704),
            .I(N__38695));
    Odrv12 I__8560 (
            .O(N__38701),
            .I(pin_out_3));
    LocalMux I__8559 (
            .O(N__38698),
            .I(pin_out_3));
    Odrv4 I__8558 (
            .O(N__38695),
            .I(pin_out_3));
    IoInMux I__8557 (
            .O(N__38688),
            .I(N__38685));
    LocalMux I__8556 (
            .O(N__38685),
            .I(N__38682));
    Span4Mux_s3_h I__8555 (
            .O(N__38682),
            .I(N__38679));
    Span4Mux_h I__8554 (
            .O(N__38679),
            .I(N__38676));
    Span4Mux_h I__8553 (
            .O(N__38676),
            .I(N__38673));
    Span4Mux_h I__8552 (
            .O(N__38673),
            .I(N__38668));
    InMux I__8551 (
            .O(N__38672),
            .I(N__38665));
    InMux I__8550 (
            .O(N__38671),
            .I(N__38662));
    Odrv4 I__8549 (
            .O(N__38668),
            .I(pin_out_2));
    LocalMux I__8548 (
            .O(N__38665),
            .I(pin_out_2));
    LocalMux I__8547 (
            .O(N__38662),
            .I(pin_out_2));
    CascadeMux I__8546 (
            .O(N__38655),
            .I(n13355_cascade_));
    InMux I__8545 (
            .O(N__38652),
            .I(N__38649));
    LocalMux I__8544 (
            .O(N__38649),
            .I(n13354));
    InMux I__8543 (
            .O(N__38646),
            .I(N__38643));
    LocalMux I__8542 (
            .O(N__38643),
            .I(n9));
    CascadeMux I__8541 (
            .O(N__38640),
            .I(n9_cascade_));
    CascadeMux I__8540 (
            .O(N__38637),
            .I(n8_adj_820_cascade_));
    CascadeMux I__8539 (
            .O(N__38634),
            .I(n6_adj_805_cascade_));
    InMux I__8538 (
            .O(N__38631),
            .I(N__38628));
    LocalMux I__8537 (
            .O(N__38628),
            .I(N__38624));
    InMux I__8536 (
            .O(N__38627),
            .I(N__38621));
    Odrv12 I__8535 (
            .O(N__38624),
            .I(n1788));
    LocalMux I__8534 (
            .O(N__38621),
            .I(n1788));
    IoInMux I__8533 (
            .O(N__38616),
            .I(N__38613));
    LocalMux I__8532 (
            .O(N__38613),
            .I(N__38610));
    Span4Mux_s3_v I__8531 (
            .O(N__38610),
            .I(N__38607));
    Span4Mux_h I__8530 (
            .O(N__38607),
            .I(N__38604));
    Span4Mux_v I__8529 (
            .O(N__38604),
            .I(N__38600));
    InMux I__8528 (
            .O(N__38603),
            .I(N__38597));
    Odrv4 I__8527 (
            .O(N__38600),
            .I(pin_oe_22));
    LocalMux I__8526 (
            .O(N__38597),
            .I(pin_oe_22));
    InMux I__8525 (
            .O(N__38592),
            .I(N__38588));
    CascadeMux I__8524 (
            .O(N__38591),
            .I(N__38585));
    LocalMux I__8523 (
            .O(N__38588),
            .I(N__38582));
    InMux I__8522 (
            .O(N__38585),
            .I(N__38579));
    Span4Mux_v I__8521 (
            .O(N__38582),
            .I(N__38574));
    LocalMux I__8520 (
            .O(N__38579),
            .I(N__38574));
    Span4Mux_h I__8519 (
            .O(N__38574),
            .I(N__38570));
    InMux I__8518 (
            .O(N__38573),
            .I(N__38567));
    Odrv4 I__8517 (
            .O(N__38570),
            .I(\nx.n2392 ));
    LocalMux I__8516 (
            .O(N__38567),
            .I(\nx.n2392 ));
    CascadeMux I__8515 (
            .O(N__38562),
            .I(N__38559));
    InMux I__8514 (
            .O(N__38559),
            .I(N__38556));
    LocalMux I__8513 (
            .O(N__38556),
            .I(\nx.n2459 ));
    CascadeMux I__8512 (
            .O(N__38553),
            .I(\nx.n2491_cascade_ ));
    InMux I__8511 (
            .O(N__38550),
            .I(N__38547));
    LocalMux I__8510 (
            .O(N__38547),
            .I(N__38544));
    Odrv12 I__8509 (
            .O(N__38544),
            .I(\nx.n33_adj_767 ));
    InMux I__8508 (
            .O(N__38541),
            .I(N__38538));
    LocalMux I__8507 (
            .O(N__38538),
            .I(\nx.n2460 ));
    CascadeMux I__8506 (
            .O(N__38535),
            .I(N__38532));
    InMux I__8505 (
            .O(N__38532),
            .I(N__38528));
    CascadeMux I__8504 (
            .O(N__38531),
            .I(N__38525));
    LocalMux I__8503 (
            .O(N__38528),
            .I(N__38522));
    InMux I__8502 (
            .O(N__38525),
            .I(N__38519));
    Span4Mux_h I__8501 (
            .O(N__38522),
            .I(N__38513));
    LocalMux I__8500 (
            .O(N__38519),
            .I(N__38513));
    InMux I__8499 (
            .O(N__38518),
            .I(N__38510));
    Odrv4 I__8498 (
            .O(N__38513),
            .I(\nx.n2393 ));
    LocalMux I__8497 (
            .O(N__38510),
            .I(\nx.n2393 ));
    CascadeMux I__8496 (
            .O(N__38505),
            .I(N__38493));
    CascadeMux I__8495 (
            .O(N__38504),
            .I(N__38489));
    InMux I__8494 (
            .O(N__38503),
            .I(N__38482));
    InMux I__8493 (
            .O(N__38502),
            .I(N__38482));
    InMux I__8492 (
            .O(N__38501),
            .I(N__38479));
    InMux I__8491 (
            .O(N__38500),
            .I(N__38475));
    CascadeMux I__8490 (
            .O(N__38499),
            .I(N__38471));
    CascadeMux I__8489 (
            .O(N__38498),
            .I(N__38466));
    CascadeMux I__8488 (
            .O(N__38497),
            .I(N__38462));
    CascadeMux I__8487 (
            .O(N__38496),
            .I(N__38457));
    InMux I__8486 (
            .O(N__38493),
            .I(N__38445));
    InMux I__8485 (
            .O(N__38492),
            .I(N__38445));
    InMux I__8484 (
            .O(N__38489),
            .I(N__38445));
    InMux I__8483 (
            .O(N__38488),
            .I(N__38445));
    InMux I__8482 (
            .O(N__38487),
            .I(N__38445));
    LocalMux I__8481 (
            .O(N__38482),
            .I(N__38440));
    LocalMux I__8480 (
            .O(N__38479),
            .I(N__38440));
    InMux I__8479 (
            .O(N__38478),
            .I(N__38437));
    LocalMux I__8478 (
            .O(N__38475),
            .I(N__38434));
    InMux I__8477 (
            .O(N__38474),
            .I(N__38431));
    InMux I__8476 (
            .O(N__38471),
            .I(N__38424));
    InMux I__8475 (
            .O(N__38470),
            .I(N__38424));
    InMux I__8474 (
            .O(N__38469),
            .I(N__38424));
    InMux I__8473 (
            .O(N__38466),
            .I(N__38419));
    InMux I__8472 (
            .O(N__38465),
            .I(N__38419));
    InMux I__8471 (
            .O(N__38462),
            .I(N__38408));
    InMux I__8470 (
            .O(N__38461),
            .I(N__38408));
    InMux I__8469 (
            .O(N__38460),
            .I(N__38408));
    InMux I__8468 (
            .O(N__38457),
            .I(N__38408));
    InMux I__8467 (
            .O(N__38456),
            .I(N__38408));
    LocalMux I__8466 (
            .O(N__38445),
            .I(\nx.n2423 ));
    Odrv4 I__8465 (
            .O(N__38440),
            .I(\nx.n2423 ));
    LocalMux I__8464 (
            .O(N__38437),
            .I(\nx.n2423 ));
    Odrv4 I__8463 (
            .O(N__38434),
            .I(\nx.n2423 ));
    LocalMux I__8462 (
            .O(N__38431),
            .I(\nx.n2423 ));
    LocalMux I__8461 (
            .O(N__38424),
            .I(\nx.n2423 ));
    LocalMux I__8460 (
            .O(N__38419),
            .I(\nx.n2423 ));
    LocalMux I__8459 (
            .O(N__38408),
            .I(\nx.n2423 ));
    SRMux I__8458 (
            .O(N__38391),
            .I(N__38387));
    SRMux I__8457 (
            .O(N__38390),
            .I(N__38384));
    LocalMux I__8456 (
            .O(N__38387),
            .I(N__38379));
    LocalMux I__8455 (
            .O(N__38384),
            .I(N__38379));
    Span4Mux_v I__8454 (
            .O(N__38379),
            .I(N__38376));
    Span4Mux_h I__8453 (
            .O(N__38376),
            .I(N__38373));
    Odrv4 I__8452 (
            .O(N__38373),
            .I(n7992));
    InMux I__8451 (
            .O(N__38370),
            .I(N__38367));
    LocalMux I__8450 (
            .O(N__38367),
            .I(n7602));
    IoInMux I__8449 (
            .O(N__38364),
            .I(N__38361));
    LocalMux I__8448 (
            .O(N__38361),
            .I(N__38358));
    IoSpan4Mux I__8447 (
            .O(N__38358),
            .I(N__38355));
    Span4Mux_s0_h I__8446 (
            .O(N__38355),
            .I(N__38352));
    Sp12to4 I__8445 (
            .O(N__38352),
            .I(N__38349));
    Span12Mux_s11_h I__8444 (
            .O(N__38349),
            .I(N__38346));
    Span12Mux_v I__8443 (
            .O(N__38346),
            .I(N__38342));
    InMux I__8442 (
            .O(N__38345),
            .I(N__38339));
    Odrv12 I__8441 (
            .O(N__38342),
            .I(pin_oe_11));
    LocalMux I__8440 (
            .O(N__38339),
            .I(pin_oe_11));
    InMux I__8439 (
            .O(N__38334),
            .I(N__38331));
    LocalMux I__8438 (
            .O(N__38331),
            .I(\nx.n2476 ));
    CascadeMux I__8437 (
            .O(N__38328),
            .I(N__38325));
    InMux I__8436 (
            .O(N__38325),
            .I(N__38322));
    LocalMux I__8435 (
            .O(N__38322),
            .I(N__38318));
    CascadeMux I__8434 (
            .O(N__38321),
            .I(N__38314));
    Span4Mux_h I__8433 (
            .O(N__38318),
            .I(N__38311));
    InMux I__8432 (
            .O(N__38317),
            .I(N__38308));
    InMux I__8431 (
            .O(N__38314),
            .I(N__38305));
    Odrv4 I__8430 (
            .O(N__38311),
            .I(\nx.n2409 ));
    LocalMux I__8429 (
            .O(N__38308),
            .I(\nx.n2409 ));
    LocalMux I__8428 (
            .O(N__38305),
            .I(\nx.n2409 ));
    InMux I__8427 (
            .O(N__38298),
            .I(N__38294));
    CascadeMux I__8426 (
            .O(N__38297),
            .I(N__38291));
    LocalMux I__8425 (
            .O(N__38294),
            .I(N__38287));
    InMux I__8424 (
            .O(N__38291),
            .I(N__38284));
    InMux I__8423 (
            .O(N__38290),
            .I(N__38281));
    Span4Mux_h I__8422 (
            .O(N__38287),
            .I(N__38278));
    LocalMux I__8421 (
            .O(N__38284),
            .I(N__38273));
    LocalMux I__8420 (
            .O(N__38281),
            .I(N__38273));
    Odrv4 I__8419 (
            .O(N__38278),
            .I(\nx.n2400 ));
    Odrv12 I__8418 (
            .O(N__38273),
            .I(\nx.n2400 ));
    CascadeMux I__8417 (
            .O(N__38268),
            .I(N__38265));
    InMux I__8416 (
            .O(N__38265),
            .I(N__38262));
    LocalMux I__8415 (
            .O(N__38262),
            .I(\nx.n2467 ));
    CascadeMux I__8414 (
            .O(N__38259),
            .I(N__38255));
    InMux I__8413 (
            .O(N__38258),
            .I(N__38251));
    InMux I__8412 (
            .O(N__38255),
            .I(N__38248));
    InMux I__8411 (
            .O(N__38254),
            .I(N__38245));
    LocalMux I__8410 (
            .O(N__38251),
            .I(N__38242));
    LocalMux I__8409 (
            .O(N__38248),
            .I(N__38239));
    LocalMux I__8408 (
            .O(N__38245),
            .I(N__38236));
    Odrv4 I__8407 (
            .O(N__38242),
            .I(\nx.n2396 ));
    Odrv4 I__8406 (
            .O(N__38239),
            .I(\nx.n2396 ));
    Odrv12 I__8405 (
            .O(N__38236),
            .I(\nx.n2396 ));
    InMux I__8404 (
            .O(N__38229),
            .I(N__38226));
    LocalMux I__8403 (
            .O(N__38226),
            .I(N__38223));
    Odrv4 I__8402 (
            .O(N__38223),
            .I(\nx.n2463 ));
    CascadeMux I__8401 (
            .O(N__38220),
            .I(\nx.n2495_cascade_ ));
    InMux I__8400 (
            .O(N__38217),
            .I(N__38214));
    LocalMux I__8399 (
            .O(N__38214),
            .I(N__38211));
    Odrv4 I__8398 (
            .O(N__38211),
            .I(\nx.n34_adj_758 ));
    InMux I__8397 (
            .O(N__38208),
            .I(N__38205));
    LocalMux I__8396 (
            .O(N__38205),
            .I(N__38201));
    CascadeMux I__8395 (
            .O(N__38204),
            .I(N__38198));
    Span4Mux_h I__8394 (
            .O(N__38201),
            .I(N__38195));
    InMux I__8393 (
            .O(N__38198),
            .I(N__38192));
    Odrv4 I__8392 (
            .O(N__38195),
            .I(\nx.n2398 ));
    LocalMux I__8391 (
            .O(N__38192),
            .I(\nx.n2398 ));
    InMux I__8390 (
            .O(N__38187),
            .I(N__38184));
    LocalMux I__8389 (
            .O(N__38184),
            .I(\nx.n2465 ));
    InMux I__8388 (
            .O(N__38181),
            .I(N__38177));
    CascadeMux I__8387 (
            .O(N__38180),
            .I(N__38174));
    LocalMux I__8386 (
            .O(N__38177),
            .I(N__38170));
    InMux I__8385 (
            .O(N__38174),
            .I(N__38167));
    InMux I__8384 (
            .O(N__38173),
            .I(N__38164));
    Odrv4 I__8383 (
            .O(N__38170),
            .I(\nx.n2395 ));
    LocalMux I__8382 (
            .O(N__38167),
            .I(\nx.n2395 ));
    LocalMux I__8381 (
            .O(N__38164),
            .I(\nx.n2395 ));
    CascadeMux I__8380 (
            .O(N__38157),
            .I(N__38154));
    InMux I__8379 (
            .O(N__38154),
            .I(N__38151));
    LocalMux I__8378 (
            .O(N__38151),
            .I(\nx.n2462 ));
    CascadeMux I__8377 (
            .O(N__38148),
            .I(N__38144));
    InMux I__8376 (
            .O(N__38147),
            .I(N__38140));
    InMux I__8375 (
            .O(N__38144),
            .I(N__38137));
    InMux I__8374 (
            .O(N__38143),
            .I(N__38134));
    LocalMux I__8373 (
            .O(N__38140),
            .I(N__38131));
    LocalMux I__8372 (
            .O(N__38137),
            .I(N__38128));
    LocalMux I__8371 (
            .O(N__38134),
            .I(N__38125));
    Odrv4 I__8370 (
            .O(N__38131),
            .I(\nx.n2397 ));
    Odrv4 I__8369 (
            .O(N__38128),
            .I(\nx.n2397 ));
    Odrv12 I__8368 (
            .O(N__38125),
            .I(\nx.n2397 ));
    CascadeMux I__8367 (
            .O(N__38118),
            .I(N__38115));
    InMux I__8366 (
            .O(N__38115),
            .I(N__38112));
    LocalMux I__8365 (
            .O(N__38112),
            .I(\nx.n2464 ));
    CascadeMux I__8364 (
            .O(N__38109),
            .I(\nx.n2496_cascade_ ));
    InMux I__8363 (
            .O(N__38106),
            .I(N__38101));
    CascadeMux I__8362 (
            .O(N__38105),
            .I(N__38098));
    InMux I__8361 (
            .O(N__38104),
            .I(N__38095));
    LocalMux I__8360 (
            .O(N__38101),
            .I(N__38092));
    InMux I__8359 (
            .O(N__38098),
            .I(N__38089));
    LocalMux I__8358 (
            .O(N__38095),
            .I(N__38086));
    Odrv4 I__8357 (
            .O(N__38092),
            .I(\nx.n2394 ));
    LocalMux I__8356 (
            .O(N__38089),
            .I(\nx.n2394 ));
    Odrv12 I__8355 (
            .O(N__38086),
            .I(\nx.n2394 ));
    CascadeMux I__8354 (
            .O(N__38079),
            .I(N__38076));
    InMux I__8353 (
            .O(N__38076),
            .I(N__38073));
    LocalMux I__8352 (
            .O(N__38073),
            .I(\nx.n2461 ));
    CascadeMux I__8351 (
            .O(N__38070),
            .I(\nx.n2592_cascade_ ));
    InMux I__8350 (
            .O(N__38067),
            .I(N__38064));
    LocalMux I__8349 (
            .O(N__38064),
            .I(\nx.n35 ));
    InMux I__8348 (
            .O(N__38061),
            .I(N__38058));
    LocalMux I__8347 (
            .O(N__38058),
            .I(N__38055));
    Span4Mux_v I__8346 (
            .O(N__38055),
            .I(N__38051));
    InMux I__8345 (
            .O(N__38054),
            .I(N__38048));
    Span4Mux_h I__8344 (
            .O(N__38051),
            .I(N__38043));
    LocalMux I__8343 (
            .O(N__38048),
            .I(N__38043));
    Odrv4 I__8342 (
            .O(N__38043),
            .I(\nx.n2391 ));
    InMux I__8341 (
            .O(N__38040),
            .I(N__38037));
    LocalMux I__8340 (
            .O(N__38037),
            .I(N__38034));
    Odrv4 I__8339 (
            .O(N__38034),
            .I(\nx.n2458 ));
    CascadeMux I__8338 (
            .O(N__38031),
            .I(\nx.n2490_cascade_ ));
    InMux I__8337 (
            .O(N__38028),
            .I(N__38025));
    LocalMux I__8336 (
            .O(N__38025),
            .I(\nx.n22_adj_755 ));
    InMux I__8335 (
            .O(N__38022),
            .I(N__38018));
    CascadeMux I__8334 (
            .O(N__38021),
            .I(N__38005));
    LocalMux I__8333 (
            .O(N__38018),
            .I(N__38001));
    CascadeMux I__8332 (
            .O(N__38017),
            .I(N__37996));
    CascadeMux I__8331 (
            .O(N__38016),
            .I(N__37992));
    CascadeMux I__8330 (
            .O(N__38015),
            .I(N__37989));
    InMux I__8329 (
            .O(N__38014),
            .I(N__37978));
    InMux I__8328 (
            .O(N__38013),
            .I(N__37978));
    InMux I__8327 (
            .O(N__38012),
            .I(N__37978));
    InMux I__8326 (
            .O(N__38011),
            .I(N__37978));
    CascadeMux I__8325 (
            .O(N__38010),
            .I(N__37975));
    CascadeMux I__8324 (
            .O(N__38009),
            .I(N__37972));
    CascadeMux I__8323 (
            .O(N__38008),
            .I(N__37969));
    InMux I__8322 (
            .O(N__38005),
            .I(N__37964));
    InMux I__8321 (
            .O(N__38004),
            .I(N__37961));
    Span4Mux_h I__8320 (
            .O(N__38001),
            .I(N__37958));
    InMux I__8319 (
            .O(N__38000),
            .I(N__37949));
    InMux I__8318 (
            .O(N__37999),
            .I(N__37949));
    InMux I__8317 (
            .O(N__37996),
            .I(N__37949));
    InMux I__8316 (
            .O(N__37995),
            .I(N__37949));
    InMux I__8315 (
            .O(N__37992),
            .I(N__37944));
    InMux I__8314 (
            .O(N__37989),
            .I(N__37944));
    InMux I__8313 (
            .O(N__37988),
            .I(N__37939));
    InMux I__8312 (
            .O(N__37987),
            .I(N__37939));
    LocalMux I__8311 (
            .O(N__37978),
            .I(N__37936));
    InMux I__8310 (
            .O(N__37975),
            .I(N__37925));
    InMux I__8309 (
            .O(N__37972),
            .I(N__37925));
    InMux I__8308 (
            .O(N__37969),
            .I(N__37925));
    InMux I__8307 (
            .O(N__37968),
            .I(N__37925));
    InMux I__8306 (
            .O(N__37967),
            .I(N__37925));
    LocalMux I__8305 (
            .O(N__37964),
            .I(N__37920));
    LocalMux I__8304 (
            .O(N__37961),
            .I(N__37920));
    Odrv4 I__8303 (
            .O(N__37958),
            .I(\nx.n2324 ));
    LocalMux I__8302 (
            .O(N__37949),
            .I(\nx.n2324 ));
    LocalMux I__8301 (
            .O(N__37944),
            .I(\nx.n2324 ));
    LocalMux I__8300 (
            .O(N__37939),
            .I(\nx.n2324 ));
    Odrv4 I__8299 (
            .O(N__37936),
            .I(\nx.n2324 ));
    LocalMux I__8298 (
            .O(N__37925),
            .I(\nx.n2324 ));
    Odrv4 I__8297 (
            .O(N__37920),
            .I(\nx.n2324 ));
    CascadeMux I__8296 (
            .O(N__37905),
            .I(N__37902));
    InMux I__8295 (
            .O(N__37902),
            .I(N__37899));
    LocalMux I__8294 (
            .O(N__37899),
            .I(N__37893));
    InMux I__8293 (
            .O(N__37898),
            .I(N__37890));
    CascadeMux I__8292 (
            .O(N__37897),
            .I(N__37887));
    InMux I__8291 (
            .O(N__37896),
            .I(N__37884));
    Span4Mux_h I__8290 (
            .O(N__37893),
            .I(N__37879));
    LocalMux I__8289 (
            .O(N__37890),
            .I(N__37879));
    InMux I__8288 (
            .O(N__37887),
            .I(N__37876));
    LocalMux I__8287 (
            .O(N__37884),
            .I(\nx.n2307 ));
    Odrv4 I__8286 (
            .O(N__37879),
            .I(\nx.n2307 ));
    LocalMux I__8285 (
            .O(N__37876),
            .I(\nx.n2307 ));
    InMux I__8284 (
            .O(N__37869),
            .I(N__37866));
    LocalMux I__8283 (
            .O(N__37866),
            .I(\nx.n13321 ));
    CascadeMux I__8282 (
            .O(N__37863),
            .I(\nx.n2505_cascade_ ));
    CascadeMux I__8281 (
            .O(N__37860),
            .I(\nx.n2606_cascade_ ));
    CascadeMux I__8280 (
            .O(N__37857),
            .I(N__37853));
    InMux I__8279 (
            .O(N__37856),
            .I(N__37850));
    InMux I__8278 (
            .O(N__37853),
            .I(N__37847));
    LocalMux I__8277 (
            .O(N__37850),
            .I(N__37843));
    LocalMux I__8276 (
            .O(N__37847),
            .I(N__37840));
    CascadeMux I__8275 (
            .O(N__37846),
            .I(N__37837));
    Span4Mux_v I__8274 (
            .O(N__37843),
            .I(N__37832));
    Span4Mux_h I__8273 (
            .O(N__37840),
            .I(N__37832));
    InMux I__8272 (
            .O(N__37837),
            .I(N__37829));
    Span4Mux_h I__8271 (
            .O(N__37832),
            .I(N__37826));
    LocalMux I__8270 (
            .O(N__37829),
            .I(\nx.n2705 ));
    Odrv4 I__8269 (
            .O(N__37826),
            .I(\nx.n2705 ));
    CascadeMux I__8268 (
            .O(N__37821),
            .I(N__37818));
    InMux I__8267 (
            .O(N__37818),
            .I(N__37814));
    InMux I__8266 (
            .O(N__37817),
            .I(N__37811));
    LocalMux I__8265 (
            .O(N__37814),
            .I(N__37808));
    LocalMux I__8264 (
            .O(N__37811),
            .I(N__37805));
    Span4Mux_h I__8263 (
            .O(N__37808),
            .I(N__37801));
    Span4Mux_h I__8262 (
            .O(N__37805),
            .I(N__37798));
    InMux I__8261 (
            .O(N__37804),
            .I(N__37795));
    Span4Mux_h I__8260 (
            .O(N__37801),
            .I(N__37792));
    Odrv4 I__8259 (
            .O(N__37798),
            .I(\nx.n2704 ));
    LocalMux I__8258 (
            .O(N__37795),
            .I(\nx.n2704 ));
    Odrv4 I__8257 (
            .O(N__37792),
            .I(\nx.n2704 ));
    CascadeMux I__8256 (
            .O(N__37785),
            .I(\nx.n37_adj_772_cascade_ ));
    InMux I__8255 (
            .O(N__37782),
            .I(N__37779));
    LocalMux I__8254 (
            .O(N__37779),
            .I(\nx.n39_adj_773 ));
    CascadeMux I__8253 (
            .O(N__37776),
            .I(\nx.n2522_cascade_ ));
    InMux I__8252 (
            .O(N__37773),
            .I(N__37770));
    LocalMux I__8251 (
            .O(N__37770),
            .I(N__37767));
    Span4Mux_h I__8250 (
            .O(N__37767),
            .I(N__37763));
    InMux I__8249 (
            .O(N__37766),
            .I(N__37759));
    Span4Mux_v I__8248 (
            .O(N__37763),
            .I(N__37756));
    InMux I__8247 (
            .O(N__37762),
            .I(N__37753));
    LocalMux I__8246 (
            .O(N__37759),
            .I(N__37750));
    Odrv4 I__8245 (
            .O(N__37756),
            .I(\nx.n2793 ));
    LocalMux I__8244 (
            .O(N__37753),
            .I(\nx.n2793 ));
    Odrv12 I__8243 (
            .O(N__37750),
            .I(\nx.n2793 ));
    CascadeMux I__8242 (
            .O(N__37743),
            .I(N__37740));
    InMux I__8241 (
            .O(N__37740),
            .I(N__37737));
    LocalMux I__8240 (
            .O(N__37737),
            .I(N__37734));
    Span4Mux_h I__8239 (
            .O(N__37734),
            .I(N__37731));
    Span4Mux_h I__8238 (
            .O(N__37731),
            .I(N__37728));
    Odrv4 I__8237 (
            .O(N__37728),
            .I(\nx.n2860 ));
    CascadeMux I__8236 (
            .O(N__37725),
            .I(N__37722));
    InMux I__8235 (
            .O(N__37722),
            .I(N__37719));
    LocalMux I__8234 (
            .O(N__37719),
            .I(N__37715));
    CascadeMux I__8233 (
            .O(N__37718),
            .I(N__37711));
    Span4Mux_h I__8232 (
            .O(N__37715),
            .I(N__37708));
    InMux I__8231 (
            .O(N__37714),
            .I(N__37705));
    InMux I__8230 (
            .O(N__37711),
            .I(N__37702));
    Odrv4 I__8229 (
            .O(N__37708),
            .I(\nx.n2892 ));
    LocalMux I__8228 (
            .O(N__37705),
            .I(\nx.n2892 ));
    LocalMux I__8227 (
            .O(N__37702),
            .I(\nx.n2892 ));
    CascadeMux I__8226 (
            .O(N__37695),
            .I(N__37692));
    InMux I__8225 (
            .O(N__37692),
            .I(N__37689));
    LocalMux I__8224 (
            .O(N__37689),
            .I(\nx.n2960 ));
    InMux I__8223 (
            .O(N__37686),
            .I(N__37682));
    InMux I__8222 (
            .O(N__37685),
            .I(N__37679));
    LocalMux I__8221 (
            .O(N__37682),
            .I(N__37674));
    LocalMux I__8220 (
            .O(N__37679),
            .I(N__37674));
    Span4Mux_h I__8219 (
            .O(N__37674),
            .I(N__37670));
    InMux I__8218 (
            .O(N__37673),
            .I(N__37667));
    Odrv4 I__8217 (
            .O(N__37670),
            .I(\nx.n2992 ));
    LocalMux I__8216 (
            .O(N__37667),
            .I(\nx.n2992 ));
    InMux I__8215 (
            .O(N__37662),
            .I(N__37659));
    LocalMux I__8214 (
            .O(N__37659),
            .I(N__37655));
    InMux I__8213 (
            .O(N__37658),
            .I(N__37651));
    Span4Mux_h I__8212 (
            .O(N__37655),
            .I(N__37648));
    CascadeMux I__8211 (
            .O(N__37654),
            .I(N__37645));
    LocalMux I__8210 (
            .O(N__37651),
            .I(N__37642));
    Span4Mux_v I__8209 (
            .O(N__37648),
            .I(N__37639));
    InMux I__8208 (
            .O(N__37645),
            .I(N__37636));
    Span4Mux_v I__8207 (
            .O(N__37642),
            .I(N__37633));
    Odrv4 I__8206 (
            .O(N__37639),
            .I(\nx.n2794 ));
    LocalMux I__8205 (
            .O(N__37636),
            .I(\nx.n2794 ));
    Odrv4 I__8204 (
            .O(N__37633),
            .I(\nx.n2794 ));
    CascadeMux I__8203 (
            .O(N__37626),
            .I(N__37623));
    InMux I__8202 (
            .O(N__37623),
            .I(N__37620));
    LocalMux I__8201 (
            .O(N__37620),
            .I(N__37617));
    Span4Mux_h I__8200 (
            .O(N__37617),
            .I(N__37614));
    Span4Mux_h I__8199 (
            .O(N__37614),
            .I(N__37611));
    Odrv4 I__8198 (
            .O(N__37611),
            .I(\nx.n2861 ));
    CascadeMux I__8197 (
            .O(N__37608),
            .I(N__37599));
    InMux I__8196 (
            .O(N__37607),
            .I(N__37592));
    CascadeMux I__8195 (
            .O(N__37606),
            .I(N__37589));
    InMux I__8194 (
            .O(N__37605),
            .I(N__37581));
    InMux I__8193 (
            .O(N__37604),
            .I(N__37581));
    InMux I__8192 (
            .O(N__37603),
            .I(N__37581));
    CascadeMux I__8191 (
            .O(N__37602),
            .I(N__37576));
    InMux I__8190 (
            .O(N__37599),
            .I(N__37570));
    InMux I__8189 (
            .O(N__37598),
            .I(N__37570));
    InMux I__8188 (
            .O(N__37597),
            .I(N__37567));
    InMux I__8187 (
            .O(N__37596),
            .I(N__37561));
    CascadeMux I__8186 (
            .O(N__37595),
            .I(N__37557));
    LocalMux I__8185 (
            .O(N__37592),
            .I(N__37552));
    InMux I__8184 (
            .O(N__37589),
            .I(N__37547));
    InMux I__8183 (
            .O(N__37588),
            .I(N__37547));
    LocalMux I__8182 (
            .O(N__37581),
            .I(N__37544));
    InMux I__8181 (
            .O(N__37580),
            .I(N__37539));
    InMux I__8180 (
            .O(N__37579),
            .I(N__37539));
    InMux I__8179 (
            .O(N__37576),
            .I(N__37534));
    InMux I__8178 (
            .O(N__37575),
            .I(N__37534));
    LocalMux I__8177 (
            .O(N__37570),
            .I(N__37531));
    LocalMux I__8176 (
            .O(N__37567),
            .I(N__37528));
    CascadeMux I__8175 (
            .O(N__37566),
            .I(N__37525));
    CascadeMux I__8174 (
            .O(N__37565),
            .I(N__37522));
    CascadeMux I__8173 (
            .O(N__37564),
            .I(N__37518));
    LocalMux I__8172 (
            .O(N__37561),
            .I(N__37514));
    InMux I__8171 (
            .O(N__37560),
            .I(N__37506));
    InMux I__8170 (
            .O(N__37557),
            .I(N__37506));
    InMux I__8169 (
            .O(N__37556),
            .I(N__37506));
    InMux I__8168 (
            .O(N__37555),
            .I(N__37503));
    Span4Mux_v I__8167 (
            .O(N__37552),
            .I(N__37500));
    LocalMux I__8166 (
            .O(N__37547),
            .I(N__37493));
    Span4Mux_h I__8165 (
            .O(N__37544),
            .I(N__37493));
    LocalMux I__8164 (
            .O(N__37539),
            .I(N__37493));
    LocalMux I__8163 (
            .O(N__37534),
            .I(N__37486));
    Span4Mux_h I__8162 (
            .O(N__37531),
            .I(N__37486));
    Span4Mux_h I__8161 (
            .O(N__37528),
            .I(N__37486));
    InMux I__8160 (
            .O(N__37525),
            .I(N__37479));
    InMux I__8159 (
            .O(N__37522),
            .I(N__37479));
    InMux I__8158 (
            .O(N__37521),
            .I(N__37479));
    InMux I__8157 (
            .O(N__37518),
            .I(N__37474));
    InMux I__8156 (
            .O(N__37517),
            .I(N__37474));
    Span4Mux_v I__8155 (
            .O(N__37514),
            .I(N__37471));
    InMux I__8154 (
            .O(N__37513),
            .I(N__37468));
    LocalMux I__8153 (
            .O(N__37506),
            .I(\nx.n2819 ));
    LocalMux I__8152 (
            .O(N__37503),
            .I(\nx.n2819 ));
    Odrv4 I__8151 (
            .O(N__37500),
            .I(\nx.n2819 ));
    Odrv4 I__8150 (
            .O(N__37493),
            .I(\nx.n2819 ));
    Odrv4 I__8149 (
            .O(N__37486),
            .I(\nx.n2819 ));
    LocalMux I__8148 (
            .O(N__37479),
            .I(\nx.n2819 ));
    LocalMux I__8147 (
            .O(N__37474),
            .I(\nx.n2819 ));
    Odrv4 I__8146 (
            .O(N__37471),
            .I(\nx.n2819 ));
    LocalMux I__8145 (
            .O(N__37468),
            .I(\nx.n2819 ));
    InMux I__8144 (
            .O(N__37449),
            .I(N__37445));
    InMux I__8143 (
            .O(N__37448),
            .I(N__37442));
    LocalMux I__8142 (
            .O(N__37445),
            .I(\nx.n2893 ));
    LocalMux I__8141 (
            .O(N__37442),
            .I(\nx.n2893 ));
    CascadeMux I__8140 (
            .O(N__37437),
            .I(N__37433));
    InMux I__8139 (
            .O(N__37436),
            .I(N__37430));
    InMux I__8138 (
            .O(N__37433),
            .I(N__37427));
    LocalMux I__8137 (
            .O(N__37430),
            .I(N__37422));
    LocalMux I__8136 (
            .O(N__37427),
            .I(N__37422));
    Odrv4 I__8135 (
            .O(N__37422),
            .I(\nx.n2898 ));
    InMux I__8134 (
            .O(N__37419),
            .I(N__37414));
    CascadeMux I__8133 (
            .O(N__37418),
            .I(N__37411));
    InMux I__8132 (
            .O(N__37417),
            .I(N__37408));
    LocalMux I__8131 (
            .O(N__37414),
            .I(N__37405));
    InMux I__8130 (
            .O(N__37411),
            .I(N__37402));
    LocalMux I__8129 (
            .O(N__37408),
            .I(\nx.n2904 ));
    Odrv4 I__8128 (
            .O(N__37405),
            .I(\nx.n2904 ));
    LocalMux I__8127 (
            .O(N__37402),
            .I(\nx.n2904 ));
    CascadeMux I__8126 (
            .O(N__37395),
            .I(\nx.n2893_cascade_ ));
    CascadeMux I__8125 (
            .O(N__37392),
            .I(N__37389));
    InMux I__8124 (
            .O(N__37389),
            .I(N__37386));
    LocalMux I__8123 (
            .O(N__37386),
            .I(N__37383));
    Span4Mux_v I__8122 (
            .O(N__37383),
            .I(N__37378));
    InMux I__8121 (
            .O(N__37382),
            .I(N__37375));
    CascadeMux I__8120 (
            .O(N__37381),
            .I(N__37372));
    Span4Mux_h I__8119 (
            .O(N__37378),
            .I(N__37367));
    LocalMux I__8118 (
            .O(N__37375),
            .I(N__37367));
    InMux I__8117 (
            .O(N__37372),
            .I(N__37364));
    Odrv4 I__8116 (
            .O(N__37367),
            .I(\nx.n2897 ));
    LocalMux I__8115 (
            .O(N__37364),
            .I(\nx.n2897 ));
    InMux I__8114 (
            .O(N__37359),
            .I(N__37356));
    LocalMux I__8113 (
            .O(N__37356),
            .I(\nx.n41_adj_768 ));
    CascadeMux I__8112 (
            .O(N__37353),
            .I(N__37350));
    InMux I__8111 (
            .O(N__37350),
            .I(N__37346));
    InMux I__8110 (
            .O(N__37349),
            .I(N__37343));
    LocalMux I__8109 (
            .O(N__37346),
            .I(N__37340));
    LocalMux I__8108 (
            .O(N__37343),
            .I(N__37336));
    Span4Mux_h I__8107 (
            .O(N__37340),
            .I(N__37333));
    InMux I__8106 (
            .O(N__37339),
            .I(N__37330));
    Odrv12 I__8105 (
            .O(N__37336),
            .I(\nx.n2894 ));
    Odrv4 I__8104 (
            .O(N__37333),
            .I(\nx.n2894 ));
    LocalMux I__8103 (
            .O(N__37330),
            .I(\nx.n2894 ));
    CascadeMux I__8102 (
            .O(N__37323),
            .I(N__37314));
    CascadeMux I__8101 (
            .O(N__37322),
            .I(N__37308));
    InMux I__8100 (
            .O(N__37321),
            .I(N__37300));
    CascadeMux I__8099 (
            .O(N__37320),
            .I(N__37295));
    InMux I__8098 (
            .O(N__37319),
            .I(N__37288));
    InMux I__8097 (
            .O(N__37318),
            .I(N__37288));
    InMux I__8096 (
            .O(N__37317),
            .I(N__37285));
    InMux I__8095 (
            .O(N__37314),
            .I(N__37280));
    InMux I__8094 (
            .O(N__37313),
            .I(N__37280));
    InMux I__8093 (
            .O(N__37312),
            .I(N__37277));
    InMux I__8092 (
            .O(N__37311),
            .I(N__37269));
    InMux I__8091 (
            .O(N__37308),
            .I(N__37269));
    InMux I__8090 (
            .O(N__37307),
            .I(N__37269));
    InMux I__8089 (
            .O(N__37306),
            .I(N__37264));
    InMux I__8088 (
            .O(N__37305),
            .I(N__37264));
    CascadeMux I__8087 (
            .O(N__37304),
            .I(N__37259));
    CascadeMux I__8086 (
            .O(N__37303),
            .I(N__37256));
    LocalMux I__8085 (
            .O(N__37300),
            .I(N__37252));
    InMux I__8084 (
            .O(N__37299),
            .I(N__37241));
    InMux I__8083 (
            .O(N__37298),
            .I(N__37241));
    InMux I__8082 (
            .O(N__37295),
            .I(N__37241));
    InMux I__8081 (
            .O(N__37294),
            .I(N__37241));
    InMux I__8080 (
            .O(N__37293),
            .I(N__37241));
    LocalMux I__8079 (
            .O(N__37288),
            .I(N__37232));
    LocalMux I__8078 (
            .O(N__37285),
            .I(N__37232));
    LocalMux I__8077 (
            .O(N__37280),
            .I(N__37232));
    LocalMux I__8076 (
            .O(N__37277),
            .I(N__37232));
    CascadeMux I__8075 (
            .O(N__37276),
            .I(N__37228));
    LocalMux I__8074 (
            .O(N__37269),
            .I(N__37224));
    LocalMux I__8073 (
            .O(N__37264),
            .I(N__37221));
    InMux I__8072 (
            .O(N__37263),
            .I(N__37218));
    InMux I__8071 (
            .O(N__37262),
            .I(N__37215));
    InMux I__8070 (
            .O(N__37259),
            .I(N__37208));
    InMux I__8069 (
            .O(N__37256),
            .I(N__37208));
    InMux I__8068 (
            .O(N__37255),
            .I(N__37208));
    Span4Mux_h I__8067 (
            .O(N__37252),
            .I(N__37201));
    LocalMux I__8066 (
            .O(N__37241),
            .I(N__37201));
    Span4Mux_v I__8065 (
            .O(N__37232),
            .I(N__37201));
    InMux I__8064 (
            .O(N__37231),
            .I(N__37194));
    InMux I__8063 (
            .O(N__37228),
            .I(N__37194));
    InMux I__8062 (
            .O(N__37227),
            .I(N__37194));
    Span4Mux_h I__8061 (
            .O(N__37224),
            .I(N__37189));
    Span4Mux_v I__8060 (
            .O(N__37221),
            .I(N__37189));
    LocalMux I__8059 (
            .O(N__37218),
            .I(N__37186));
    LocalMux I__8058 (
            .O(N__37215),
            .I(\nx.n2918 ));
    LocalMux I__8057 (
            .O(N__37208),
            .I(\nx.n2918 ));
    Odrv4 I__8056 (
            .O(N__37201),
            .I(\nx.n2918 ));
    LocalMux I__8055 (
            .O(N__37194),
            .I(\nx.n2918 ));
    Odrv4 I__8054 (
            .O(N__37189),
            .I(\nx.n2918 ));
    Odrv4 I__8053 (
            .O(N__37186),
            .I(\nx.n2918 ));
    InMux I__8052 (
            .O(N__37173),
            .I(N__37170));
    LocalMux I__8051 (
            .O(N__37170),
            .I(\nx.n2961 ));
    InMux I__8050 (
            .O(N__37167),
            .I(N__37163));
    InMux I__8049 (
            .O(N__37166),
            .I(N__37160));
    LocalMux I__8048 (
            .O(N__37163),
            .I(N__37154));
    LocalMux I__8047 (
            .O(N__37160),
            .I(N__37154));
    InMux I__8046 (
            .O(N__37159),
            .I(N__37151));
    Odrv12 I__8045 (
            .O(N__37154),
            .I(\nx.n2993 ));
    LocalMux I__8044 (
            .O(N__37151),
            .I(\nx.n2993 ));
    InMux I__8043 (
            .O(N__37146),
            .I(N__37143));
    LocalMux I__8042 (
            .O(N__37143),
            .I(N__37140));
    Span4Mux_h I__8041 (
            .O(N__37140),
            .I(N__37137));
    Odrv4 I__8040 (
            .O(N__37137),
            .I(\nx.n40 ));
    CascadeMux I__8039 (
            .O(N__37134),
            .I(\nx.n2609_cascade_ ));
    CascadeMux I__8038 (
            .O(N__37131),
            .I(N__37128));
    InMux I__8037 (
            .O(N__37128),
            .I(N__37125));
    LocalMux I__8036 (
            .O(N__37125),
            .I(\nx.n28 ));
    CascadeMux I__8035 (
            .O(N__37122),
            .I(n6_adj_813_cascade_));
    InMux I__8034 (
            .O(N__37119),
            .I(N__37116));
    LocalMux I__8033 (
            .O(N__37116),
            .I(N__37113));
    Span4Mux_v I__8032 (
            .O(N__37113),
            .I(N__37110));
    Odrv4 I__8031 (
            .O(N__37110),
            .I(n11974));
    CascadeMux I__8030 (
            .O(N__37107),
            .I(N__37104));
    InMux I__8029 (
            .O(N__37104),
            .I(N__37099));
    CascadeMux I__8028 (
            .O(N__37103),
            .I(N__37096));
    InMux I__8027 (
            .O(N__37102),
            .I(N__37093));
    LocalMux I__8026 (
            .O(N__37099),
            .I(N__37090));
    InMux I__8025 (
            .O(N__37096),
            .I(N__37087));
    LocalMux I__8024 (
            .O(N__37093),
            .I(N__37084));
    Span4Mux_h I__8023 (
            .O(N__37090),
            .I(N__37081));
    LocalMux I__8022 (
            .O(N__37087),
            .I(N__37076));
    Span4Mux_h I__8021 (
            .O(N__37084),
            .I(N__37076));
    Span4Mux_h I__8020 (
            .O(N__37081),
            .I(N__37073));
    Span4Mux_h I__8019 (
            .O(N__37076),
            .I(N__37070));
    Odrv4 I__8018 (
            .O(N__37073),
            .I(\nx.n2890 ));
    Odrv4 I__8017 (
            .O(N__37070),
            .I(\nx.n2890 ));
    CascadeMux I__8016 (
            .O(N__37065),
            .I(N__37062));
    InMux I__8015 (
            .O(N__37062),
            .I(N__37059));
    LocalMux I__8014 (
            .O(N__37059),
            .I(N__37056));
    Span4Mux_v I__8013 (
            .O(N__37056),
            .I(N__37053));
    Span4Mux_h I__8012 (
            .O(N__37053),
            .I(N__37050));
    Odrv4 I__8011 (
            .O(N__37050),
            .I(\nx.n30_adj_759 ));
    InMux I__8010 (
            .O(N__37047),
            .I(N__37044));
    LocalMux I__8009 (
            .O(N__37044),
            .I(N__37041));
    Span4Mux_v I__8008 (
            .O(N__37041),
            .I(N__37038));
    Odrv4 I__8007 (
            .O(N__37038),
            .I(\nx.n39_adj_761 ));
    InMux I__8006 (
            .O(N__37035),
            .I(N__37032));
    LocalMux I__8005 (
            .O(N__37032),
            .I(N__37029));
    Span4Mux_v I__8004 (
            .O(N__37029),
            .I(N__37026));
    Span4Mux_h I__8003 (
            .O(N__37026),
            .I(N__37023));
    Odrv4 I__8002 (
            .O(N__37023),
            .I(\nx.n42_adj_765 ));
    CascadeMux I__8001 (
            .O(N__37020),
            .I(\nx.n45_adj_769_cascade_ ));
    InMux I__8000 (
            .O(N__37017),
            .I(N__37014));
    LocalMux I__7999 (
            .O(N__37014),
            .I(\nx.n47_adj_770 ));
    CascadeMux I__7998 (
            .O(N__37011),
            .I(N__37008));
    InMux I__7997 (
            .O(N__37008),
            .I(N__37004));
    InMux I__7996 (
            .O(N__37007),
            .I(N__37001));
    LocalMux I__7995 (
            .O(N__37004),
            .I(N__36998));
    LocalMux I__7994 (
            .O(N__37001),
            .I(\nx.n2896 ));
    Odrv4 I__7993 (
            .O(N__36998),
            .I(\nx.n2896 ));
    CascadeMux I__7992 (
            .O(N__36993),
            .I(\nx.n2918_cascade_ ));
    InMux I__7991 (
            .O(N__36990),
            .I(N__36987));
    LocalMux I__7990 (
            .O(N__36987),
            .I(\nx.n2963 ));
    InMux I__7989 (
            .O(N__36984),
            .I(N__36981));
    LocalMux I__7988 (
            .O(N__36981),
            .I(\nx.n2970 ));
    InMux I__7987 (
            .O(N__36978),
            .I(N__36974));
    InMux I__7986 (
            .O(N__36977),
            .I(N__36971));
    LocalMux I__7985 (
            .O(N__36974),
            .I(N__36966));
    LocalMux I__7984 (
            .O(N__36971),
            .I(N__36966));
    Span4Mux_h I__7983 (
            .O(N__36966),
            .I(N__36963));
    Odrv4 I__7982 (
            .O(N__36963),
            .I(\nx.n3002 ));
    InMux I__7981 (
            .O(N__36960),
            .I(N__36956));
    InMux I__7980 (
            .O(N__36959),
            .I(N__36953));
    LocalMux I__7979 (
            .O(N__36956),
            .I(N__36948));
    LocalMux I__7978 (
            .O(N__36953),
            .I(N__36948));
    Span4Mux_h I__7977 (
            .O(N__36948),
            .I(N__36944));
    InMux I__7976 (
            .O(N__36947),
            .I(N__36941));
    Odrv4 I__7975 (
            .O(N__36944),
            .I(\nx.n2995 ));
    LocalMux I__7974 (
            .O(N__36941),
            .I(\nx.n2995 ));
    CascadeMux I__7973 (
            .O(N__36936),
            .I(\nx.n3002_cascade_ ));
    InMux I__7972 (
            .O(N__36933),
            .I(N__36930));
    LocalMux I__7971 (
            .O(N__36930),
            .I(N__36927));
    Span4Mux_h I__7970 (
            .O(N__36927),
            .I(N__36924));
    Odrv4 I__7969 (
            .O(N__36924),
            .I(\nx.n42 ));
    InMux I__7968 (
            .O(N__36921),
            .I(N__36918));
    LocalMux I__7967 (
            .O(N__36918),
            .I(\nx.n2958 ));
    CascadeMux I__7966 (
            .O(N__36915),
            .I(N__36912));
    InMux I__7965 (
            .O(N__36912),
            .I(N__36908));
    CascadeMux I__7964 (
            .O(N__36911),
            .I(N__36905));
    LocalMux I__7963 (
            .O(N__36908),
            .I(N__36901));
    InMux I__7962 (
            .O(N__36905),
            .I(N__36898));
    CascadeMux I__7961 (
            .O(N__36904),
            .I(N__36895));
    Span4Mux_h I__7960 (
            .O(N__36901),
            .I(N__36892));
    LocalMux I__7959 (
            .O(N__36898),
            .I(N__36889));
    InMux I__7958 (
            .O(N__36895),
            .I(N__36886));
    Span4Mux_h I__7957 (
            .O(N__36892),
            .I(N__36883));
    Span4Mux_h I__7956 (
            .O(N__36889),
            .I(N__36878));
    LocalMux I__7955 (
            .O(N__36886),
            .I(N__36878));
    Odrv4 I__7954 (
            .O(N__36883),
            .I(\nx.n2891 ));
    Odrv4 I__7953 (
            .O(N__36878),
            .I(\nx.n2891 ));
    InMux I__7952 (
            .O(N__36873),
            .I(N__36868));
    InMux I__7951 (
            .O(N__36872),
            .I(N__36865));
    InMux I__7950 (
            .O(N__36871),
            .I(N__36862));
    LocalMux I__7949 (
            .O(N__36868),
            .I(N__36857));
    LocalMux I__7948 (
            .O(N__36865),
            .I(N__36857));
    LocalMux I__7947 (
            .O(N__36862),
            .I(N__36854));
    Odrv12 I__7946 (
            .O(N__36857),
            .I(\nx.n2990 ));
    Odrv4 I__7945 (
            .O(N__36854),
            .I(\nx.n2990 ));
    InMux I__7944 (
            .O(N__36849),
            .I(N__36846));
    LocalMux I__7943 (
            .O(N__36846),
            .I(N__36842));
    CascadeMux I__7942 (
            .O(N__36845),
            .I(N__36838));
    Span12Mux_h I__7941 (
            .O(N__36842),
            .I(N__36835));
    InMux I__7940 (
            .O(N__36841),
            .I(N__36832));
    InMux I__7939 (
            .O(N__36838),
            .I(N__36829));
    Odrv12 I__7938 (
            .O(N__36835),
            .I(\nx.n2804 ));
    LocalMux I__7937 (
            .O(N__36832),
            .I(\nx.n2804 ));
    LocalMux I__7936 (
            .O(N__36829),
            .I(\nx.n2804 ));
    CascadeMux I__7935 (
            .O(N__36822),
            .I(N__36819));
    InMux I__7934 (
            .O(N__36819),
            .I(N__36816));
    LocalMux I__7933 (
            .O(N__36816),
            .I(N__36813));
    Span4Mux_h I__7932 (
            .O(N__36813),
            .I(N__36810));
    Span4Mux_h I__7931 (
            .O(N__36810),
            .I(N__36807));
    Odrv4 I__7930 (
            .O(N__36807),
            .I(\nx.n2871 ));
    CascadeMux I__7929 (
            .O(N__36804),
            .I(N__36799));
    InMux I__7928 (
            .O(N__36803),
            .I(N__36796));
    CascadeMux I__7927 (
            .O(N__36802),
            .I(N__36793));
    InMux I__7926 (
            .O(N__36799),
            .I(N__36790));
    LocalMux I__7925 (
            .O(N__36796),
            .I(N__36787));
    InMux I__7924 (
            .O(N__36793),
            .I(N__36784));
    LocalMux I__7923 (
            .O(N__36790),
            .I(\nx.n2903 ));
    Odrv4 I__7922 (
            .O(N__36787),
            .I(\nx.n2903 ));
    LocalMux I__7921 (
            .O(N__36784),
            .I(\nx.n2903 ));
    IoInMux I__7920 (
            .O(N__36777),
            .I(N__36774));
    LocalMux I__7919 (
            .O(N__36774),
            .I(N__36771));
    Span12Mux_s4_v I__7918 (
            .O(N__36771),
            .I(N__36768));
    Span12Mux_h I__7917 (
            .O(N__36768),
            .I(N__36764));
    InMux I__7916 (
            .O(N__36767),
            .I(N__36761));
    Odrv12 I__7915 (
            .O(N__36764),
            .I(pin_oe_9));
    LocalMux I__7914 (
            .O(N__36761),
            .I(pin_oe_9));
    IoInMux I__7913 (
            .O(N__36756),
            .I(N__36753));
    LocalMux I__7912 (
            .O(N__36753),
            .I(N__36750));
    Span12Mux_s6_v I__7911 (
            .O(N__36750),
            .I(N__36747));
    Span12Mux_h I__7910 (
            .O(N__36747),
            .I(N__36743));
    InMux I__7909 (
            .O(N__36746),
            .I(N__36740));
    Odrv12 I__7908 (
            .O(N__36743),
            .I(pin_oe_10));
    LocalMux I__7907 (
            .O(N__36740),
            .I(pin_oe_10));
    InMux I__7906 (
            .O(N__36735),
            .I(N__36732));
    LocalMux I__7905 (
            .O(N__36732),
            .I(n11960));
    InMux I__7904 (
            .O(N__36729),
            .I(N__36726));
    LocalMux I__7903 (
            .O(N__36726),
            .I(n2618));
    IoInMux I__7902 (
            .O(N__36723),
            .I(N__36720));
    LocalMux I__7901 (
            .O(N__36720),
            .I(N__36717));
    Span12Mux_s2_h I__7900 (
            .O(N__36717),
            .I(N__36714));
    Span12Mux_h I__7899 (
            .O(N__36714),
            .I(N__36710));
    InMux I__7898 (
            .O(N__36713),
            .I(N__36707));
    Odrv12 I__7897 (
            .O(N__36710),
            .I(pin_oe_3));
    LocalMux I__7896 (
            .O(N__36707),
            .I(pin_oe_3));
    CascadeMux I__7895 (
            .O(N__36702),
            .I(n8_adj_825_cascade_));
    IoInMux I__7894 (
            .O(N__36699),
            .I(N__36696));
    LocalMux I__7893 (
            .O(N__36696),
            .I(N__36693));
    Span12Mux_s7_v I__7892 (
            .O(N__36693),
            .I(N__36690));
    Span12Mux_h I__7891 (
            .O(N__36690),
            .I(N__36685));
    InMux I__7890 (
            .O(N__36689),
            .I(N__36682));
    InMux I__7889 (
            .O(N__36688),
            .I(N__36679));
    Odrv12 I__7888 (
            .O(N__36685),
            .I(pin_out_9));
    LocalMux I__7887 (
            .O(N__36682),
            .I(pin_out_9));
    LocalMux I__7886 (
            .O(N__36679),
            .I(pin_out_9));
    InMux I__7885 (
            .O(N__36672),
            .I(N__36668));
    CascadeMux I__7884 (
            .O(N__36671),
            .I(N__36665));
    LocalMux I__7883 (
            .O(N__36668),
            .I(N__36661));
    InMux I__7882 (
            .O(N__36665),
            .I(N__36658));
    InMux I__7881 (
            .O(N__36664),
            .I(N__36655));
    Odrv4 I__7880 (
            .O(N__36661),
            .I(\nx.n2297 ));
    LocalMux I__7879 (
            .O(N__36658),
            .I(\nx.n2297 ));
    LocalMux I__7878 (
            .O(N__36655),
            .I(\nx.n2297 ));
    CascadeMux I__7877 (
            .O(N__36648),
            .I(N__36645));
    InMux I__7876 (
            .O(N__36645),
            .I(N__36642));
    LocalMux I__7875 (
            .O(N__36642),
            .I(\nx.n2364 ));
    InMux I__7874 (
            .O(N__36639),
            .I(N__36635));
    CascadeMux I__7873 (
            .O(N__36638),
            .I(N__36632));
    LocalMux I__7872 (
            .O(N__36635),
            .I(N__36628));
    InMux I__7871 (
            .O(N__36632),
            .I(N__36625));
    InMux I__7870 (
            .O(N__36631),
            .I(N__36622));
    Odrv4 I__7869 (
            .O(N__36628),
            .I(\nx.n2298 ));
    LocalMux I__7868 (
            .O(N__36625),
            .I(\nx.n2298 ));
    LocalMux I__7867 (
            .O(N__36622),
            .I(\nx.n2298 ));
    CascadeMux I__7866 (
            .O(N__36615),
            .I(N__36612));
    InMux I__7865 (
            .O(N__36612),
            .I(N__36609));
    LocalMux I__7864 (
            .O(N__36609),
            .I(\nx.n2365 ));
    InMux I__7863 (
            .O(N__36606),
            .I(N__36603));
    LocalMux I__7862 (
            .O(N__36603),
            .I(N__36600));
    Span4Mux_h I__7861 (
            .O(N__36600),
            .I(N__36597));
    Odrv4 I__7860 (
            .O(N__36597),
            .I(\nx.n2168 ));
    CascadeMux I__7859 (
            .O(N__36594),
            .I(N__36590));
    CascadeMux I__7858 (
            .O(N__36593),
            .I(N__36587));
    InMux I__7857 (
            .O(N__36590),
            .I(N__36584));
    InMux I__7856 (
            .O(N__36587),
            .I(N__36581));
    LocalMux I__7855 (
            .O(N__36584),
            .I(N__36577));
    LocalMux I__7854 (
            .O(N__36581),
            .I(N__36574));
    InMux I__7853 (
            .O(N__36580),
            .I(N__36571));
    Odrv12 I__7852 (
            .O(N__36577),
            .I(\nx.n2101 ));
    Odrv4 I__7851 (
            .O(N__36574),
            .I(\nx.n2101 ));
    LocalMux I__7850 (
            .O(N__36571),
            .I(\nx.n2101 ));
    CascadeMux I__7849 (
            .O(N__36564),
            .I(N__36554));
    CascadeMux I__7848 (
            .O(N__36563),
            .I(N__36549));
    InMux I__7847 (
            .O(N__36562),
            .I(N__36545));
    CascadeMux I__7846 (
            .O(N__36561),
            .I(N__36542));
    CascadeMux I__7845 (
            .O(N__36560),
            .I(N__36539));
    CascadeMux I__7844 (
            .O(N__36559),
            .I(N__36535));
    CascadeMux I__7843 (
            .O(N__36558),
            .I(N__36529));
    CascadeMux I__7842 (
            .O(N__36557),
            .I(N__36526));
    InMux I__7841 (
            .O(N__36554),
            .I(N__36519));
    InMux I__7840 (
            .O(N__36553),
            .I(N__36519));
    InMux I__7839 (
            .O(N__36552),
            .I(N__36512));
    InMux I__7838 (
            .O(N__36549),
            .I(N__36512));
    InMux I__7837 (
            .O(N__36548),
            .I(N__36512));
    LocalMux I__7836 (
            .O(N__36545),
            .I(N__36509));
    InMux I__7835 (
            .O(N__36542),
            .I(N__36506));
    InMux I__7834 (
            .O(N__36539),
            .I(N__36501));
    InMux I__7833 (
            .O(N__36538),
            .I(N__36501));
    InMux I__7832 (
            .O(N__36535),
            .I(N__36496));
    InMux I__7831 (
            .O(N__36534),
            .I(N__36496));
    InMux I__7830 (
            .O(N__36533),
            .I(N__36491));
    InMux I__7829 (
            .O(N__36532),
            .I(N__36491));
    InMux I__7828 (
            .O(N__36529),
            .I(N__36482));
    InMux I__7827 (
            .O(N__36526),
            .I(N__36482));
    InMux I__7826 (
            .O(N__36525),
            .I(N__36482));
    InMux I__7825 (
            .O(N__36524),
            .I(N__36482));
    LocalMux I__7824 (
            .O(N__36519),
            .I(N__36475));
    LocalMux I__7823 (
            .O(N__36512),
            .I(N__36475));
    Span4Mux_v I__7822 (
            .O(N__36509),
            .I(N__36475));
    LocalMux I__7821 (
            .O(N__36506),
            .I(N__36472));
    LocalMux I__7820 (
            .O(N__36501),
            .I(\nx.n2126 ));
    LocalMux I__7819 (
            .O(N__36496),
            .I(\nx.n2126 ));
    LocalMux I__7818 (
            .O(N__36491),
            .I(\nx.n2126 ));
    LocalMux I__7817 (
            .O(N__36482),
            .I(\nx.n2126 ));
    Odrv4 I__7816 (
            .O(N__36475),
            .I(\nx.n2126 ));
    Odrv12 I__7815 (
            .O(N__36472),
            .I(\nx.n2126 ));
    CascadeMux I__7814 (
            .O(N__36459),
            .I(N__36456));
    InMux I__7813 (
            .O(N__36456),
            .I(N__36451));
    InMux I__7812 (
            .O(N__36455),
            .I(N__36448));
    InMux I__7811 (
            .O(N__36454),
            .I(N__36445));
    LocalMux I__7810 (
            .O(N__36451),
            .I(N__36442));
    LocalMux I__7809 (
            .O(N__36448),
            .I(N__36439));
    LocalMux I__7808 (
            .O(N__36445),
            .I(N__36436));
    Span4Mux_h I__7807 (
            .O(N__36442),
            .I(N__36433));
    Span4Mux_h I__7806 (
            .O(N__36439),
            .I(N__36430));
    Odrv4 I__7805 (
            .O(N__36436),
            .I(\nx.n2200 ));
    Odrv4 I__7804 (
            .O(N__36433),
            .I(\nx.n2200 ));
    Odrv4 I__7803 (
            .O(N__36430),
            .I(\nx.n2200 ));
    InMux I__7802 (
            .O(N__36423),
            .I(N__36419));
    CascadeMux I__7801 (
            .O(N__36422),
            .I(N__36416));
    LocalMux I__7800 (
            .O(N__36419),
            .I(N__36412));
    InMux I__7799 (
            .O(N__36416),
            .I(N__36409));
    InMux I__7798 (
            .O(N__36415),
            .I(N__36406));
    Span4Mux_h I__7797 (
            .O(N__36412),
            .I(N__36401));
    LocalMux I__7796 (
            .O(N__36409),
            .I(N__36401));
    LocalMux I__7795 (
            .O(N__36406),
            .I(\nx.n2301 ));
    Odrv4 I__7794 (
            .O(N__36401),
            .I(\nx.n2301 ));
    CascadeMux I__7793 (
            .O(N__36396),
            .I(N__36393));
    InMux I__7792 (
            .O(N__36393),
            .I(N__36390));
    LocalMux I__7791 (
            .O(N__36390),
            .I(\nx.n2368 ));
    CascadeMux I__7790 (
            .O(N__36387),
            .I(n7602_cascade_));
    CascadeMux I__7789 (
            .O(N__36384),
            .I(n7730_cascade_));
    InMux I__7788 (
            .O(N__36381),
            .I(\nx.n10931 ));
    InMux I__7787 (
            .O(N__36378),
            .I(\nx.n10932 ));
    InMux I__7786 (
            .O(N__36375),
            .I(bfn_14_26_0_));
    InMux I__7785 (
            .O(N__36372),
            .I(\nx.n10934 ));
    InMux I__7784 (
            .O(N__36369),
            .I(\nx.n10935 ));
    InMux I__7783 (
            .O(N__36366),
            .I(\nx.n10936 ));
    CascadeMux I__7782 (
            .O(N__36363),
            .I(N__36360));
    InMux I__7781 (
            .O(N__36360),
            .I(N__36356));
    InMux I__7780 (
            .O(N__36359),
            .I(N__36353));
    LocalMux I__7779 (
            .O(N__36356),
            .I(N__36350));
    LocalMux I__7778 (
            .O(N__36353),
            .I(N__36347));
    Odrv4 I__7777 (
            .O(N__36350),
            .I(\nx.n2390 ));
    Odrv4 I__7776 (
            .O(N__36347),
            .I(\nx.n2390 ));
    InMux I__7775 (
            .O(N__36342),
            .I(\nx.n10937 ));
    IoInMux I__7774 (
            .O(N__36339),
            .I(N__36336));
    LocalMux I__7773 (
            .O(N__36336),
            .I(N__36333));
    Span12Mux_s6_v I__7772 (
            .O(N__36333),
            .I(N__36330));
    Span12Mux_h I__7771 (
            .O(N__36330),
            .I(N__36326));
    InMux I__7770 (
            .O(N__36329),
            .I(N__36323));
    Odrv12 I__7769 (
            .O(N__36326),
            .I(pin_oe_18));
    LocalMux I__7768 (
            .O(N__36323),
            .I(pin_oe_18));
    CascadeMux I__7767 (
            .O(N__36318),
            .I(N__36314));
    InMux I__7766 (
            .O(N__36317),
            .I(N__36311));
    InMux I__7765 (
            .O(N__36314),
            .I(N__36308));
    LocalMux I__7764 (
            .O(N__36311),
            .I(N__36302));
    LocalMux I__7763 (
            .O(N__36308),
            .I(N__36302));
    InMux I__7762 (
            .O(N__36307),
            .I(N__36299));
    Odrv4 I__7761 (
            .O(N__36302),
            .I(\nx.n2295 ));
    LocalMux I__7760 (
            .O(N__36299),
            .I(\nx.n2295 ));
    CascadeMux I__7759 (
            .O(N__36294),
            .I(N__36291));
    InMux I__7758 (
            .O(N__36291),
            .I(N__36288));
    LocalMux I__7757 (
            .O(N__36288),
            .I(\nx.n2362 ));
    InMux I__7756 (
            .O(N__36285),
            .I(\nx.n10922 ));
    CascadeMux I__7755 (
            .O(N__36282),
            .I(N__36278));
    CascadeMux I__7754 (
            .O(N__36281),
            .I(N__36275));
    InMux I__7753 (
            .O(N__36278),
            .I(N__36271));
    InMux I__7752 (
            .O(N__36275),
            .I(N__36268));
    InMux I__7751 (
            .O(N__36274),
            .I(N__36265));
    LocalMux I__7750 (
            .O(N__36271),
            .I(\nx.n2404 ));
    LocalMux I__7749 (
            .O(N__36268),
            .I(\nx.n2404 ));
    LocalMux I__7748 (
            .O(N__36265),
            .I(\nx.n2404 ));
    InMux I__7747 (
            .O(N__36258),
            .I(N__36255));
    LocalMux I__7746 (
            .O(N__36255),
            .I(\nx.n2471 ));
    InMux I__7745 (
            .O(N__36252),
            .I(\nx.n10923 ));
    CascadeMux I__7744 (
            .O(N__36249),
            .I(N__36246));
    InMux I__7743 (
            .O(N__36246),
            .I(N__36242));
    CascadeMux I__7742 (
            .O(N__36245),
            .I(N__36239));
    LocalMux I__7741 (
            .O(N__36242),
            .I(N__36235));
    InMux I__7740 (
            .O(N__36239),
            .I(N__36232));
    InMux I__7739 (
            .O(N__36238),
            .I(N__36229));
    Odrv4 I__7738 (
            .O(N__36235),
            .I(\nx.n2403 ));
    LocalMux I__7737 (
            .O(N__36232),
            .I(\nx.n2403 ));
    LocalMux I__7736 (
            .O(N__36229),
            .I(\nx.n2403 ));
    InMux I__7735 (
            .O(N__36222),
            .I(N__36219));
    LocalMux I__7734 (
            .O(N__36219),
            .I(\nx.n2470 ));
    InMux I__7733 (
            .O(N__36216),
            .I(\nx.n10924 ));
    CascadeMux I__7732 (
            .O(N__36213),
            .I(N__36209));
    InMux I__7731 (
            .O(N__36212),
            .I(N__36206));
    InMux I__7730 (
            .O(N__36209),
            .I(N__36203));
    LocalMux I__7729 (
            .O(N__36206),
            .I(N__36199));
    LocalMux I__7728 (
            .O(N__36203),
            .I(N__36196));
    InMux I__7727 (
            .O(N__36202),
            .I(N__36193));
    Odrv4 I__7726 (
            .O(N__36199),
            .I(\nx.n2402 ));
    Odrv4 I__7725 (
            .O(N__36196),
            .I(\nx.n2402 ));
    LocalMux I__7724 (
            .O(N__36193),
            .I(\nx.n2402 ));
    InMux I__7723 (
            .O(N__36186),
            .I(N__36183));
    LocalMux I__7722 (
            .O(N__36183),
            .I(N__36180));
    Odrv4 I__7721 (
            .O(N__36180),
            .I(\nx.n2469 ));
    InMux I__7720 (
            .O(N__36177),
            .I(bfn_14_25_0_));
    CascadeMux I__7719 (
            .O(N__36174),
            .I(N__36171));
    InMux I__7718 (
            .O(N__36171),
            .I(N__36167));
    CascadeMux I__7717 (
            .O(N__36170),
            .I(N__36164));
    LocalMux I__7716 (
            .O(N__36167),
            .I(N__36161));
    InMux I__7715 (
            .O(N__36164),
            .I(N__36158));
    Span4Mux_h I__7714 (
            .O(N__36161),
            .I(N__36155));
    LocalMux I__7713 (
            .O(N__36158),
            .I(N__36152));
    Odrv4 I__7712 (
            .O(N__36155),
            .I(\nx.n2401 ));
    Odrv4 I__7711 (
            .O(N__36152),
            .I(\nx.n2401 ));
    InMux I__7710 (
            .O(N__36147),
            .I(N__36144));
    LocalMux I__7709 (
            .O(N__36144),
            .I(N__36141));
    Odrv4 I__7708 (
            .O(N__36141),
            .I(\nx.n2468 ));
    InMux I__7707 (
            .O(N__36138),
            .I(\nx.n10926 ));
    InMux I__7706 (
            .O(N__36135),
            .I(\nx.n10927 ));
    CascadeMux I__7705 (
            .O(N__36132),
            .I(N__36128));
    CascadeMux I__7704 (
            .O(N__36131),
            .I(N__36124));
    InMux I__7703 (
            .O(N__36128),
            .I(N__36121));
    CascadeMux I__7702 (
            .O(N__36127),
            .I(N__36118));
    InMux I__7701 (
            .O(N__36124),
            .I(N__36115));
    LocalMux I__7700 (
            .O(N__36121),
            .I(N__36112));
    InMux I__7699 (
            .O(N__36118),
            .I(N__36109));
    LocalMux I__7698 (
            .O(N__36115),
            .I(N__36106));
    Odrv4 I__7697 (
            .O(N__36112),
            .I(\nx.n2399 ));
    LocalMux I__7696 (
            .O(N__36109),
            .I(\nx.n2399 ));
    Odrv4 I__7695 (
            .O(N__36106),
            .I(\nx.n2399 ));
    InMux I__7694 (
            .O(N__36099),
            .I(N__36096));
    LocalMux I__7693 (
            .O(N__36096),
            .I(N__36093));
    Span4Mux_h I__7692 (
            .O(N__36093),
            .I(N__36090));
    Odrv4 I__7691 (
            .O(N__36090),
            .I(\nx.n2466 ));
    InMux I__7690 (
            .O(N__36087),
            .I(\nx.n10928 ));
    InMux I__7689 (
            .O(N__36084),
            .I(\nx.n10929 ));
    InMux I__7688 (
            .O(N__36081),
            .I(\nx.n10930 ));
    CascadeMux I__7687 (
            .O(N__36078),
            .I(\nx.n2423_cascade_ ));
    InMux I__7686 (
            .O(N__36075),
            .I(N__36072));
    LocalMux I__7685 (
            .O(N__36072),
            .I(N__36068));
    InMux I__7684 (
            .O(N__36071),
            .I(N__36065));
    Odrv4 I__7683 (
            .O(N__36068),
            .I(\nx.n2374 ));
    LocalMux I__7682 (
            .O(N__36065),
            .I(\nx.n2374 ));
    InMux I__7681 (
            .O(N__36060),
            .I(N__36054));
    InMux I__7680 (
            .O(N__36059),
            .I(N__36049));
    InMux I__7679 (
            .O(N__36058),
            .I(N__36049));
    InMux I__7678 (
            .O(N__36057),
            .I(N__36046));
    LocalMux I__7677 (
            .O(N__36054),
            .I(N__36042));
    LocalMux I__7676 (
            .O(N__36049),
            .I(N__36039));
    LocalMux I__7675 (
            .O(N__36046),
            .I(N__36036));
    InMux I__7674 (
            .O(N__36045),
            .I(N__36033));
    Span4Mux_v I__7673 (
            .O(N__36042),
            .I(N__36030));
    Span12Mux_h I__7672 (
            .O(N__36039),
            .I(N__36027));
    Span12Mux_h I__7671 (
            .O(N__36036),
            .I(N__36024));
    LocalMux I__7670 (
            .O(N__36033),
            .I(\nx.bit_ctr_11 ));
    Odrv4 I__7669 (
            .O(N__36030),
            .I(\nx.bit_ctr_11 ));
    Odrv12 I__7668 (
            .O(N__36027),
            .I(\nx.bit_ctr_11 ));
    Odrv12 I__7667 (
            .O(N__36024),
            .I(\nx.bit_ctr_11 ));
    InMux I__7666 (
            .O(N__36015),
            .I(N__36012));
    LocalMux I__7665 (
            .O(N__36012),
            .I(\nx.n2477 ));
    InMux I__7664 (
            .O(N__36009),
            .I(bfn_14_24_0_));
    InMux I__7663 (
            .O(N__36006),
            .I(\nx.n10918 ));
    CascadeMux I__7662 (
            .O(N__36003),
            .I(N__35999));
    CascadeMux I__7661 (
            .O(N__36002),
            .I(N__35996));
    InMux I__7660 (
            .O(N__35999),
            .I(N__35992));
    InMux I__7659 (
            .O(N__35996),
            .I(N__35989));
    InMux I__7658 (
            .O(N__35995),
            .I(N__35986));
    LocalMux I__7657 (
            .O(N__35992),
            .I(\nx.n2408 ));
    LocalMux I__7656 (
            .O(N__35989),
            .I(\nx.n2408 ));
    LocalMux I__7655 (
            .O(N__35986),
            .I(\nx.n2408 ));
    InMux I__7654 (
            .O(N__35979),
            .I(N__35976));
    LocalMux I__7653 (
            .O(N__35976),
            .I(\nx.n2475 ));
    InMux I__7652 (
            .O(N__35973),
            .I(\nx.n10919 ));
    CascadeMux I__7651 (
            .O(N__35970),
            .I(N__35965));
    CascadeMux I__7650 (
            .O(N__35969),
            .I(N__35962));
    InMux I__7649 (
            .O(N__35968),
            .I(N__35957));
    InMux I__7648 (
            .O(N__35965),
            .I(N__35957));
    InMux I__7647 (
            .O(N__35962),
            .I(N__35954));
    LocalMux I__7646 (
            .O(N__35957),
            .I(\nx.n2407 ));
    LocalMux I__7645 (
            .O(N__35954),
            .I(\nx.n2407 ));
    InMux I__7644 (
            .O(N__35949),
            .I(N__35946));
    LocalMux I__7643 (
            .O(N__35946),
            .I(\nx.n2474 ));
    InMux I__7642 (
            .O(N__35943),
            .I(\nx.n10920 ));
    CascadeMux I__7641 (
            .O(N__35940),
            .I(N__35937));
    InMux I__7640 (
            .O(N__35937),
            .I(N__35933));
    InMux I__7639 (
            .O(N__35936),
            .I(N__35930));
    LocalMux I__7638 (
            .O(N__35933),
            .I(\nx.n2406 ));
    LocalMux I__7637 (
            .O(N__35930),
            .I(\nx.n2406 ));
    CascadeMux I__7636 (
            .O(N__35925),
            .I(N__35922));
    InMux I__7635 (
            .O(N__35922),
            .I(N__35919));
    LocalMux I__7634 (
            .O(N__35919),
            .I(\nx.n2473 ));
    InMux I__7633 (
            .O(N__35916),
            .I(\nx.n10921 ));
    InMux I__7632 (
            .O(N__35913),
            .I(N__35909));
    CascadeMux I__7631 (
            .O(N__35912),
            .I(N__35906));
    LocalMux I__7630 (
            .O(N__35909),
            .I(N__35902));
    InMux I__7629 (
            .O(N__35906),
            .I(N__35899));
    InMux I__7628 (
            .O(N__35905),
            .I(N__35896));
    Odrv4 I__7627 (
            .O(N__35902),
            .I(\nx.n2405 ));
    LocalMux I__7626 (
            .O(N__35899),
            .I(\nx.n2405 ));
    LocalMux I__7625 (
            .O(N__35896),
            .I(\nx.n2405 ));
    InMux I__7624 (
            .O(N__35889),
            .I(N__35886));
    LocalMux I__7623 (
            .O(N__35886),
            .I(\nx.n2472 ));
    InMux I__7622 (
            .O(N__35883),
            .I(N__35880));
    LocalMux I__7621 (
            .O(N__35880),
            .I(N__35877));
    Odrv12 I__7620 (
            .O(N__35877),
            .I(\nx.n2953 ));
    InMux I__7619 (
            .O(N__35874),
            .I(bfn_14_22_0_));
    CascadeMux I__7618 (
            .O(N__35871),
            .I(N__35868));
    InMux I__7617 (
            .O(N__35868),
            .I(N__35865));
    LocalMux I__7616 (
            .O(N__35865),
            .I(N__35862));
    Span4Mux_v I__7615 (
            .O(N__35862),
            .I(N__35858));
    InMux I__7614 (
            .O(N__35861),
            .I(N__35855));
    Span4Mux_h I__7613 (
            .O(N__35858),
            .I(N__35850));
    LocalMux I__7612 (
            .O(N__35855),
            .I(N__35850));
    Odrv4 I__7611 (
            .O(N__35850),
            .I(\nx.n2885 ));
    InMux I__7610 (
            .O(N__35847),
            .I(\nx.n11052 ));
    InMux I__7609 (
            .O(N__35844),
            .I(N__35840));
    InMux I__7608 (
            .O(N__35843),
            .I(N__35837));
    LocalMux I__7607 (
            .O(N__35840),
            .I(N__35831));
    LocalMux I__7606 (
            .O(N__35837),
            .I(N__35831));
    InMux I__7605 (
            .O(N__35836),
            .I(N__35828));
    Span4Mux_v I__7604 (
            .O(N__35831),
            .I(N__35823));
    LocalMux I__7603 (
            .O(N__35828),
            .I(N__35823));
    Span4Mux_h I__7602 (
            .O(N__35823),
            .I(N__35820));
    Odrv4 I__7601 (
            .O(N__35820),
            .I(\nx.n2984 ));
    InMux I__7600 (
            .O(N__35817),
            .I(N__35814));
    LocalMux I__7599 (
            .O(N__35814),
            .I(\nx.n27_adj_757 ));
    InMux I__7598 (
            .O(N__35811),
            .I(N__35808));
    LocalMux I__7597 (
            .O(N__35808),
            .I(\nx.n36_adj_756 ));
    InMux I__7596 (
            .O(N__35805),
            .I(N__35800));
    InMux I__7595 (
            .O(N__35804),
            .I(N__35797));
    CascadeMux I__7594 (
            .O(N__35803),
            .I(N__35794));
    LocalMux I__7593 (
            .O(N__35800),
            .I(N__35791));
    LocalMux I__7592 (
            .O(N__35797),
            .I(N__35788));
    InMux I__7591 (
            .O(N__35794),
            .I(N__35785));
    Span4Mux_v I__7590 (
            .O(N__35791),
            .I(N__35778));
    Span4Mux_v I__7589 (
            .O(N__35788),
            .I(N__35778));
    LocalMux I__7588 (
            .O(N__35785),
            .I(N__35778));
    Odrv4 I__7587 (
            .O(N__35778),
            .I(\nx.n2708 ));
    CascadeMux I__7586 (
            .O(N__35775),
            .I(N__35772));
    InMux I__7585 (
            .O(N__35772),
            .I(N__35768));
    InMux I__7584 (
            .O(N__35771),
            .I(N__35765));
    LocalMux I__7583 (
            .O(N__35768),
            .I(N__35761));
    LocalMux I__7582 (
            .O(N__35765),
            .I(N__35758));
    InMux I__7581 (
            .O(N__35764),
            .I(N__35755));
    Span4Mux_h I__7580 (
            .O(N__35761),
            .I(N__35752));
    Odrv12 I__7579 (
            .O(N__35758),
            .I(\nx.n2703 ));
    LocalMux I__7578 (
            .O(N__35755),
            .I(\nx.n2703 ));
    Odrv4 I__7577 (
            .O(N__35752),
            .I(\nx.n2703 ));
    InMux I__7576 (
            .O(N__35745),
            .I(N__35742));
    LocalMux I__7575 (
            .O(N__35742),
            .I(N__35739));
    Odrv12 I__7574 (
            .O(N__35739),
            .I(\nx.n39_adj_689 ));
    CascadeMux I__7573 (
            .O(N__35736),
            .I(\nx.n25_adj_702_cascade_ ));
    InMux I__7572 (
            .O(N__35733),
            .I(N__35730));
    LocalMux I__7571 (
            .O(N__35730),
            .I(N__35727));
    Span4Mux_h I__7570 (
            .O(N__35727),
            .I(N__35724));
    Odrv4 I__7569 (
            .O(N__35724),
            .I(\nx.n34_adj_701 ));
    InMux I__7568 (
            .O(N__35721),
            .I(N__35718));
    LocalMux I__7567 (
            .O(N__35718),
            .I(N__35715));
    Odrv4 I__7566 (
            .O(N__35715),
            .I(\nx.n35_adj_708 ));
    InMux I__7565 (
            .O(N__35712),
            .I(N__35709));
    LocalMux I__7564 (
            .O(N__35709),
            .I(\nx.n32_adj_703 ));
    CascadeMux I__7563 (
            .O(N__35706),
            .I(\nx.n37_adj_709_cascade_ ));
    InMux I__7562 (
            .O(N__35703),
            .I(N__35700));
    LocalMux I__7561 (
            .O(N__35700),
            .I(N__35697));
    Span4Mux_v I__7560 (
            .O(N__35697),
            .I(N__35694));
    Odrv4 I__7559 (
            .O(N__35694),
            .I(\nx.n31_adj_707 ));
    InMux I__7558 (
            .O(N__35691),
            .I(bfn_14_21_0_));
    InMux I__7557 (
            .O(N__35688),
            .I(\nx.n11044 ));
    InMux I__7556 (
            .O(N__35685),
            .I(N__35682));
    LocalMux I__7555 (
            .O(N__35682),
            .I(\nx.n2959 ));
    InMux I__7554 (
            .O(N__35679),
            .I(\nx.n11045 ));
    InMux I__7553 (
            .O(N__35676),
            .I(\nx.n11046 ));
    InMux I__7552 (
            .O(N__35673),
            .I(N__35670));
    LocalMux I__7551 (
            .O(N__35670),
            .I(N__35667));
    Span4Mux_h I__7550 (
            .O(N__35667),
            .I(N__35664));
    Odrv4 I__7549 (
            .O(N__35664),
            .I(\nx.n2957 ));
    InMux I__7548 (
            .O(N__35661),
            .I(\nx.n11047 ));
    CascadeMux I__7547 (
            .O(N__35658),
            .I(N__35654));
    InMux I__7546 (
            .O(N__35657),
            .I(N__35651));
    InMux I__7545 (
            .O(N__35654),
            .I(N__35648));
    LocalMux I__7544 (
            .O(N__35651),
            .I(N__35643));
    LocalMux I__7543 (
            .O(N__35648),
            .I(N__35643));
    Span4Mux_h I__7542 (
            .O(N__35643),
            .I(N__35640));
    Odrv4 I__7541 (
            .O(N__35640),
            .I(\nx.n2889 ));
    CascadeMux I__7540 (
            .O(N__35637),
            .I(N__35634));
    InMux I__7539 (
            .O(N__35634),
            .I(N__35631));
    LocalMux I__7538 (
            .O(N__35631),
            .I(N__35628));
    Odrv4 I__7537 (
            .O(N__35628),
            .I(\nx.n2956 ));
    InMux I__7536 (
            .O(N__35625),
            .I(\nx.n11048 ));
    CascadeMux I__7535 (
            .O(N__35622),
            .I(N__35619));
    InMux I__7534 (
            .O(N__35619),
            .I(N__35616));
    LocalMux I__7533 (
            .O(N__35616),
            .I(N__35613));
    Span4Mux_v I__7532 (
            .O(N__35613),
            .I(N__35608));
    InMux I__7531 (
            .O(N__35612),
            .I(N__35605));
    InMux I__7530 (
            .O(N__35611),
            .I(N__35602));
    Span4Mux_h I__7529 (
            .O(N__35608),
            .I(N__35599));
    LocalMux I__7528 (
            .O(N__35605),
            .I(N__35596));
    LocalMux I__7527 (
            .O(N__35602),
            .I(\nx.n2888 ));
    Odrv4 I__7526 (
            .O(N__35599),
            .I(\nx.n2888 ));
    Odrv4 I__7525 (
            .O(N__35596),
            .I(\nx.n2888 ));
    CascadeMux I__7524 (
            .O(N__35589),
            .I(N__35586));
    InMux I__7523 (
            .O(N__35586),
            .I(N__35583));
    LocalMux I__7522 (
            .O(N__35583),
            .I(N__35580));
    Span4Mux_h I__7521 (
            .O(N__35580),
            .I(N__35577));
    Odrv4 I__7520 (
            .O(N__35577),
            .I(\nx.n2955 ));
    InMux I__7519 (
            .O(N__35574),
            .I(\nx.n11049 ));
    CascadeMux I__7518 (
            .O(N__35571),
            .I(N__35567));
    InMux I__7517 (
            .O(N__35570),
            .I(N__35564));
    InMux I__7516 (
            .O(N__35567),
            .I(N__35561));
    LocalMux I__7515 (
            .O(N__35564),
            .I(N__35555));
    LocalMux I__7514 (
            .O(N__35561),
            .I(N__35555));
    InMux I__7513 (
            .O(N__35560),
            .I(N__35552));
    Odrv4 I__7512 (
            .O(N__35555),
            .I(\nx.n2887 ));
    LocalMux I__7511 (
            .O(N__35552),
            .I(\nx.n2887 ));
    CascadeMux I__7510 (
            .O(N__35547),
            .I(N__35544));
    InMux I__7509 (
            .O(N__35544),
            .I(N__35541));
    LocalMux I__7508 (
            .O(N__35541),
            .I(\nx.n2954 ));
    InMux I__7507 (
            .O(N__35538),
            .I(\nx.n11050 ));
    CascadeMux I__7506 (
            .O(N__35535),
            .I(N__35532));
    InMux I__7505 (
            .O(N__35532),
            .I(N__35529));
    LocalMux I__7504 (
            .O(N__35529),
            .I(N__35525));
    InMux I__7503 (
            .O(N__35528),
            .I(N__35522));
    Odrv4 I__7502 (
            .O(N__35525),
            .I(\nx.n2886 ));
    LocalMux I__7501 (
            .O(N__35522),
            .I(\nx.n2886 ));
    CascadeMux I__7500 (
            .O(N__35517),
            .I(N__35512));
    CascadeMux I__7499 (
            .O(N__35516),
            .I(N__35509));
    InMux I__7498 (
            .O(N__35515),
            .I(N__35506));
    InMux I__7497 (
            .O(N__35512),
            .I(N__35503));
    InMux I__7496 (
            .O(N__35509),
            .I(N__35500));
    LocalMux I__7495 (
            .O(N__35506),
            .I(N__35497));
    LocalMux I__7494 (
            .O(N__35503),
            .I(N__35494));
    LocalMux I__7493 (
            .O(N__35500),
            .I(N__35491));
    Span4Mux_v I__7492 (
            .O(N__35497),
            .I(N__35486));
    Span4Mux_h I__7491 (
            .O(N__35494),
            .I(N__35486));
    Odrv4 I__7490 (
            .O(N__35491),
            .I(\nx.n2902 ));
    Odrv4 I__7489 (
            .O(N__35486),
            .I(\nx.n2902 ));
    CascadeMux I__7488 (
            .O(N__35481),
            .I(N__35478));
    InMux I__7487 (
            .O(N__35478),
            .I(N__35475));
    LocalMux I__7486 (
            .O(N__35475),
            .I(N__35472));
    Span4Mux_v I__7485 (
            .O(N__35472),
            .I(N__35469));
    Odrv4 I__7484 (
            .O(N__35469),
            .I(\nx.n2969 ));
    InMux I__7483 (
            .O(N__35466),
            .I(bfn_14_20_0_));
    CascadeMux I__7482 (
            .O(N__35463),
            .I(N__35459));
    InMux I__7481 (
            .O(N__35462),
            .I(N__35456));
    InMux I__7480 (
            .O(N__35459),
            .I(N__35453));
    LocalMux I__7479 (
            .O(N__35456),
            .I(N__35450));
    LocalMux I__7478 (
            .O(N__35453),
            .I(N__35446));
    Span4Mux_v I__7477 (
            .O(N__35450),
            .I(N__35443));
    InMux I__7476 (
            .O(N__35449),
            .I(N__35440));
    Span4Mux_h I__7475 (
            .O(N__35446),
            .I(N__35437));
    Odrv4 I__7474 (
            .O(N__35443),
            .I(\nx.n2901 ));
    LocalMux I__7473 (
            .O(N__35440),
            .I(\nx.n2901 ));
    Odrv4 I__7472 (
            .O(N__35437),
            .I(\nx.n2901 ));
    CascadeMux I__7471 (
            .O(N__35430),
            .I(N__35427));
    InMux I__7470 (
            .O(N__35427),
            .I(N__35424));
    LocalMux I__7469 (
            .O(N__35424),
            .I(N__35421));
    Span4Mux_v I__7468 (
            .O(N__35421),
            .I(N__35418));
    Odrv4 I__7467 (
            .O(N__35418),
            .I(\nx.n2968 ));
    InMux I__7466 (
            .O(N__35415),
            .I(\nx.n11036 ));
    InMux I__7465 (
            .O(N__35412),
            .I(N__35408));
    CascadeMux I__7464 (
            .O(N__35411),
            .I(N__35405));
    LocalMux I__7463 (
            .O(N__35408),
            .I(N__35402));
    InMux I__7462 (
            .O(N__35405),
            .I(N__35398));
    Span4Mux_v I__7461 (
            .O(N__35402),
            .I(N__35395));
    InMux I__7460 (
            .O(N__35401),
            .I(N__35392));
    LocalMux I__7459 (
            .O(N__35398),
            .I(N__35389));
    Odrv4 I__7458 (
            .O(N__35395),
            .I(\nx.n2900 ));
    LocalMux I__7457 (
            .O(N__35392),
            .I(\nx.n2900 ));
    Odrv12 I__7456 (
            .O(N__35389),
            .I(\nx.n2900 ));
    InMux I__7455 (
            .O(N__35382),
            .I(N__35379));
    LocalMux I__7454 (
            .O(N__35379),
            .I(N__35376));
    Odrv4 I__7453 (
            .O(N__35376),
            .I(\nx.n2967 ));
    InMux I__7452 (
            .O(N__35373),
            .I(\nx.n11037 ));
    CascadeMux I__7451 (
            .O(N__35370),
            .I(N__35366));
    InMux I__7450 (
            .O(N__35369),
            .I(N__35363));
    InMux I__7449 (
            .O(N__35366),
            .I(N__35360));
    LocalMux I__7448 (
            .O(N__35363),
            .I(N__35357));
    LocalMux I__7447 (
            .O(N__35360),
            .I(N__35353));
    Span4Mux_h I__7446 (
            .O(N__35357),
            .I(N__35350));
    InMux I__7445 (
            .O(N__35356),
            .I(N__35347));
    Span4Mux_h I__7444 (
            .O(N__35353),
            .I(N__35344));
    Span4Mux_v I__7443 (
            .O(N__35350),
            .I(N__35341));
    LocalMux I__7442 (
            .O(N__35347),
            .I(\nx.n2899 ));
    Odrv4 I__7441 (
            .O(N__35344),
            .I(\nx.n2899 ));
    Odrv4 I__7440 (
            .O(N__35341),
            .I(\nx.n2899 ));
    InMux I__7439 (
            .O(N__35334),
            .I(N__35331));
    LocalMux I__7438 (
            .O(N__35331),
            .I(N__35328));
    Span4Mux_h I__7437 (
            .O(N__35328),
            .I(N__35325));
    Odrv4 I__7436 (
            .O(N__35325),
            .I(\nx.n2966 ));
    InMux I__7435 (
            .O(N__35322),
            .I(\nx.n11038 ));
    InMux I__7434 (
            .O(N__35319),
            .I(N__35316));
    LocalMux I__7433 (
            .O(N__35316),
            .I(N__35313));
    Odrv12 I__7432 (
            .O(N__35313),
            .I(\nx.n2965 ));
    InMux I__7431 (
            .O(N__35310),
            .I(\nx.n11039 ));
    InMux I__7430 (
            .O(N__35307),
            .I(N__35304));
    LocalMux I__7429 (
            .O(N__35304),
            .I(N__35301));
    Span4Mux_v I__7428 (
            .O(N__35301),
            .I(N__35298));
    Odrv4 I__7427 (
            .O(N__35298),
            .I(\nx.n2964 ));
    InMux I__7426 (
            .O(N__35295),
            .I(\nx.n11040 ));
    InMux I__7425 (
            .O(N__35292),
            .I(\nx.n11041 ));
    CascadeMux I__7424 (
            .O(N__35289),
            .I(N__35286));
    InMux I__7423 (
            .O(N__35286),
            .I(N__35283));
    LocalMux I__7422 (
            .O(N__35283),
            .I(N__35279));
    InMux I__7421 (
            .O(N__35282),
            .I(N__35276));
    Odrv4 I__7420 (
            .O(N__35279),
            .I(\nx.n2895 ));
    LocalMux I__7419 (
            .O(N__35276),
            .I(\nx.n2895 ));
    InMux I__7418 (
            .O(N__35271),
            .I(N__35268));
    LocalMux I__7417 (
            .O(N__35268),
            .I(N__35265));
    Odrv4 I__7416 (
            .O(N__35265),
            .I(\nx.n2962 ));
    InMux I__7415 (
            .O(N__35262),
            .I(\nx.n11042 ));
    InMux I__7414 (
            .O(N__35259),
            .I(N__35254));
    InMux I__7413 (
            .O(N__35258),
            .I(N__35251));
    InMux I__7412 (
            .O(N__35257),
            .I(N__35248));
    LocalMux I__7411 (
            .O(N__35254),
            .I(N__35245));
    LocalMux I__7410 (
            .O(N__35251),
            .I(N__35242));
    LocalMux I__7409 (
            .O(N__35248),
            .I(N__35239));
    Span4Mux_h I__7408 (
            .O(N__35245),
            .I(N__35234));
    Span4Mux_h I__7407 (
            .O(N__35242),
            .I(N__35234));
    Span4Mux_h I__7406 (
            .O(N__35239),
            .I(N__35229));
    Span4Mux_v I__7405 (
            .O(N__35234),
            .I(N__35226));
    InMux I__7404 (
            .O(N__35233),
            .I(N__35223));
    InMux I__7403 (
            .O(N__35232),
            .I(N__35220));
    Span4Mux_h I__7402 (
            .O(N__35229),
            .I(N__35217));
    Span4Mux_h I__7401 (
            .O(N__35226),
            .I(N__35214));
    LocalMux I__7400 (
            .O(N__35223),
            .I(\nx.bit_ctr_6 ));
    LocalMux I__7399 (
            .O(N__35220),
            .I(\nx.bit_ctr_6 ));
    Odrv4 I__7398 (
            .O(N__35217),
            .I(\nx.bit_ctr_6 ));
    Odrv4 I__7397 (
            .O(N__35214),
            .I(\nx.bit_ctr_6 ));
    InMux I__7396 (
            .O(N__35205),
            .I(N__35202));
    LocalMux I__7395 (
            .O(N__35202),
            .I(N__35199));
    Span4Mux_h I__7394 (
            .O(N__35199),
            .I(N__35196));
    Odrv4 I__7393 (
            .O(N__35196),
            .I(\nx.n2977 ));
    InMux I__7392 (
            .O(N__35193),
            .I(bfn_14_19_0_));
    CascadeMux I__7391 (
            .O(N__35190),
            .I(N__35187));
    InMux I__7390 (
            .O(N__35187),
            .I(N__35182));
    InMux I__7389 (
            .O(N__35186),
            .I(N__35179));
    InMux I__7388 (
            .O(N__35185),
            .I(N__35176));
    LocalMux I__7387 (
            .O(N__35182),
            .I(N__35173));
    LocalMux I__7386 (
            .O(N__35179),
            .I(\nx.n2909 ));
    LocalMux I__7385 (
            .O(N__35176),
            .I(\nx.n2909 ));
    Odrv12 I__7384 (
            .O(N__35173),
            .I(\nx.n2909 ));
    InMux I__7383 (
            .O(N__35166),
            .I(N__35163));
    LocalMux I__7382 (
            .O(N__35163),
            .I(N__35160));
    Span4Mux_h I__7381 (
            .O(N__35160),
            .I(N__35157));
    Odrv4 I__7380 (
            .O(N__35157),
            .I(\nx.n2976 ));
    InMux I__7379 (
            .O(N__35154),
            .I(\nx.n11028 ));
    InMux I__7378 (
            .O(N__35151),
            .I(N__35147));
    CascadeMux I__7377 (
            .O(N__35150),
            .I(N__35143));
    LocalMux I__7376 (
            .O(N__35147),
            .I(N__35140));
    CascadeMux I__7375 (
            .O(N__35146),
            .I(N__35137));
    InMux I__7374 (
            .O(N__35143),
            .I(N__35134));
    Span4Mux_v I__7373 (
            .O(N__35140),
            .I(N__35131));
    InMux I__7372 (
            .O(N__35137),
            .I(N__35128));
    LocalMux I__7371 (
            .O(N__35134),
            .I(N__35121));
    Sp12to4 I__7370 (
            .O(N__35131),
            .I(N__35121));
    LocalMux I__7369 (
            .O(N__35128),
            .I(N__35121));
    Odrv12 I__7368 (
            .O(N__35121),
            .I(\nx.n2908 ));
    InMux I__7367 (
            .O(N__35118),
            .I(N__35115));
    LocalMux I__7366 (
            .O(N__35115),
            .I(N__35112));
    Odrv12 I__7365 (
            .O(N__35112),
            .I(\nx.n2975 ));
    InMux I__7364 (
            .O(N__35109),
            .I(\nx.n11029 ));
    InMux I__7363 (
            .O(N__35106),
            .I(N__35100));
    InMux I__7362 (
            .O(N__35105),
            .I(N__35100));
    LocalMux I__7361 (
            .O(N__35100),
            .I(N__35096));
    CascadeMux I__7360 (
            .O(N__35099),
            .I(N__35093));
    Span4Mux_v I__7359 (
            .O(N__35096),
            .I(N__35090));
    InMux I__7358 (
            .O(N__35093),
            .I(N__35087));
    Sp12to4 I__7357 (
            .O(N__35090),
            .I(N__35082));
    LocalMux I__7356 (
            .O(N__35087),
            .I(N__35082));
    Odrv12 I__7355 (
            .O(N__35082),
            .I(\nx.n2907 ));
    InMux I__7354 (
            .O(N__35079),
            .I(N__35076));
    LocalMux I__7353 (
            .O(N__35076),
            .I(\nx.n2974 ));
    InMux I__7352 (
            .O(N__35073),
            .I(\nx.n11030 ));
    CascadeMux I__7351 (
            .O(N__35070),
            .I(N__35066));
    InMux I__7350 (
            .O(N__35069),
            .I(N__35062));
    InMux I__7349 (
            .O(N__35066),
            .I(N__35059));
    CascadeMux I__7348 (
            .O(N__35065),
            .I(N__35056));
    LocalMux I__7347 (
            .O(N__35062),
            .I(N__35051));
    LocalMux I__7346 (
            .O(N__35059),
            .I(N__35051));
    InMux I__7345 (
            .O(N__35056),
            .I(N__35048));
    Span4Mux_h I__7344 (
            .O(N__35051),
            .I(N__35045));
    LocalMux I__7343 (
            .O(N__35048),
            .I(\nx.n2906 ));
    Odrv4 I__7342 (
            .O(N__35045),
            .I(\nx.n2906 ));
    InMux I__7341 (
            .O(N__35040),
            .I(N__35037));
    LocalMux I__7340 (
            .O(N__35037),
            .I(N__35034));
    Odrv4 I__7339 (
            .O(N__35034),
            .I(\nx.n2973 ));
    InMux I__7338 (
            .O(N__35031),
            .I(\nx.n11031 ));
    InMux I__7337 (
            .O(N__35028),
            .I(N__35021));
    InMux I__7336 (
            .O(N__35027),
            .I(N__35021));
    InMux I__7335 (
            .O(N__35026),
            .I(N__35018));
    LocalMux I__7334 (
            .O(N__35021),
            .I(\nx.n2905 ));
    LocalMux I__7333 (
            .O(N__35018),
            .I(\nx.n2905 ));
    CascadeMux I__7332 (
            .O(N__35013),
            .I(N__35010));
    InMux I__7331 (
            .O(N__35010),
            .I(N__35007));
    LocalMux I__7330 (
            .O(N__35007),
            .I(\nx.n2972 ));
    InMux I__7329 (
            .O(N__35004),
            .I(\nx.n11032 ));
    CascadeMux I__7328 (
            .O(N__35001),
            .I(N__34998));
    InMux I__7327 (
            .O(N__34998),
            .I(N__34995));
    LocalMux I__7326 (
            .O(N__34995),
            .I(N__34992));
    Odrv4 I__7325 (
            .O(N__34992),
            .I(\nx.n2971 ));
    InMux I__7324 (
            .O(N__34989),
            .I(\nx.n11033 ));
    InMux I__7323 (
            .O(N__34986),
            .I(\nx.n11034 ));
    CascadeMux I__7322 (
            .O(N__34983),
            .I(N__34980));
    InMux I__7321 (
            .O(N__34980),
            .I(N__34977));
    LocalMux I__7320 (
            .O(N__34977),
            .I(N__34974));
    Span4Mux_h I__7319 (
            .O(N__34974),
            .I(N__34970));
    InMux I__7318 (
            .O(N__34973),
            .I(N__34967));
    Odrv4 I__7317 (
            .O(N__34970),
            .I(\nx.n2291 ));
    LocalMux I__7316 (
            .O(N__34967),
            .I(\nx.n2291 ));
    InMux I__7315 (
            .O(N__34962),
            .I(\nx.n10917 ));
    InMux I__7314 (
            .O(N__34959),
            .I(N__34955));
    InMux I__7313 (
            .O(N__34958),
            .I(N__34952));
    LocalMux I__7312 (
            .O(N__34955),
            .I(N__34947));
    LocalMux I__7311 (
            .O(N__34952),
            .I(N__34947));
    Odrv12 I__7310 (
            .O(N__34947),
            .I(\nx.n3006 ));
    InMux I__7309 (
            .O(N__34944),
            .I(N__34940));
    InMux I__7308 (
            .O(N__34943),
            .I(N__34937));
    LocalMux I__7307 (
            .O(N__34940),
            .I(N__34931));
    LocalMux I__7306 (
            .O(N__34937),
            .I(N__34931));
    InMux I__7305 (
            .O(N__34936),
            .I(N__34928));
    Odrv12 I__7304 (
            .O(N__34931),
            .I(\nx.n3004 ));
    LocalMux I__7303 (
            .O(N__34928),
            .I(\nx.n3004 ));
    CascadeMux I__7302 (
            .O(N__34923),
            .I(\nx.n3006_cascade_ ));
    InMux I__7301 (
            .O(N__34920),
            .I(N__34917));
    LocalMux I__7300 (
            .O(N__34917),
            .I(N__34914));
    Span4Mux_h I__7299 (
            .O(N__34914),
            .I(N__34911));
    Odrv4 I__7298 (
            .O(N__34911),
            .I(\nx.n43 ));
    InMux I__7297 (
            .O(N__34908),
            .I(N__34904));
    InMux I__7296 (
            .O(N__34907),
            .I(N__34901));
    LocalMux I__7295 (
            .O(N__34904),
            .I(N__34896));
    LocalMux I__7294 (
            .O(N__34901),
            .I(N__34896));
    Span4Mux_h I__7293 (
            .O(N__34896),
            .I(N__34892));
    InMux I__7292 (
            .O(N__34895),
            .I(N__34889));
    Odrv4 I__7291 (
            .O(N__34892),
            .I(\nx.n2999 ));
    LocalMux I__7290 (
            .O(N__34889),
            .I(\nx.n2999 ));
    InMux I__7289 (
            .O(N__34884),
            .I(N__34879));
    CascadeMux I__7288 (
            .O(N__34883),
            .I(N__34876));
    CascadeMux I__7287 (
            .O(N__34882),
            .I(N__34873));
    LocalMux I__7286 (
            .O(N__34879),
            .I(N__34870));
    InMux I__7285 (
            .O(N__34876),
            .I(N__34867));
    InMux I__7284 (
            .O(N__34873),
            .I(N__34864));
    Span4Mux_h I__7283 (
            .O(N__34870),
            .I(N__34859));
    LocalMux I__7282 (
            .O(N__34867),
            .I(N__34859));
    LocalMux I__7281 (
            .O(N__34864),
            .I(N__34856));
    Odrv4 I__7280 (
            .O(N__34859),
            .I(\nx.n2797 ));
    Odrv4 I__7279 (
            .O(N__34856),
            .I(\nx.n2797 ));
    InMux I__7278 (
            .O(N__34851),
            .I(N__34848));
    LocalMux I__7277 (
            .O(N__34848),
            .I(N__34845));
    Span4Mux_h I__7276 (
            .O(N__34845),
            .I(N__34842));
    Span4Mux_h I__7275 (
            .O(N__34842),
            .I(N__34839));
    Odrv4 I__7274 (
            .O(N__34839),
            .I(\nx.n2864 ));
    CascadeMux I__7273 (
            .O(N__34836),
            .I(\nx.n2896_cascade_ ));
    CascadeMux I__7272 (
            .O(N__34833),
            .I(\nx.n43_adj_763_cascade_ ));
    InMux I__7271 (
            .O(N__34830),
            .I(N__34827));
    LocalMux I__7270 (
            .O(N__34827),
            .I(N__34824));
    Span4Mux_h I__7269 (
            .O(N__34824),
            .I(N__34821));
    Odrv4 I__7268 (
            .O(N__34821),
            .I(\nx.n38_adj_762 ));
    InMux I__7267 (
            .O(N__34818),
            .I(N__34814));
    CascadeMux I__7266 (
            .O(N__34817),
            .I(N__34811));
    LocalMux I__7265 (
            .O(N__34814),
            .I(N__34808));
    InMux I__7264 (
            .O(N__34811),
            .I(N__34805));
    Span4Mux_v I__7263 (
            .O(N__34808),
            .I(N__34801));
    LocalMux I__7262 (
            .O(N__34805),
            .I(N__34798));
    InMux I__7261 (
            .O(N__34804),
            .I(N__34795));
    Span4Mux_h I__7260 (
            .O(N__34801),
            .I(N__34790));
    Span4Mux_h I__7259 (
            .O(N__34798),
            .I(N__34790));
    LocalMux I__7258 (
            .O(N__34795),
            .I(\nx.n2806 ));
    Odrv4 I__7257 (
            .O(N__34790),
            .I(\nx.n2806 ));
    CascadeMux I__7256 (
            .O(N__34785),
            .I(N__34782));
    InMux I__7255 (
            .O(N__34782),
            .I(N__34779));
    LocalMux I__7254 (
            .O(N__34779),
            .I(N__34776));
    Span4Mux_v I__7253 (
            .O(N__34776),
            .I(N__34773));
    Span4Mux_h I__7252 (
            .O(N__34773),
            .I(N__34770));
    Odrv4 I__7251 (
            .O(N__34770),
            .I(\nx.n2873 ));
    InMux I__7250 (
            .O(N__34767),
            .I(N__34764));
    LocalMux I__7249 (
            .O(N__34764),
            .I(N__34761));
    Span4Mux_v I__7248 (
            .O(N__34761),
            .I(N__34757));
    InMux I__7247 (
            .O(N__34760),
            .I(N__34754));
    Odrv4 I__7246 (
            .O(N__34757),
            .I(\nx.n2299 ));
    LocalMux I__7245 (
            .O(N__34754),
            .I(\nx.n2299 ));
    InMux I__7244 (
            .O(N__34749),
            .I(N__34746));
    LocalMux I__7243 (
            .O(N__34746),
            .I(N__34743));
    Odrv4 I__7242 (
            .O(N__34743),
            .I(\nx.n2366 ));
    InMux I__7241 (
            .O(N__34740),
            .I(\nx.n10909 ));
    InMux I__7240 (
            .O(N__34737),
            .I(\nx.n10910 ));
    InMux I__7239 (
            .O(N__34734),
            .I(\nx.n10911 ));
    CascadeMux I__7238 (
            .O(N__34731),
            .I(N__34727));
    CascadeMux I__7237 (
            .O(N__34730),
            .I(N__34724));
    InMux I__7236 (
            .O(N__34727),
            .I(N__34721));
    InMux I__7235 (
            .O(N__34724),
            .I(N__34718));
    LocalMux I__7234 (
            .O(N__34721),
            .I(N__34714));
    LocalMux I__7233 (
            .O(N__34718),
            .I(N__34711));
    InMux I__7232 (
            .O(N__34717),
            .I(N__34708));
    Span4Mux_v I__7231 (
            .O(N__34714),
            .I(N__34701));
    Span4Mux_v I__7230 (
            .O(N__34711),
            .I(N__34701));
    LocalMux I__7229 (
            .O(N__34708),
            .I(N__34701));
    Span4Mux_h I__7228 (
            .O(N__34701),
            .I(N__34698));
    Odrv4 I__7227 (
            .O(N__34698),
            .I(\nx.n2296 ));
    InMux I__7226 (
            .O(N__34695),
            .I(N__34692));
    LocalMux I__7225 (
            .O(N__34692),
            .I(N__34689));
    Odrv12 I__7224 (
            .O(N__34689),
            .I(\nx.n2363 ));
    InMux I__7223 (
            .O(N__34686),
            .I(\nx.n10912 ));
    InMux I__7222 (
            .O(N__34683),
            .I(\nx.n10913 ));
    CascadeMux I__7221 (
            .O(N__34680),
            .I(N__34675));
    CascadeMux I__7220 (
            .O(N__34679),
            .I(N__34672));
    InMux I__7219 (
            .O(N__34678),
            .I(N__34667));
    InMux I__7218 (
            .O(N__34675),
            .I(N__34667));
    InMux I__7217 (
            .O(N__34672),
            .I(N__34664));
    LocalMux I__7216 (
            .O(N__34667),
            .I(N__34661));
    LocalMux I__7215 (
            .O(N__34664),
            .I(\nx.n2294 ));
    Odrv4 I__7214 (
            .O(N__34661),
            .I(\nx.n2294 ));
    InMux I__7213 (
            .O(N__34656),
            .I(N__34653));
    LocalMux I__7212 (
            .O(N__34653),
            .I(N__34650));
    Odrv4 I__7211 (
            .O(N__34650),
            .I(\nx.n2361 ));
    InMux I__7210 (
            .O(N__34647),
            .I(bfn_13_28_0_));
    CascadeMux I__7209 (
            .O(N__34644),
            .I(N__34639));
    InMux I__7208 (
            .O(N__34643),
            .I(N__34636));
    InMux I__7207 (
            .O(N__34642),
            .I(N__34633));
    InMux I__7206 (
            .O(N__34639),
            .I(N__34630));
    LocalMux I__7205 (
            .O(N__34636),
            .I(N__34627));
    LocalMux I__7204 (
            .O(N__34633),
            .I(\nx.n2293 ));
    LocalMux I__7203 (
            .O(N__34630),
            .I(\nx.n2293 ));
    Odrv4 I__7202 (
            .O(N__34627),
            .I(\nx.n2293 ));
    InMux I__7201 (
            .O(N__34620),
            .I(N__34617));
    LocalMux I__7200 (
            .O(N__34617),
            .I(\nx.n2360 ));
    InMux I__7199 (
            .O(N__34614),
            .I(\nx.n10915 ));
    CascadeMux I__7198 (
            .O(N__34611),
            .I(N__34608));
    InMux I__7197 (
            .O(N__34608),
            .I(N__34605));
    LocalMux I__7196 (
            .O(N__34605),
            .I(N__34602));
    Span4Mux_h I__7195 (
            .O(N__34602),
            .I(N__34597));
    InMux I__7194 (
            .O(N__34601),
            .I(N__34592));
    InMux I__7193 (
            .O(N__34600),
            .I(N__34592));
    Odrv4 I__7192 (
            .O(N__34597),
            .I(\nx.n2292 ));
    LocalMux I__7191 (
            .O(N__34592),
            .I(\nx.n2292 ));
    InMux I__7190 (
            .O(N__34587),
            .I(N__34584));
    LocalMux I__7189 (
            .O(N__34584),
            .I(N__34581));
    Odrv4 I__7188 (
            .O(N__34581),
            .I(\nx.n2359 ));
    InMux I__7187 (
            .O(N__34578),
            .I(\nx.n10916 ));
    InMux I__7186 (
            .O(N__34575),
            .I(\nx.n10901 ));
    CascadeMux I__7185 (
            .O(N__34572),
            .I(N__34567));
    InMux I__7184 (
            .O(N__34571),
            .I(N__34564));
    InMux I__7183 (
            .O(N__34570),
            .I(N__34561));
    InMux I__7182 (
            .O(N__34567),
            .I(N__34558));
    LocalMux I__7181 (
            .O(N__34564),
            .I(N__34555));
    LocalMux I__7180 (
            .O(N__34561),
            .I(\nx.n2306 ));
    LocalMux I__7179 (
            .O(N__34558),
            .I(\nx.n2306 ));
    Odrv4 I__7178 (
            .O(N__34555),
            .I(\nx.n2306 ));
    CascadeMux I__7177 (
            .O(N__34548),
            .I(N__34545));
    InMux I__7176 (
            .O(N__34545),
            .I(N__34542));
    LocalMux I__7175 (
            .O(N__34542),
            .I(\nx.n2373 ));
    InMux I__7174 (
            .O(N__34539),
            .I(\nx.n10902 ));
    CascadeMux I__7173 (
            .O(N__34536),
            .I(N__34532));
    CascadeMux I__7172 (
            .O(N__34535),
            .I(N__34529));
    InMux I__7171 (
            .O(N__34532),
            .I(N__34525));
    InMux I__7170 (
            .O(N__34529),
            .I(N__34522));
    InMux I__7169 (
            .O(N__34528),
            .I(N__34519));
    LocalMux I__7168 (
            .O(N__34525),
            .I(N__34516));
    LocalMux I__7167 (
            .O(N__34522),
            .I(\nx.n2305 ));
    LocalMux I__7166 (
            .O(N__34519),
            .I(\nx.n2305 ));
    Odrv4 I__7165 (
            .O(N__34516),
            .I(\nx.n2305 ));
    InMux I__7164 (
            .O(N__34509),
            .I(N__34506));
    LocalMux I__7163 (
            .O(N__34506),
            .I(\nx.n2372 ));
    InMux I__7162 (
            .O(N__34503),
            .I(\nx.n10903 ));
    CascadeMux I__7161 (
            .O(N__34500),
            .I(N__34495));
    InMux I__7160 (
            .O(N__34499),
            .I(N__34492));
    InMux I__7159 (
            .O(N__34498),
            .I(N__34489));
    InMux I__7158 (
            .O(N__34495),
            .I(N__34486));
    LocalMux I__7157 (
            .O(N__34492),
            .I(\nx.n2304 ));
    LocalMux I__7156 (
            .O(N__34489),
            .I(\nx.n2304 ));
    LocalMux I__7155 (
            .O(N__34486),
            .I(\nx.n2304 ));
    InMux I__7154 (
            .O(N__34479),
            .I(N__34476));
    LocalMux I__7153 (
            .O(N__34476),
            .I(\nx.n2371 ));
    InMux I__7152 (
            .O(N__34473),
            .I(\nx.n10904 ));
    CascadeMux I__7151 (
            .O(N__34470),
            .I(N__34466));
    InMux I__7150 (
            .O(N__34469),
            .I(N__34463));
    InMux I__7149 (
            .O(N__34466),
            .I(N__34460));
    LocalMux I__7148 (
            .O(N__34463),
            .I(\nx.n2303 ));
    LocalMux I__7147 (
            .O(N__34460),
            .I(\nx.n2303 ));
    InMux I__7146 (
            .O(N__34455),
            .I(N__34452));
    LocalMux I__7145 (
            .O(N__34452),
            .I(\nx.n2370 ));
    InMux I__7144 (
            .O(N__34449),
            .I(\nx.n10905 ));
    CascadeMux I__7143 (
            .O(N__34446),
            .I(N__34443));
    InMux I__7142 (
            .O(N__34443),
            .I(N__34439));
    InMux I__7141 (
            .O(N__34442),
            .I(N__34436));
    LocalMux I__7140 (
            .O(N__34439),
            .I(N__34433));
    LocalMux I__7139 (
            .O(N__34436),
            .I(\nx.n2302 ));
    Odrv4 I__7138 (
            .O(N__34433),
            .I(\nx.n2302 ));
    InMux I__7137 (
            .O(N__34428),
            .I(N__34425));
    LocalMux I__7136 (
            .O(N__34425),
            .I(N__34422));
    Odrv4 I__7135 (
            .O(N__34422),
            .I(\nx.n2369 ));
    InMux I__7134 (
            .O(N__34419),
            .I(bfn_13_27_0_));
    InMux I__7133 (
            .O(N__34416),
            .I(\nx.n10907 ));
    InMux I__7132 (
            .O(N__34413),
            .I(N__34409));
    CascadeMux I__7131 (
            .O(N__34412),
            .I(N__34406));
    LocalMux I__7130 (
            .O(N__34409),
            .I(N__34402));
    InMux I__7129 (
            .O(N__34406),
            .I(N__34399));
    InMux I__7128 (
            .O(N__34405),
            .I(N__34396));
    Odrv4 I__7127 (
            .O(N__34402),
            .I(\nx.n2300 ));
    LocalMux I__7126 (
            .O(N__34399),
            .I(\nx.n2300 ));
    LocalMux I__7125 (
            .O(N__34396),
            .I(\nx.n2300 ));
    InMux I__7124 (
            .O(N__34389),
            .I(N__34386));
    LocalMux I__7123 (
            .O(N__34386),
            .I(N__34383));
    Odrv4 I__7122 (
            .O(N__34383),
            .I(\nx.n2367 ));
    InMux I__7121 (
            .O(N__34380),
            .I(\nx.n10908 ));
    CascadeMux I__7120 (
            .O(N__34377),
            .I(\nx.n2398_cascade_ ));
    InMux I__7119 (
            .O(N__34374),
            .I(N__34371));
    LocalMux I__7118 (
            .O(N__34371),
            .I(N__34368));
    Odrv4 I__7117 (
            .O(N__34368),
            .I(\nx.n31_adj_700 ));
    InMux I__7116 (
            .O(N__34365),
            .I(N__34362));
    LocalMux I__7115 (
            .O(N__34362),
            .I(\nx.n32_adj_698 ));
    CascadeMux I__7114 (
            .O(N__34359),
            .I(N__34356));
    InMux I__7113 (
            .O(N__34356),
            .I(N__34353));
    LocalMux I__7112 (
            .O(N__34353),
            .I(\nx.n33_adj_699 ));
    InMux I__7111 (
            .O(N__34350),
            .I(N__34347));
    LocalMux I__7110 (
            .O(N__34347),
            .I(\nx.n34_adj_697 ));
    CascadeMux I__7109 (
            .O(N__34344),
            .I(\nx.n2324_cascade_ ));
    InMux I__7108 (
            .O(N__34341),
            .I(N__34337));
    InMux I__7107 (
            .O(N__34340),
            .I(N__34334));
    LocalMux I__7106 (
            .O(N__34337),
            .I(N__34330));
    LocalMux I__7105 (
            .O(N__34334),
            .I(N__34325));
    InMux I__7104 (
            .O(N__34333),
            .I(N__34322));
    Span4Mux_v I__7103 (
            .O(N__34330),
            .I(N__34319));
    InMux I__7102 (
            .O(N__34329),
            .I(N__34316));
    InMux I__7101 (
            .O(N__34328),
            .I(N__34313));
    Span4Mux_h I__7100 (
            .O(N__34325),
            .I(N__34310));
    LocalMux I__7099 (
            .O(N__34322),
            .I(N__34303));
    Sp12to4 I__7098 (
            .O(N__34319),
            .I(N__34303));
    LocalMux I__7097 (
            .O(N__34316),
            .I(N__34303));
    LocalMux I__7096 (
            .O(N__34313),
            .I(\nx.bit_ctr_12 ));
    Odrv4 I__7095 (
            .O(N__34310),
            .I(\nx.bit_ctr_12 ));
    Odrv12 I__7094 (
            .O(N__34303),
            .I(\nx.bit_ctr_12 ));
    InMux I__7093 (
            .O(N__34296),
            .I(N__34293));
    LocalMux I__7092 (
            .O(N__34293),
            .I(N__34290));
    Odrv4 I__7091 (
            .O(N__34290),
            .I(\nx.n2377 ));
    InMux I__7090 (
            .O(N__34287),
            .I(bfn_13_26_0_));
    CascadeMux I__7089 (
            .O(N__34284),
            .I(N__34281));
    InMux I__7088 (
            .O(N__34281),
            .I(N__34277));
    InMux I__7087 (
            .O(N__34280),
            .I(N__34274));
    LocalMux I__7086 (
            .O(N__34277),
            .I(N__34271));
    LocalMux I__7085 (
            .O(N__34274),
            .I(\nx.n2309 ));
    Odrv4 I__7084 (
            .O(N__34271),
            .I(\nx.n2309 ));
    InMux I__7083 (
            .O(N__34266),
            .I(N__34263));
    LocalMux I__7082 (
            .O(N__34263),
            .I(N__34260));
    Odrv4 I__7081 (
            .O(N__34260),
            .I(\nx.n2376 ));
    InMux I__7080 (
            .O(N__34257),
            .I(\nx.n10899 ));
    CascadeMux I__7079 (
            .O(N__34254),
            .I(N__34251));
    InMux I__7078 (
            .O(N__34251),
            .I(N__34246));
    InMux I__7077 (
            .O(N__34250),
            .I(N__34243));
    InMux I__7076 (
            .O(N__34249),
            .I(N__34240));
    LocalMux I__7075 (
            .O(N__34246),
            .I(N__34237));
    LocalMux I__7074 (
            .O(N__34243),
            .I(\nx.n2308 ));
    LocalMux I__7073 (
            .O(N__34240),
            .I(\nx.n2308 ));
    Odrv4 I__7072 (
            .O(N__34237),
            .I(\nx.n2308 ));
    CascadeMux I__7071 (
            .O(N__34230),
            .I(N__34227));
    InMux I__7070 (
            .O(N__34227),
            .I(N__34224));
    LocalMux I__7069 (
            .O(N__34224),
            .I(N__34221));
    Odrv4 I__7068 (
            .O(N__34221),
            .I(\nx.n2375 ));
    InMux I__7067 (
            .O(N__34218),
            .I(\nx.n10900 ));
    CascadeMux I__7066 (
            .O(N__34215),
            .I(\nx.n2507_cascade_ ));
    CascadeMux I__7065 (
            .O(N__34212),
            .I(\nx.n2603_cascade_ ));
    InMux I__7064 (
            .O(N__34209),
            .I(N__34205));
    CascadeMux I__7063 (
            .O(N__34208),
            .I(N__34202));
    LocalMux I__7062 (
            .O(N__34205),
            .I(N__34198));
    InMux I__7061 (
            .O(N__34202),
            .I(N__34195));
    InMux I__7060 (
            .O(N__34201),
            .I(N__34192));
    Span4Mux_h I__7059 (
            .O(N__34198),
            .I(N__34187));
    LocalMux I__7058 (
            .O(N__34195),
            .I(N__34187));
    LocalMux I__7057 (
            .O(N__34192),
            .I(N__34184));
    Span4Mux_h I__7056 (
            .O(N__34187),
            .I(N__34181));
    Odrv4 I__7055 (
            .O(N__34184),
            .I(\nx.n2702 ));
    Odrv4 I__7054 (
            .O(N__34181),
            .I(\nx.n2702 ));
    InMux I__7053 (
            .O(N__34176),
            .I(N__34173));
    LocalMux I__7052 (
            .O(N__34173),
            .I(N__34169));
    CascadeMux I__7051 (
            .O(N__34172),
            .I(N__34165));
    Span4Mux_h I__7050 (
            .O(N__34169),
            .I(N__34162));
    InMux I__7049 (
            .O(N__34168),
            .I(N__34159));
    InMux I__7048 (
            .O(N__34165),
            .I(N__34156));
    Odrv4 I__7047 (
            .O(N__34162),
            .I(\nx.n2803 ));
    LocalMux I__7046 (
            .O(N__34159),
            .I(\nx.n2803 ));
    LocalMux I__7045 (
            .O(N__34156),
            .I(\nx.n2803 ));
    CascadeMux I__7044 (
            .O(N__34149),
            .I(N__34146));
    InMux I__7043 (
            .O(N__34146),
            .I(N__34143));
    LocalMux I__7042 (
            .O(N__34143),
            .I(N__34140));
    Span4Mux_h I__7041 (
            .O(N__34140),
            .I(N__34137));
    Odrv4 I__7040 (
            .O(N__34137),
            .I(\nx.n2870 ));
    CascadeMux I__7039 (
            .O(N__34134),
            .I(\nx.n2501_cascade_ ));
    InMux I__7038 (
            .O(N__34131),
            .I(N__34128));
    LocalMux I__7037 (
            .O(N__34128),
            .I(N__34123));
    InMux I__7036 (
            .O(N__34127),
            .I(N__34120));
    InMux I__7035 (
            .O(N__34126),
            .I(N__34117));
    Span4Mux_h I__7034 (
            .O(N__34123),
            .I(N__34112));
    LocalMux I__7033 (
            .O(N__34120),
            .I(N__34112));
    LocalMux I__7032 (
            .O(N__34117),
            .I(N__34109));
    Span4Mux_v I__7031 (
            .O(N__34112),
            .I(N__34106));
    Span4Mux_h I__7030 (
            .O(N__34109),
            .I(N__34103));
    Odrv4 I__7029 (
            .O(N__34106),
            .I(\nx.n3085 ));
    Odrv4 I__7028 (
            .O(N__34103),
            .I(\nx.n3085 ));
    InMux I__7027 (
            .O(N__34098),
            .I(N__34095));
    LocalMux I__7026 (
            .O(N__34095),
            .I(N__34092));
    Span4Mux_h I__7025 (
            .O(N__34092),
            .I(N__34089));
    Span4Mux_h I__7024 (
            .O(N__34089),
            .I(N__34086));
    Odrv4 I__7023 (
            .O(N__34086),
            .I(\nx.n3152 ));
    InMux I__7022 (
            .O(N__34083),
            .I(\nx.n11103 ));
    InMux I__7021 (
            .O(N__34080),
            .I(N__34075));
    InMux I__7020 (
            .O(N__34079),
            .I(N__34072));
    InMux I__7019 (
            .O(N__34078),
            .I(N__34069));
    LocalMux I__7018 (
            .O(N__34075),
            .I(N__34066));
    LocalMux I__7017 (
            .O(N__34072),
            .I(N__34063));
    LocalMux I__7016 (
            .O(N__34069),
            .I(N__34060));
    Span4Mux_v I__7015 (
            .O(N__34066),
            .I(N__34055));
    Span4Mux_v I__7014 (
            .O(N__34063),
            .I(N__34055));
    Span4Mux_h I__7013 (
            .O(N__34060),
            .I(N__34052));
    Odrv4 I__7012 (
            .O(N__34055),
            .I(\nx.n3084 ));
    Odrv4 I__7011 (
            .O(N__34052),
            .I(\nx.n3084 ));
    InMux I__7010 (
            .O(N__34047),
            .I(N__34044));
    LocalMux I__7009 (
            .O(N__34044),
            .I(N__34041));
    Span12Mux_h I__7008 (
            .O(N__34041),
            .I(N__34038));
    Odrv12 I__7007 (
            .O(N__34038),
            .I(\nx.n3151 ));
    InMux I__7006 (
            .O(N__34035),
            .I(\nx.n11104 ));
    CascadeMux I__7005 (
            .O(N__34032),
            .I(N__34029));
    InMux I__7004 (
            .O(N__34029),
            .I(N__34017));
    InMux I__7003 (
            .O(N__34028),
            .I(N__34017));
    InMux I__7002 (
            .O(N__34027),
            .I(N__34017));
    InMux I__7001 (
            .O(N__34026),
            .I(N__34014));
    CascadeMux I__7000 (
            .O(N__34025),
            .I(N__34011));
    CascadeMux I__6999 (
            .O(N__34024),
            .I(N__34008));
    LocalMux I__6998 (
            .O(N__34017),
            .I(N__33998));
    LocalMux I__6997 (
            .O(N__34014),
            .I(N__33995));
    InMux I__6996 (
            .O(N__34011),
            .I(N__33990));
    InMux I__6995 (
            .O(N__34008),
            .I(N__33990));
    CascadeMux I__6994 (
            .O(N__34007),
            .I(N__33981));
    CascadeMux I__6993 (
            .O(N__34006),
            .I(N__33978));
    CascadeMux I__6992 (
            .O(N__34005),
            .I(N__33974));
    CascadeMux I__6991 (
            .O(N__34004),
            .I(N__33969));
    CascadeMux I__6990 (
            .O(N__34003),
            .I(N__33963));
    CascadeMux I__6989 (
            .O(N__34002),
            .I(N__33959));
    CascadeMux I__6988 (
            .O(N__34001),
            .I(N__33956));
    Span4Mux_v I__6987 (
            .O(N__33998),
            .I(N__33948));
    Span4Mux_v I__6986 (
            .O(N__33995),
            .I(N__33948));
    LocalMux I__6985 (
            .O(N__33990),
            .I(N__33948));
    InMux I__6984 (
            .O(N__33989),
            .I(N__33943));
    InMux I__6983 (
            .O(N__33988),
            .I(N__33943));
    InMux I__6982 (
            .O(N__33987),
            .I(N__33930));
    InMux I__6981 (
            .O(N__33986),
            .I(N__33930));
    InMux I__6980 (
            .O(N__33985),
            .I(N__33930));
    InMux I__6979 (
            .O(N__33984),
            .I(N__33930));
    InMux I__6978 (
            .O(N__33981),
            .I(N__33930));
    InMux I__6977 (
            .O(N__33978),
            .I(N__33930));
    InMux I__6976 (
            .O(N__33977),
            .I(N__33915));
    InMux I__6975 (
            .O(N__33974),
            .I(N__33915));
    InMux I__6974 (
            .O(N__33973),
            .I(N__33915));
    InMux I__6973 (
            .O(N__33972),
            .I(N__33915));
    InMux I__6972 (
            .O(N__33969),
            .I(N__33915));
    InMux I__6971 (
            .O(N__33968),
            .I(N__33915));
    InMux I__6970 (
            .O(N__33967),
            .I(N__33915));
    InMux I__6969 (
            .O(N__33966),
            .I(N__33902));
    InMux I__6968 (
            .O(N__33963),
            .I(N__33902));
    InMux I__6967 (
            .O(N__33962),
            .I(N__33902));
    InMux I__6966 (
            .O(N__33959),
            .I(N__33902));
    InMux I__6965 (
            .O(N__33956),
            .I(N__33902));
    InMux I__6964 (
            .O(N__33955),
            .I(N__33902));
    Odrv4 I__6963 (
            .O(N__33948),
            .I(\nx.n3116 ));
    LocalMux I__6962 (
            .O(N__33943),
            .I(\nx.n3116 ));
    LocalMux I__6961 (
            .O(N__33930),
            .I(\nx.n3116 ));
    LocalMux I__6960 (
            .O(N__33915),
            .I(\nx.n3116 ));
    LocalMux I__6959 (
            .O(N__33902),
            .I(\nx.n3116 ));
    CascadeMux I__6958 (
            .O(N__33891),
            .I(N__33888));
    InMux I__6957 (
            .O(N__33888),
            .I(N__33884));
    InMux I__6956 (
            .O(N__33887),
            .I(N__33881));
    LocalMux I__6955 (
            .O(N__33884),
            .I(N__33878));
    LocalMux I__6954 (
            .O(N__33881),
            .I(N__33875));
    Span4Mux_h I__6953 (
            .O(N__33878),
            .I(N__33872));
    Span4Mux_h I__6952 (
            .O(N__33875),
            .I(N__33869));
    Odrv4 I__6951 (
            .O(N__33872),
            .I(\nx.n3083 ));
    Odrv4 I__6950 (
            .O(N__33869),
            .I(\nx.n3083 ));
    InMux I__6949 (
            .O(N__33864),
            .I(\nx.n11105 ));
    InMux I__6948 (
            .O(N__33861),
            .I(N__33858));
    LocalMux I__6947 (
            .O(N__33858),
            .I(N__33855));
    Span4Mux_v I__6946 (
            .O(N__33855),
            .I(N__33852));
    Odrv4 I__6945 (
            .O(N__33852),
            .I(\nx.n13280 ));
    InMux I__6944 (
            .O(N__33849),
            .I(N__33846));
    LocalMux I__6943 (
            .O(N__33846),
            .I(N__33841));
    InMux I__6942 (
            .O(N__33845),
            .I(N__33838));
    CascadeMux I__6941 (
            .O(N__33844),
            .I(N__33835));
    Span4Mux_h I__6940 (
            .O(N__33841),
            .I(N__33832));
    LocalMux I__6939 (
            .O(N__33838),
            .I(N__33829));
    InMux I__6938 (
            .O(N__33835),
            .I(N__33826));
    Odrv4 I__6937 (
            .O(N__33832),
            .I(\nx.n2805 ));
    Odrv4 I__6936 (
            .O(N__33829),
            .I(\nx.n2805 ));
    LocalMux I__6935 (
            .O(N__33826),
            .I(\nx.n2805 ));
    CascadeMux I__6934 (
            .O(N__33819),
            .I(N__33816));
    InMux I__6933 (
            .O(N__33816),
            .I(N__33813));
    LocalMux I__6932 (
            .O(N__33813),
            .I(N__33810));
    Span4Mux_h I__6931 (
            .O(N__33810),
            .I(N__33807));
    Odrv4 I__6930 (
            .O(N__33807),
            .I(\nx.n2872 ));
    CascadeMux I__6929 (
            .O(N__33804),
            .I(N__33800));
    InMux I__6928 (
            .O(N__33803),
            .I(N__33797));
    InMux I__6927 (
            .O(N__33800),
            .I(N__33793));
    LocalMux I__6926 (
            .O(N__33797),
            .I(N__33790));
    InMux I__6925 (
            .O(N__33796),
            .I(N__33787));
    LocalMux I__6924 (
            .O(N__33793),
            .I(N__33784));
    Span4Mux_h I__6923 (
            .O(N__33790),
            .I(N__33779));
    LocalMux I__6922 (
            .O(N__33787),
            .I(N__33779));
    Span4Mux_h I__6921 (
            .O(N__33784),
            .I(N__33776));
    Odrv4 I__6920 (
            .O(N__33779),
            .I(\nx.n2798 ));
    Odrv4 I__6919 (
            .O(N__33776),
            .I(\nx.n2798 ));
    CascadeMux I__6918 (
            .O(N__33771),
            .I(N__33768));
    InMux I__6917 (
            .O(N__33768),
            .I(N__33765));
    LocalMux I__6916 (
            .O(N__33765),
            .I(N__33762));
    Span4Mux_v I__6915 (
            .O(N__33762),
            .I(N__33759));
    Span4Mux_h I__6914 (
            .O(N__33759),
            .I(N__33756));
    Odrv4 I__6913 (
            .O(N__33756),
            .I(\nx.n2865 ));
    InMux I__6912 (
            .O(N__33753),
            .I(N__33749));
    InMux I__6911 (
            .O(N__33752),
            .I(N__33746));
    LocalMux I__6910 (
            .O(N__33749),
            .I(N__33740));
    LocalMux I__6909 (
            .O(N__33746),
            .I(N__33740));
    InMux I__6908 (
            .O(N__33745),
            .I(N__33737));
    Odrv4 I__6907 (
            .O(N__33740),
            .I(\nx.n2986 ));
    LocalMux I__6906 (
            .O(N__33737),
            .I(\nx.n2986 ));
    InMux I__6905 (
            .O(N__33732),
            .I(N__33728));
    InMux I__6904 (
            .O(N__33731),
            .I(N__33725));
    LocalMux I__6903 (
            .O(N__33728),
            .I(N__33720));
    LocalMux I__6902 (
            .O(N__33725),
            .I(N__33720));
    Span4Mux_h I__6901 (
            .O(N__33720),
            .I(N__33716));
    InMux I__6900 (
            .O(N__33719),
            .I(N__33713));
    Odrv4 I__6899 (
            .O(N__33716),
            .I(\nx.n2991 ));
    LocalMux I__6898 (
            .O(N__33713),
            .I(\nx.n2991 ));
    InMux I__6897 (
            .O(N__33708),
            .I(N__33705));
    LocalMux I__6896 (
            .O(N__33705),
            .I(N__33702));
    Span4Mux_h I__6895 (
            .O(N__33702),
            .I(N__33699));
    Odrv4 I__6894 (
            .O(N__33699),
            .I(\nx.n3160 ));
    InMux I__6893 (
            .O(N__33696),
            .I(\nx.n11095 ));
    InMux I__6892 (
            .O(N__33693),
            .I(N__33689));
    CascadeMux I__6891 (
            .O(N__33692),
            .I(N__33686));
    LocalMux I__6890 (
            .O(N__33689),
            .I(N__33682));
    InMux I__6889 (
            .O(N__33686),
            .I(N__33679));
    InMux I__6888 (
            .O(N__33685),
            .I(N__33676));
    Span4Mux_v I__6887 (
            .O(N__33682),
            .I(N__33673));
    LocalMux I__6886 (
            .O(N__33679),
            .I(N__33668));
    LocalMux I__6885 (
            .O(N__33676),
            .I(N__33668));
    Odrv4 I__6884 (
            .O(N__33673),
            .I(\nx.n3092 ));
    Odrv4 I__6883 (
            .O(N__33668),
            .I(\nx.n3092 ));
    InMux I__6882 (
            .O(N__33663),
            .I(N__33660));
    LocalMux I__6881 (
            .O(N__33660),
            .I(N__33657));
    Span4Mux_v I__6880 (
            .O(N__33657),
            .I(N__33654));
    Odrv4 I__6879 (
            .O(N__33654),
            .I(\nx.n3159 ));
    InMux I__6878 (
            .O(N__33651),
            .I(\nx.n11096 ));
    InMux I__6877 (
            .O(N__33648),
            .I(N__33644));
    InMux I__6876 (
            .O(N__33647),
            .I(N__33641));
    LocalMux I__6875 (
            .O(N__33644),
            .I(N__33637));
    LocalMux I__6874 (
            .O(N__33641),
            .I(N__33634));
    InMux I__6873 (
            .O(N__33640),
            .I(N__33631));
    Span4Mux_v I__6872 (
            .O(N__33637),
            .I(N__33626));
    Span4Mux_h I__6871 (
            .O(N__33634),
            .I(N__33626));
    LocalMux I__6870 (
            .O(N__33631),
            .I(N__33623));
    Odrv4 I__6869 (
            .O(N__33626),
            .I(\nx.n3091 ));
    Odrv4 I__6868 (
            .O(N__33623),
            .I(\nx.n3091 ));
    InMux I__6867 (
            .O(N__33618),
            .I(N__33615));
    LocalMux I__6866 (
            .O(N__33615),
            .I(N__33612));
    Span4Mux_v I__6865 (
            .O(N__33612),
            .I(N__33609));
    Odrv4 I__6864 (
            .O(N__33609),
            .I(\nx.n3158 ));
    InMux I__6863 (
            .O(N__33606),
            .I(\nx.n11097 ));
    InMux I__6862 (
            .O(N__33603),
            .I(N__33599));
    InMux I__6861 (
            .O(N__33602),
            .I(N__33596));
    LocalMux I__6860 (
            .O(N__33599),
            .I(N__33592));
    LocalMux I__6859 (
            .O(N__33596),
            .I(N__33589));
    InMux I__6858 (
            .O(N__33595),
            .I(N__33586));
    Span4Mux_v I__6857 (
            .O(N__33592),
            .I(N__33581));
    Span4Mux_h I__6856 (
            .O(N__33589),
            .I(N__33581));
    LocalMux I__6855 (
            .O(N__33586),
            .I(N__33578));
    Odrv4 I__6854 (
            .O(N__33581),
            .I(\nx.n3090 ));
    Odrv4 I__6853 (
            .O(N__33578),
            .I(\nx.n3090 ));
    InMux I__6852 (
            .O(N__33573),
            .I(N__33570));
    LocalMux I__6851 (
            .O(N__33570),
            .I(N__33567));
    Span4Mux_h I__6850 (
            .O(N__33567),
            .I(N__33564));
    Odrv4 I__6849 (
            .O(N__33564),
            .I(\nx.n3157 ));
    InMux I__6848 (
            .O(N__33561),
            .I(\nx.n11098 ));
    InMux I__6847 (
            .O(N__33558),
            .I(N__33555));
    LocalMux I__6846 (
            .O(N__33555),
            .I(N__33550));
    InMux I__6845 (
            .O(N__33554),
            .I(N__33547));
    InMux I__6844 (
            .O(N__33553),
            .I(N__33544));
    Span4Mux_h I__6843 (
            .O(N__33550),
            .I(N__33541));
    LocalMux I__6842 (
            .O(N__33547),
            .I(N__33536));
    LocalMux I__6841 (
            .O(N__33544),
            .I(N__33536));
    Odrv4 I__6840 (
            .O(N__33541),
            .I(\nx.n3089 ));
    Odrv4 I__6839 (
            .O(N__33536),
            .I(\nx.n3089 ));
    InMux I__6838 (
            .O(N__33531),
            .I(N__33528));
    LocalMux I__6837 (
            .O(N__33528),
            .I(N__33525));
    Span4Mux_h I__6836 (
            .O(N__33525),
            .I(N__33522));
    Odrv4 I__6835 (
            .O(N__33522),
            .I(\nx.n3156 ));
    InMux I__6834 (
            .O(N__33519),
            .I(\nx.n11099 ));
    InMux I__6833 (
            .O(N__33516),
            .I(N__33512));
    InMux I__6832 (
            .O(N__33515),
            .I(N__33509));
    LocalMux I__6831 (
            .O(N__33512),
            .I(N__33505));
    LocalMux I__6830 (
            .O(N__33509),
            .I(N__33502));
    InMux I__6829 (
            .O(N__33508),
            .I(N__33499));
    Span4Mux_v I__6828 (
            .O(N__33505),
            .I(N__33496));
    Span4Mux_h I__6827 (
            .O(N__33502),
            .I(N__33493));
    LocalMux I__6826 (
            .O(N__33499),
            .I(N__33490));
    Odrv4 I__6825 (
            .O(N__33496),
            .I(\nx.n3088 ));
    Odrv4 I__6824 (
            .O(N__33493),
            .I(\nx.n3088 ));
    Odrv4 I__6823 (
            .O(N__33490),
            .I(\nx.n3088 ));
    InMux I__6822 (
            .O(N__33483),
            .I(N__33480));
    LocalMux I__6821 (
            .O(N__33480),
            .I(N__33477));
    Span4Mux_h I__6820 (
            .O(N__33477),
            .I(N__33474));
    Odrv4 I__6819 (
            .O(N__33474),
            .I(\nx.n3155 ));
    InMux I__6818 (
            .O(N__33471),
            .I(\nx.n11100 ));
    InMux I__6817 (
            .O(N__33468),
            .I(N__33463));
    InMux I__6816 (
            .O(N__33467),
            .I(N__33460));
    CascadeMux I__6815 (
            .O(N__33466),
            .I(N__33457));
    LocalMux I__6814 (
            .O(N__33463),
            .I(N__33454));
    LocalMux I__6813 (
            .O(N__33460),
            .I(N__33451));
    InMux I__6812 (
            .O(N__33457),
            .I(N__33448));
    Span4Mux_h I__6811 (
            .O(N__33454),
            .I(N__33445));
    Span4Mux_h I__6810 (
            .O(N__33451),
            .I(N__33442));
    LocalMux I__6809 (
            .O(N__33448),
            .I(N__33439));
    Odrv4 I__6808 (
            .O(N__33445),
            .I(\nx.n3087 ));
    Odrv4 I__6807 (
            .O(N__33442),
            .I(\nx.n3087 ));
    Odrv12 I__6806 (
            .O(N__33439),
            .I(\nx.n3087 ));
    InMux I__6805 (
            .O(N__33432),
            .I(N__33429));
    LocalMux I__6804 (
            .O(N__33429),
            .I(N__33426));
    Span4Mux_h I__6803 (
            .O(N__33426),
            .I(N__33423));
    Odrv4 I__6802 (
            .O(N__33423),
            .I(\nx.n3154 ));
    InMux I__6801 (
            .O(N__33420),
            .I(\nx.n11101 ));
    InMux I__6800 (
            .O(N__33417),
            .I(N__33414));
    LocalMux I__6799 (
            .O(N__33414),
            .I(N__33409));
    InMux I__6798 (
            .O(N__33413),
            .I(N__33406));
    InMux I__6797 (
            .O(N__33412),
            .I(N__33403));
    Span4Mux_h I__6796 (
            .O(N__33409),
            .I(N__33400));
    LocalMux I__6795 (
            .O(N__33406),
            .I(N__33397));
    LocalMux I__6794 (
            .O(N__33403),
            .I(N__33394));
    Odrv4 I__6793 (
            .O(N__33400),
            .I(\nx.n3086 ));
    Odrv12 I__6792 (
            .O(N__33397),
            .I(\nx.n3086 ));
    Odrv12 I__6791 (
            .O(N__33394),
            .I(\nx.n3086 ));
    InMux I__6790 (
            .O(N__33387),
            .I(N__33384));
    LocalMux I__6789 (
            .O(N__33384),
            .I(N__33381));
    Span4Mux_h I__6788 (
            .O(N__33381),
            .I(N__33378));
    Odrv4 I__6787 (
            .O(N__33378),
            .I(\nx.n3153 ));
    InMux I__6786 (
            .O(N__33375),
            .I(bfn_13_20_0_));
    CascadeMux I__6785 (
            .O(N__33372),
            .I(N__33369));
    InMux I__6784 (
            .O(N__33369),
            .I(N__33366));
    LocalMux I__6783 (
            .O(N__33366),
            .I(N__33362));
    InMux I__6782 (
            .O(N__33365),
            .I(N__33358));
    Span4Mux_v I__6781 (
            .O(N__33362),
            .I(N__33355));
    InMux I__6780 (
            .O(N__33361),
            .I(N__33352));
    LocalMux I__6779 (
            .O(N__33358),
            .I(\nx.n3100 ));
    Odrv4 I__6778 (
            .O(N__33355),
            .I(\nx.n3100 ));
    LocalMux I__6777 (
            .O(N__33352),
            .I(\nx.n3100 ));
    InMux I__6776 (
            .O(N__33345),
            .I(N__33342));
    LocalMux I__6775 (
            .O(N__33342),
            .I(\nx.n3167 ));
    InMux I__6774 (
            .O(N__33339),
            .I(\nx.n11088 ));
    CascadeMux I__6773 (
            .O(N__33336),
            .I(N__33333));
    InMux I__6772 (
            .O(N__33333),
            .I(N__33330));
    LocalMux I__6771 (
            .O(N__33330),
            .I(N__33325));
    InMux I__6770 (
            .O(N__33329),
            .I(N__33322));
    InMux I__6769 (
            .O(N__33328),
            .I(N__33319));
    Span4Mux_h I__6768 (
            .O(N__33325),
            .I(N__33316));
    LocalMux I__6767 (
            .O(N__33322),
            .I(N__33311));
    LocalMux I__6766 (
            .O(N__33319),
            .I(N__33311));
    Odrv4 I__6765 (
            .O(N__33316),
            .I(\nx.n3099 ));
    Odrv4 I__6764 (
            .O(N__33311),
            .I(\nx.n3099 ));
    InMux I__6763 (
            .O(N__33306),
            .I(N__33303));
    LocalMux I__6762 (
            .O(N__33303),
            .I(\nx.n3166 ));
    InMux I__6761 (
            .O(N__33300),
            .I(\nx.n11089 ));
    CascadeMux I__6760 (
            .O(N__33297),
            .I(N__33294));
    InMux I__6759 (
            .O(N__33294),
            .I(N__33290));
    InMux I__6758 (
            .O(N__33293),
            .I(N__33287));
    LocalMux I__6757 (
            .O(N__33290),
            .I(N__33283));
    LocalMux I__6756 (
            .O(N__33287),
            .I(N__33280));
    InMux I__6755 (
            .O(N__33286),
            .I(N__33277));
    Span4Mux_h I__6754 (
            .O(N__33283),
            .I(N__33274));
    Span4Mux_v I__6753 (
            .O(N__33280),
            .I(N__33271));
    LocalMux I__6752 (
            .O(N__33277),
            .I(\nx.n3098 ));
    Odrv4 I__6751 (
            .O(N__33274),
            .I(\nx.n3098 ));
    Odrv4 I__6750 (
            .O(N__33271),
            .I(\nx.n3098 ));
    InMux I__6749 (
            .O(N__33264),
            .I(N__33261));
    LocalMux I__6748 (
            .O(N__33261),
            .I(N__33258));
    Odrv12 I__6747 (
            .O(N__33258),
            .I(\nx.n3165 ));
    InMux I__6746 (
            .O(N__33255),
            .I(\nx.n11090 ));
    CascadeMux I__6745 (
            .O(N__33252),
            .I(N__33249));
    InMux I__6744 (
            .O(N__33249),
            .I(N__33245));
    InMux I__6743 (
            .O(N__33248),
            .I(N__33242));
    LocalMux I__6742 (
            .O(N__33245),
            .I(N__33239));
    LocalMux I__6741 (
            .O(N__33242),
            .I(N__33235));
    Span4Mux_h I__6740 (
            .O(N__33239),
            .I(N__33232));
    InMux I__6739 (
            .O(N__33238),
            .I(N__33229));
    Odrv4 I__6738 (
            .O(N__33235),
            .I(\nx.n3097 ));
    Odrv4 I__6737 (
            .O(N__33232),
            .I(\nx.n3097 ));
    LocalMux I__6736 (
            .O(N__33229),
            .I(\nx.n3097 ));
    InMux I__6735 (
            .O(N__33222),
            .I(N__33219));
    LocalMux I__6734 (
            .O(N__33219),
            .I(\nx.n3164 ));
    InMux I__6733 (
            .O(N__33216),
            .I(\nx.n11091 ));
    CascadeMux I__6732 (
            .O(N__33213),
            .I(N__33210));
    InMux I__6731 (
            .O(N__33210),
            .I(N__33206));
    InMux I__6730 (
            .O(N__33209),
            .I(N__33202));
    LocalMux I__6729 (
            .O(N__33206),
            .I(N__33199));
    CascadeMux I__6728 (
            .O(N__33205),
            .I(N__33196));
    LocalMux I__6727 (
            .O(N__33202),
            .I(N__33193));
    Span4Mux_h I__6726 (
            .O(N__33199),
            .I(N__33190));
    InMux I__6725 (
            .O(N__33196),
            .I(N__33187));
    Odrv4 I__6724 (
            .O(N__33193),
            .I(\nx.n3096 ));
    Odrv4 I__6723 (
            .O(N__33190),
            .I(\nx.n3096 ));
    LocalMux I__6722 (
            .O(N__33187),
            .I(\nx.n3096 ));
    InMux I__6721 (
            .O(N__33180),
            .I(N__33177));
    LocalMux I__6720 (
            .O(N__33177),
            .I(\nx.n3163 ));
    InMux I__6719 (
            .O(N__33174),
            .I(\nx.n11092 ));
    CascadeMux I__6718 (
            .O(N__33171),
            .I(N__33168));
    InMux I__6717 (
            .O(N__33168),
            .I(N__33165));
    LocalMux I__6716 (
            .O(N__33165),
            .I(N__33160));
    InMux I__6715 (
            .O(N__33164),
            .I(N__33157));
    InMux I__6714 (
            .O(N__33163),
            .I(N__33154));
    Span4Mux_h I__6713 (
            .O(N__33160),
            .I(N__33151));
    LocalMux I__6712 (
            .O(N__33157),
            .I(N__33148));
    LocalMux I__6711 (
            .O(N__33154),
            .I(\nx.n3095 ));
    Odrv4 I__6710 (
            .O(N__33151),
            .I(\nx.n3095 ));
    Odrv12 I__6709 (
            .O(N__33148),
            .I(\nx.n3095 ));
    InMux I__6708 (
            .O(N__33141),
            .I(N__33138));
    LocalMux I__6707 (
            .O(N__33138),
            .I(\nx.n3162 ));
    InMux I__6706 (
            .O(N__33135),
            .I(\nx.n11093 ));
    InMux I__6705 (
            .O(N__33132),
            .I(N__33128));
    InMux I__6704 (
            .O(N__33131),
            .I(N__33125));
    LocalMux I__6703 (
            .O(N__33128),
            .I(N__33121));
    LocalMux I__6702 (
            .O(N__33125),
            .I(N__33118));
    InMux I__6701 (
            .O(N__33124),
            .I(N__33115));
    Span4Mux_h I__6700 (
            .O(N__33121),
            .I(N__33110));
    Span4Mux_h I__6699 (
            .O(N__33118),
            .I(N__33110));
    LocalMux I__6698 (
            .O(N__33115),
            .I(\nx.n3094 ));
    Odrv4 I__6697 (
            .O(N__33110),
            .I(\nx.n3094 ));
    CascadeMux I__6696 (
            .O(N__33105),
            .I(N__33102));
    InMux I__6695 (
            .O(N__33102),
            .I(N__33099));
    LocalMux I__6694 (
            .O(N__33099),
            .I(\nx.n3161 ));
    InMux I__6693 (
            .O(N__33096),
            .I(bfn_13_19_0_));
    CascadeMux I__6692 (
            .O(N__33093),
            .I(N__33089));
    InMux I__6691 (
            .O(N__33092),
            .I(N__33086));
    InMux I__6690 (
            .O(N__33089),
            .I(N__33082));
    LocalMux I__6689 (
            .O(N__33086),
            .I(N__33079));
    InMux I__6688 (
            .O(N__33085),
            .I(N__33076));
    LocalMux I__6687 (
            .O(N__33082),
            .I(N__33073));
    Span4Mux_v I__6686 (
            .O(N__33079),
            .I(N__33070));
    LocalMux I__6685 (
            .O(N__33076),
            .I(N__33067));
    Span4Mux_v I__6684 (
            .O(N__33073),
            .I(N__33064));
    Span4Mux_h I__6683 (
            .O(N__33070),
            .I(N__33061));
    Odrv4 I__6682 (
            .O(N__33067),
            .I(\nx.n3093 ));
    Odrv4 I__6681 (
            .O(N__33064),
            .I(\nx.n3093 ));
    Odrv4 I__6680 (
            .O(N__33061),
            .I(\nx.n3093 ));
    CascadeMux I__6679 (
            .O(N__33054),
            .I(N__33051));
    InMux I__6678 (
            .O(N__33051),
            .I(N__33047));
    CascadeMux I__6677 (
            .O(N__33050),
            .I(N__33044));
    LocalMux I__6676 (
            .O(N__33047),
            .I(N__33040));
    InMux I__6675 (
            .O(N__33044),
            .I(N__33035));
    InMux I__6674 (
            .O(N__33043),
            .I(N__33035));
    Span4Mux_v I__6673 (
            .O(N__33040),
            .I(N__33032));
    LocalMux I__6672 (
            .O(N__33035),
            .I(\nx.n3108 ));
    Odrv4 I__6671 (
            .O(N__33032),
            .I(\nx.n3108 ));
    InMux I__6670 (
            .O(N__33027),
            .I(N__33024));
    LocalMux I__6669 (
            .O(N__33024),
            .I(N__33021));
    Span4Mux_h I__6668 (
            .O(N__33021),
            .I(N__33018));
    Odrv4 I__6667 (
            .O(N__33018),
            .I(\nx.n3175 ));
    InMux I__6666 (
            .O(N__33015),
            .I(\nx.n11080 ));
    CascadeMux I__6665 (
            .O(N__33012),
            .I(N__33009));
    InMux I__6664 (
            .O(N__33009),
            .I(N__33006));
    LocalMux I__6663 (
            .O(N__33006),
            .I(N__33001));
    InMux I__6662 (
            .O(N__33005),
            .I(N__32998));
    InMux I__6661 (
            .O(N__33004),
            .I(N__32995));
    Span4Mux_h I__6660 (
            .O(N__33001),
            .I(N__32992));
    LocalMux I__6659 (
            .O(N__32998),
            .I(\nx.n3107 ));
    LocalMux I__6658 (
            .O(N__32995),
            .I(\nx.n3107 ));
    Odrv4 I__6657 (
            .O(N__32992),
            .I(\nx.n3107 ));
    InMux I__6656 (
            .O(N__32985),
            .I(N__32982));
    LocalMux I__6655 (
            .O(N__32982),
            .I(\nx.n3174 ));
    InMux I__6654 (
            .O(N__32979),
            .I(\nx.n11081 ));
    CascadeMux I__6653 (
            .O(N__32976),
            .I(N__32972));
    InMux I__6652 (
            .O(N__32975),
            .I(N__32969));
    InMux I__6651 (
            .O(N__32972),
            .I(N__32966));
    LocalMux I__6650 (
            .O(N__32969),
            .I(N__32963));
    LocalMux I__6649 (
            .O(N__32966),
            .I(N__32959));
    Span4Mux_v I__6648 (
            .O(N__32963),
            .I(N__32956));
    InMux I__6647 (
            .O(N__32962),
            .I(N__32953));
    Span4Mux_h I__6646 (
            .O(N__32959),
            .I(N__32948));
    Span4Mux_h I__6645 (
            .O(N__32956),
            .I(N__32948));
    LocalMux I__6644 (
            .O(N__32953),
            .I(\nx.n3106 ));
    Odrv4 I__6643 (
            .O(N__32948),
            .I(\nx.n3106 ));
    InMux I__6642 (
            .O(N__32943),
            .I(N__32940));
    LocalMux I__6641 (
            .O(N__32940),
            .I(N__32937));
    Odrv4 I__6640 (
            .O(N__32937),
            .I(\nx.n3173 ));
    InMux I__6639 (
            .O(N__32934),
            .I(\nx.n11082 ));
    CascadeMux I__6638 (
            .O(N__32931),
            .I(N__32928));
    InMux I__6637 (
            .O(N__32928),
            .I(N__32925));
    LocalMux I__6636 (
            .O(N__32925),
            .I(N__32920));
    InMux I__6635 (
            .O(N__32924),
            .I(N__32917));
    InMux I__6634 (
            .O(N__32923),
            .I(N__32914));
    Span4Mux_h I__6633 (
            .O(N__32920),
            .I(N__32911));
    LocalMux I__6632 (
            .O(N__32917),
            .I(\nx.n3105 ));
    LocalMux I__6631 (
            .O(N__32914),
            .I(\nx.n3105 ));
    Odrv4 I__6630 (
            .O(N__32911),
            .I(\nx.n3105 ));
    InMux I__6629 (
            .O(N__32904),
            .I(N__32901));
    LocalMux I__6628 (
            .O(N__32901),
            .I(N__32898));
    Odrv4 I__6627 (
            .O(N__32898),
            .I(\nx.n3172 ));
    InMux I__6626 (
            .O(N__32895),
            .I(\nx.n11083 ));
    CascadeMux I__6625 (
            .O(N__32892),
            .I(N__32888));
    InMux I__6624 (
            .O(N__32891),
            .I(N__32885));
    InMux I__6623 (
            .O(N__32888),
            .I(N__32881));
    LocalMux I__6622 (
            .O(N__32885),
            .I(N__32878));
    InMux I__6621 (
            .O(N__32884),
            .I(N__32875));
    LocalMux I__6620 (
            .O(N__32881),
            .I(N__32872));
    Span4Mux_v I__6619 (
            .O(N__32878),
            .I(N__32869));
    LocalMux I__6618 (
            .O(N__32875),
            .I(N__32866));
    Span4Mux_h I__6617 (
            .O(N__32872),
            .I(N__32861));
    Span4Mux_h I__6616 (
            .O(N__32869),
            .I(N__32861));
    Odrv4 I__6615 (
            .O(N__32866),
            .I(\nx.n3104 ));
    Odrv4 I__6614 (
            .O(N__32861),
            .I(\nx.n3104 ));
    InMux I__6613 (
            .O(N__32856),
            .I(N__32853));
    LocalMux I__6612 (
            .O(N__32853),
            .I(\nx.n3171 ));
    InMux I__6611 (
            .O(N__32850),
            .I(\nx.n11084 ));
    CascadeMux I__6610 (
            .O(N__32847),
            .I(N__32844));
    InMux I__6609 (
            .O(N__32844),
            .I(N__32840));
    InMux I__6608 (
            .O(N__32843),
            .I(N__32837));
    LocalMux I__6607 (
            .O(N__32840),
            .I(N__32834));
    LocalMux I__6606 (
            .O(N__32837),
            .I(N__32830));
    Span4Mux_v I__6605 (
            .O(N__32834),
            .I(N__32827));
    InMux I__6604 (
            .O(N__32833),
            .I(N__32824));
    Span4Mux_h I__6603 (
            .O(N__32830),
            .I(N__32821));
    Span4Mux_h I__6602 (
            .O(N__32827),
            .I(N__32818));
    LocalMux I__6601 (
            .O(N__32824),
            .I(\nx.n3103 ));
    Odrv4 I__6600 (
            .O(N__32821),
            .I(\nx.n3103 ));
    Odrv4 I__6599 (
            .O(N__32818),
            .I(\nx.n3103 ));
    InMux I__6598 (
            .O(N__32811),
            .I(N__32808));
    LocalMux I__6597 (
            .O(N__32808),
            .I(\nx.n3170 ));
    InMux I__6596 (
            .O(N__32805),
            .I(\nx.n11085 ));
    CascadeMux I__6595 (
            .O(N__32802),
            .I(N__32799));
    InMux I__6594 (
            .O(N__32799),
            .I(N__32795));
    InMux I__6593 (
            .O(N__32798),
            .I(N__32791));
    LocalMux I__6592 (
            .O(N__32795),
            .I(N__32788));
    InMux I__6591 (
            .O(N__32794),
            .I(N__32785));
    LocalMux I__6590 (
            .O(N__32791),
            .I(\nx.n3102 ));
    Odrv4 I__6589 (
            .O(N__32788),
            .I(\nx.n3102 ));
    LocalMux I__6588 (
            .O(N__32785),
            .I(\nx.n3102 ));
    InMux I__6587 (
            .O(N__32778),
            .I(N__32775));
    LocalMux I__6586 (
            .O(N__32775),
            .I(\nx.n3169 ));
    InMux I__6585 (
            .O(N__32772),
            .I(bfn_13_18_0_));
    CascadeMux I__6584 (
            .O(N__32769),
            .I(N__32764));
    CascadeMux I__6583 (
            .O(N__32768),
            .I(N__32761));
    CascadeMux I__6582 (
            .O(N__32767),
            .I(N__32758));
    InMux I__6581 (
            .O(N__32764),
            .I(N__32755));
    InMux I__6580 (
            .O(N__32761),
            .I(N__32752));
    InMux I__6579 (
            .O(N__32758),
            .I(N__32749));
    LocalMux I__6578 (
            .O(N__32755),
            .I(N__32746));
    LocalMux I__6577 (
            .O(N__32752),
            .I(N__32743));
    LocalMux I__6576 (
            .O(N__32749),
            .I(N__32740));
    Span4Mux_h I__6575 (
            .O(N__32746),
            .I(N__32737));
    Span4Mux_v I__6574 (
            .O(N__32743),
            .I(N__32732));
    Span4Mux_h I__6573 (
            .O(N__32740),
            .I(N__32732));
    Odrv4 I__6572 (
            .O(N__32737),
            .I(\nx.n3101 ));
    Odrv4 I__6571 (
            .O(N__32732),
            .I(\nx.n3101 ));
    InMux I__6570 (
            .O(N__32727),
            .I(N__32724));
    LocalMux I__6569 (
            .O(N__32724),
            .I(\nx.n3168 ));
    InMux I__6568 (
            .O(N__32721),
            .I(\nx.n11087 ));
    InMux I__6567 (
            .O(N__32718),
            .I(N__32715));
    LocalMux I__6566 (
            .O(N__32715),
            .I(N__32712));
    Odrv4 I__6565 (
            .O(N__32712),
            .I(\nx.n2169 ));
    CascadeMux I__6564 (
            .O(N__32709),
            .I(N__32704));
    CascadeMux I__6563 (
            .O(N__32708),
            .I(N__32701));
    CascadeMux I__6562 (
            .O(N__32707),
            .I(N__32698));
    InMux I__6561 (
            .O(N__32704),
            .I(N__32695));
    InMux I__6560 (
            .O(N__32701),
            .I(N__32692));
    InMux I__6559 (
            .O(N__32698),
            .I(N__32689));
    LocalMux I__6558 (
            .O(N__32695),
            .I(N__32684));
    LocalMux I__6557 (
            .O(N__32692),
            .I(N__32684));
    LocalMux I__6556 (
            .O(N__32689),
            .I(N__32681));
    Span4Mux_v I__6555 (
            .O(N__32684),
            .I(N__32678));
    Odrv12 I__6554 (
            .O(N__32681),
            .I(\nx.n2102 ));
    Odrv4 I__6553 (
            .O(N__32678),
            .I(\nx.n2102 ));
    CascadeMux I__6552 (
            .O(N__32673),
            .I(N__32670));
    InMux I__6551 (
            .O(N__32670),
            .I(N__32666));
    InMux I__6550 (
            .O(N__32669),
            .I(N__32662));
    LocalMux I__6549 (
            .O(N__32666),
            .I(N__32659));
    InMux I__6548 (
            .O(N__32665),
            .I(N__32656));
    LocalMux I__6547 (
            .O(N__32662),
            .I(\nx.n2201 ));
    Odrv4 I__6546 (
            .O(N__32659),
            .I(\nx.n2201 ));
    LocalMux I__6545 (
            .O(N__32656),
            .I(\nx.n2201 ));
    InMux I__6544 (
            .O(N__32649),
            .I(N__32646));
    LocalMux I__6543 (
            .O(N__32646),
            .I(\nx.n2261 ));
    CascadeMux I__6542 (
            .O(N__32643),
            .I(N__32639));
    InMux I__6541 (
            .O(N__32642),
            .I(N__32635));
    InMux I__6540 (
            .O(N__32639),
            .I(N__32632));
    InMux I__6539 (
            .O(N__32638),
            .I(N__32629));
    LocalMux I__6538 (
            .O(N__32635),
            .I(\nx.n2194 ));
    LocalMux I__6537 (
            .O(N__32632),
            .I(\nx.n2194 ));
    LocalMux I__6536 (
            .O(N__32629),
            .I(\nx.n2194 ));
    InMux I__6535 (
            .O(N__32622),
            .I(N__32619));
    LocalMux I__6534 (
            .O(N__32619),
            .I(N__32616));
    Odrv4 I__6533 (
            .O(N__32616),
            .I(\nx.n2262 ));
    CascadeMux I__6532 (
            .O(N__32613),
            .I(N__32610));
    InMux I__6531 (
            .O(N__32610),
            .I(N__32606));
    CascadeMux I__6530 (
            .O(N__32609),
            .I(N__32603));
    LocalMux I__6529 (
            .O(N__32606),
            .I(N__32600));
    InMux I__6528 (
            .O(N__32603),
            .I(N__32597));
    Span4Mux_v I__6527 (
            .O(N__32600),
            .I(N__32593));
    LocalMux I__6526 (
            .O(N__32597),
            .I(N__32590));
    InMux I__6525 (
            .O(N__32596),
            .I(N__32587));
    Odrv4 I__6524 (
            .O(N__32593),
            .I(\nx.n2195 ));
    Odrv4 I__6523 (
            .O(N__32590),
            .I(\nx.n2195 ));
    LocalMux I__6522 (
            .O(N__32587),
            .I(\nx.n2195 ));
    CascadeMux I__6521 (
            .O(N__32580),
            .I(N__32573));
    InMux I__6520 (
            .O(N__32579),
            .I(N__32566));
    CascadeMux I__6519 (
            .O(N__32578),
            .I(N__32563));
    CascadeMux I__6518 (
            .O(N__32577),
            .I(N__32555));
    CascadeMux I__6517 (
            .O(N__32576),
            .I(N__32549));
    InMux I__6516 (
            .O(N__32573),
            .I(N__32542));
    InMux I__6515 (
            .O(N__32572),
            .I(N__32542));
    InMux I__6514 (
            .O(N__32571),
            .I(N__32542));
    CascadeMux I__6513 (
            .O(N__32570),
            .I(N__32539));
    CascadeMux I__6512 (
            .O(N__32569),
            .I(N__32535));
    LocalMux I__6511 (
            .O(N__32566),
            .I(N__32532));
    InMux I__6510 (
            .O(N__32563),
            .I(N__32525));
    InMux I__6509 (
            .O(N__32562),
            .I(N__32525));
    InMux I__6508 (
            .O(N__32561),
            .I(N__32525));
    InMux I__6507 (
            .O(N__32560),
            .I(N__32518));
    InMux I__6506 (
            .O(N__32559),
            .I(N__32518));
    InMux I__6505 (
            .O(N__32558),
            .I(N__32518));
    InMux I__6504 (
            .O(N__32555),
            .I(N__32511));
    InMux I__6503 (
            .O(N__32554),
            .I(N__32511));
    InMux I__6502 (
            .O(N__32553),
            .I(N__32511));
    InMux I__6501 (
            .O(N__32552),
            .I(N__32506));
    InMux I__6500 (
            .O(N__32549),
            .I(N__32506));
    LocalMux I__6499 (
            .O(N__32542),
            .I(N__32503));
    InMux I__6498 (
            .O(N__32539),
            .I(N__32496));
    InMux I__6497 (
            .O(N__32538),
            .I(N__32496));
    InMux I__6496 (
            .O(N__32535),
            .I(N__32496));
    Span4Mux_h I__6495 (
            .O(N__32532),
            .I(N__32493));
    LocalMux I__6494 (
            .O(N__32525),
            .I(N__32490));
    LocalMux I__6493 (
            .O(N__32518),
            .I(\nx.n2225 ));
    LocalMux I__6492 (
            .O(N__32511),
            .I(\nx.n2225 ));
    LocalMux I__6491 (
            .O(N__32506),
            .I(\nx.n2225 ));
    Odrv4 I__6490 (
            .O(N__32503),
            .I(\nx.n2225 ));
    LocalMux I__6489 (
            .O(N__32496),
            .I(\nx.n2225 ));
    Odrv4 I__6488 (
            .O(N__32493),
            .I(\nx.n2225 ));
    Odrv12 I__6487 (
            .O(N__32490),
            .I(\nx.n2225 ));
    IoInMux I__6486 (
            .O(N__32475),
            .I(N__32472));
    LocalMux I__6485 (
            .O(N__32472),
            .I(N__32469));
    IoSpan4Mux I__6484 (
            .O(N__32469),
            .I(N__32466));
    Sp12to4 I__6483 (
            .O(N__32466),
            .I(N__32463));
    Span12Mux_h I__6482 (
            .O(N__32463),
            .I(N__32459));
    InMux I__6481 (
            .O(N__32462),
            .I(N__32456));
    Odrv12 I__6480 (
            .O(N__32459),
            .I(pin_oe_4));
    LocalMux I__6479 (
            .O(N__32456),
            .I(pin_oe_4));
    CascadeMux I__6478 (
            .O(N__32451),
            .I(n11970_cascade_));
    IoInMux I__6477 (
            .O(N__32448),
            .I(N__32445));
    LocalMux I__6476 (
            .O(N__32445),
            .I(N__32442));
    Span12Mux_s4_v I__6475 (
            .O(N__32442),
            .I(N__32439));
    Span12Mux_h I__6474 (
            .O(N__32439),
            .I(N__32436));
    Span12Mux_v I__6473 (
            .O(N__32436),
            .I(N__32432));
    InMux I__6472 (
            .O(N__32435),
            .I(N__32429));
    Odrv12 I__6471 (
            .O(N__32432),
            .I(pin_oe_0));
    LocalMux I__6470 (
            .O(N__32429),
            .I(pin_oe_0));
    InMux I__6469 (
            .O(N__32424),
            .I(N__32421));
    LocalMux I__6468 (
            .O(N__32421),
            .I(N__32418));
    Span4Mux_h I__6467 (
            .O(N__32418),
            .I(N__32415));
    Odrv4 I__6466 (
            .O(N__32415),
            .I(n11968));
    InMux I__6465 (
            .O(N__32412),
            .I(N__32408));
    InMux I__6464 (
            .O(N__32411),
            .I(N__32405));
    LocalMux I__6463 (
            .O(N__32408),
            .I(N__32400));
    LocalMux I__6462 (
            .O(N__32405),
            .I(N__32400));
    Span4Mux_h I__6461 (
            .O(N__32400),
            .I(N__32396));
    InMux I__6460 (
            .O(N__32399),
            .I(N__32393));
    Sp12to4 I__6459 (
            .O(N__32396),
            .I(N__32386));
    LocalMux I__6458 (
            .O(N__32393),
            .I(N__32386));
    InMux I__6457 (
            .O(N__32392),
            .I(N__32383));
    InMux I__6456 (
            .O(N__32391),
            .I(N__32380));
    Span12Mux_v I__6455 (
            .O(N__32386),
            .I(N__32377));
    LocalMux I__6454 (
            .O(N__32383),
            .I(\nx.bit_ctr_4 ));
    LocalMux I__6453 (
            .O(N__32380),
            .I(\nx.bit_ctr_4 ));
    Odrv12 I__6452 (
            .O(N__32377),
            .I(\nx.bit_ctr_4 ));
    InMux I__6451 (
            .O(N__32370),
            .I(N__32367));
    LocalMux I__6450 (
            .O(N__32367),
            .I(N__32364));
    Odrv4 I__6449 (
            .O(N__32364),
            .I(\nx.n3177 ));
    InMux I__6448 (
            .O(N__32361),
            .I(bfn_13_17_0_));
    CascadeMux I__6447 (
            .O(N__32358),
            .I(N__32355));
    InMux I__6446 (
            .O(N__32355),
            .I(N__32350));
    CascadeMux I__6445 (
            .O(N__32354),
            .I(N__32347));
    CascadeMux I__6444 (
            .O(N__32353),
            .I(N__32344));
    LocalMux I__6443 (
            .O(N__32350),
            .I(N__32341));
    InMux I__6442 (
            .O(N__32347),
            .I(N__32338));
    InMux I__6441 (
            .O(N__32344),
            .I(N__32335));
    Span4Mux_v I__6440 (
            .O(N__32341),
            .I(N__32332));
    LocalMux I__6439 (
            .O(N__32338),
            .I(\nx.n3109 ));
    LocalMux I__6438 (
            .O(N__32335),
            .I(\nx.n3109 ));
    Odrv4 I__6437 (
            .O(N__32332),
            .I(\nx.n3109 ));
    InMux I__6436 (
            .O(N__32325),
            .I(N__32322));
    LocalMux I__6435 (
            .O(N__32322),
            .I(\nx.n3176 ));
    InMux I__6434 (
            .O(N__32319),
            .I(\nx.n11079 ));
    CascadeMux I__6433 (
            .O(N__32316),
            .I(\nx.n2299_cascade_ ));
    CascadeMux I__6432 (
            .O(N__32313),
            .I(N__32310));
    InMux I__6431 (
            .O(N__32310),
            .I(N__32307));
    LocalMux I__6430 (
            .O(N__32307),
            .I(\nx.n2265 ));
    CascadeMux I__6429 (
            .O(N__32304),
            .I(N__32301));
    InMux I__6428 (
            .O(N__32301),
            .I(N__32298));
    LocalMux I__6427 (
            .O(N__32298),
            .I(N__32294));
    CascadeMux I__6426 (
            .O(N__32297),
            .I(N__32291));
    Span4Mux_h I__6425 (
            .O(N__32294),
            .I(N__32287));
    InMux I__6424 (
            .O(N__32291),
            .I(N__32284));
    InMux I__6423 (
            .O(N__32290),
            .I(N__32281));
    Odrv4 I__6422 (
            .O(N__32287),
            .I(\nx.n2197 ));
    LocalMux I__6421 (
            .O(N__32284),
            .I(\nx.n2197 ));
    LocalMux I__6420 (
            .O(N__32281),
            .I(\nx.n2197 ));
    CascadeMux I__6419 (
            .O(N__32274),
            .I(N__32271));
    InMux I__6418 (
            .O(N__32271),
            .I(N__32267));
    InMux I__6417 (
            .O(N__32270),
            .I(N__32264));
    LocalMux I__6416 (
            .O(N__32267),
            .I(\nx.n2196 ));
    LocalMux I__6415 (
            .O(N__32264),
            .I(\nx.n2196 ));
    InMux I__6414 (
            .O(N__32259),
            .I(N__32256));
    LocalMux I__6413 (
            .O(N__32256),
            .I(\nx.n30_adj_694 ));
    InMux I__6412 (
            .O(N__32253),
            .I(N__32250));
    LocalMux I__6411 (
            .O(N__32250),
            .I(N__32247));
    Span4Mux_h I__6410 (
            .O(N__32247),
            .I(N__32244));
    Odrv4 I__6409 (
            .O(N__32244),
            .I(\nx.n22_adj_693 ));
    CascadeMux I__6408 (
            .O(N__32241),
            .I(\nx.n21_cascade_ ));
    InMux I__6407 (
            .O(N__32238),
            .I(N__32235));
    LocalMux I__6406 (
            .O(N__32235),
            .I(\nx.n34_adj_695 ));
    InMux I__6405 (
            .O(N__32232),
            .I(N__32229));
    LocalMux I__6404 (
            .O(N__32229),
            .I(\nx.n2268 ));
    CascadeMux I__6403 (
            .O(N__32226),
            .I(\nx.n2225_cascade_ ));
    InMux I__6402 (
            .O(N__32223),
            .I(N__32215));
    InMux I__6401 (
            .O(N__32222),
            .I(N__32215));
    InMux I__6400 (
            .O(N__32221),
            .I(N__32212));
    InMux I__6399 (
            .O(N__32220),
            .I(N__32209));
    LocalMux I__6398 (
            .O(N__32215),
            .I(N__32204));
    LocalMux I__6397 (
            .O(N__32212),
            .I(N__32204));
    LocalMux I__6396 (
            .O(N__32209),
            .I(N__32200));
    Sp12to4 I__6395 (
            .O(N__32204),
            .I(N__32197));
    InMux I__6394 (
            .O(N__32203),
            .I(N__32194));
    Span12Mux_s11_h I__6393 (
            .O(N__32200),
            .I(N__32191));
    Span12Mux_v I__6392 (
            .O(N__32197),
            .I(N__32188));
    LocalMux I__6391 (
            .O(N__32194),
            .I(neopxl_color_4));
    Odrv12 I__6390 (
            .O(N__32191),
            .I(neopxl_color_4));
    Odrv12 I__6389 (
            .O(N__32188),
            .I(neopxl_color_4));
    SRMux I__6388 (
            .O(N__32181),
            .I(N__32178));
    LocalMux I__6387 (
            .O(N__32178),
            .I(N__32175));
    Span4Mux_h I__6386 (
            .O(N__32175),
            .I(N__32172));
    Span4Mux_v I__6385 (
            .O(N__32172),
            .I(N__32169));
    Odrv4 I__6384 (
            .O(N__32169),
            .I(n22_adj_787));
    CascadeMux I__6383 (
            .O(N__32166),
            .I(N__32163));
    InMux I__6382 (
            .O(N__32163),
            .I(N__32159));
    InMux I__6381 (
            .O(N__32162),
            .I(N__32156));
    LocalMux I__6380 (
            .O(N__32159),
            .I(N__32153));
    LocalMux I__6379 (
            .O(N__32156),
            .I(N__32150));
    Span4Mux_h I__6378 (
            .O(N__32153),
            .I(N__32147));
    Odrv12 I__6377 (
            .O(N__32150),
            .I(\nx.n2099 ));
    Odrv4 I__6376 (
            .O(N__32147),
            .I(\nx.n2099 ));
    InMux I__6375 (
            .O(N__32142),
            .I(N__32139));
    LocalMux I__6374 (
            .O(N__32139),
            .I(N__32136));
    Odrv4 I__6373 (
            .O(N__32136),
            .I(\nx.n2166 ));
    InMux I__6372 (
            .O(N__32133),
            .I(N__32129));
    InMux I__6371 (
            .O(N__32132),
            .I(N__32125));
    LocalMux I__6370 (
            .O(N__32129),
            .I(N__32122));
    InMux I__6369 (
            .O(N__32128),
            .I(N__32119));
    LocalMux I__6368 (
            .O(N__32125),
            .I(\nx.n2198 ));
    Odrv4 I__6367 (
            .O(N__32122),
            .I(\nx.n2198 ));
    LocalMux I__6366 (
            .O(N__32119),
            .I(\nx.n2198 ));
    InMux I__6365 (
            .O(N__32112),
            .I(N__32109));
    LocalMux I__6364 (
            .O(N__32109),
            .I(\nx.n2274 ));
    CascadeMux I__6363 (
            .O(N__32106),
            .I(N__32102));
    InMux I__6362 (
            .O(N__32105),
            .I(N__32099));
    InMux I__6361 (
            .O(N__32102),
            .I(N__32096));
    LocalMux I__6360 (
            .O(N__32099),
            .I(N__32093));
    LocalMux I__6359 (
            .O(N__32096),
            .I(N__32089));
    Span4Mux_v I__6358 (
            .O(N__32093),
            .I(N__32086));
    InMux I__6357 (
            .O(N__32092),
            .I(N__32083));
    Span4Mux_h I__6356 (
            .O(N__32089),
            .I(N__32080));
    Odrv4 I__6355 (
            .O(N__32086),
            .I(\nx.n2207 ));
    LocalMux I__6354 (
            .O(N__32083),
            .I(\nx.n2207 ));
    Odrv4 I__6353 (
            .O(N__32080),
            .I(\nx.n2207 ));
    InMux I__6352 (
            .O(N__32073),
            .I(N__32069));
    CascadeMux I__6351 (
            .O(N__32072),
            .I(N__32066));
    LocalMux I__6350 (
            .O(N__32069),
            .I(N__32063));
    InMux I__6349 (
            .O(N__32066),
            .I(N__32059));
    Span4Mux_h I__6348 (
            .O(N__32063),
            .I(N__32056));
    InMux I__6347 (
            .O(N__32062),
            .I(N__32053));
    LocalMux I__6346 (
            .O(N__32059),
            .I(N__32050));
    Odrv4 I__6345 (
            .O(N__32056),
            .I(\nx.n2208 ));
    LocalMux I__6344 (
            .O(N__32053),
            .I(\nx.n2208 ));
    Odrv4 I__6343 (
            .O(N__32050),
            .I(\nx.n2208 ));
    CascadeMux I__6342 (
            .O(N__32043),
            .I(N__32040));
    InMux I__6341 (
            .O(N__32040),
            .I(N__32037));
    LocalMux I__6340 (
            .O(N__32037),
            .I(N__32034));
    Odrv4 I__6339 (
            .O(N__32034),
            .I(\nx.n2275 ));
    InMux I__6338 (
            .O(N__32031),
            .I(N__32028));
    LocalMux I__6337 (
            .O(N__32028),
            .I(\nx.n2272 ));
    CascadeMux I__6336 (
            .O(N__32025),
            .I(N__32021));
    InMux I__6335 (
            .O(N__32024),
            .I(N__32018));
    InMux I__6334 (
            .O(N__32021),
            .I(N__32015));
    LocalMux I__6333 (
            .O(N__32018),
            .I(N__32012));
    LocalMux I__6332 (
            .O(N__32015),
            .I(N__32008));
    Span4Mux_h I__6331 (
            .O(N__32012),
            .I(N__32005));
    InMux I__6330 (
            .O(N__32011),
            .I(N__32002));
    Span4Mux_v I__6329 (
            .O(N__32008),
            .I(N__31999));
    Odrv4 I__6328 (
            .O(N__32005),
            .I(\nx.n2205 ));
    LocalMux I__6327 (
            .O(N__32002),
            .I(\nx.n2205 ));
    Odrv4 I__6326 (
            .O(N__31999),
            .I(\nx.n2205 ));
    CascadeMux I__6325 (
            .O(N__31992),
            .I(\nx.n2391_cascade_ ));
    CascadeMux I__6324 (
            .O(N__31989),
            .I(\nx.n30_adj_696_cascade_ ));
    InMux I__6323 (
            .O(N__31986),
            .I(N__31983));
    LocalMux I__6322 (
            .O(N__31983),
            .I(\nx.n2266 ));
    CascadeMux I__6321 (
            .O(N__31980),
            .I(N__31976));
    InMux I__6320 (
            .O(N__31979),
            .I(N__31973));
    InMux I__6319 (
            .O(N__31976),
            .I(N__31970));
    LocalMux I__6318 (
            .O(N__31973),
            .I(N__31967));
    LocalMux I__6317 (
            .O(N__31970),
            .I(\nx.n2199 ));
    Odrv4 I__6316 (
            .O(N__31967),
            .I(\nx.n2199 ));
    InMux I__6315 (
            .O(N__31962),
            .I(N__31959));
    LocalMux I__6314 (
            .O(N__31959),
            .I(\nx.n2267 ));
    InMux I__6313 (
            .O(N__31956),
            .I(N__31952));
    CascadeMux I__6312 (
            .O(N__31955),
            .I(N__31948));
    LocalMux I__6311 (
            .O(N__31952),
            .I(N__31945));
    CascadeMux I__6310 (
            .O(N__31951),
            .I(N__31942));
    InMux I__6309 (
            .O(N__31948),
            .I(N__31939));
    Span4Mux_h I__6308 (
            .O(N__31945),
            .I(N__31936));
    InMux I__6307 (
            .O(N__31942),
            .I(N__31933));
    LocalMux I__6306 (
            .O(N__31939),
            .I(N__31930));
    Odrv4 I__6305 (
            .O(N__31936),
            .I(\nx.n2204 ));
    LocalMux I__6304 (
            .O(N__31933),
            .I(\nx.n2204 ));
    Odrv4 I__6303 (
            .O(N__31930),
            .I(\nx.n2204 ));
    CascadeMux I__6302 (
            .O(N__31923),
            .I(N__31920));
    InMux I__6301 (
            .O(N__31920),
            .I(N__31917));
    LocalMux I__6300 (
            .O(N__31917),
            .I(\nx.n2271 ));
    CascadeMux I__6299 (
            .O(N__31914),
            .I(\nx.n2303_cascade_ ));
    InMux I__6298 (
            .O(N__31911),
            .I(N__31908));
    LocalMux I__6297 (
            .O(N__31908),
            .I(\nx.n2269 ));
    InMux I__6296 (
            .O(N__31905),
            .I(N__31901));
    CascadeMux I__6295 (
            .O(N__31904),
            .I(N__31898));
    LocalMux I__6294 (
            .O(N__31901),
            .I(N__31895));
    InMux I__6293 (
            .O(N__31898),
            .I(N__31892));
    Span4Mux_h I__6292 (
            .O(N__31895),
            .I(N__31887));
    LocalMux I__6291 (
            .O(N__31892),
            .I(N__31887));
    Odrv4 I__6290 (
            .O(N__31887),
            .I(\nx.n2202 ));
    InMux I__6289 (
            .O(N__31884),
            .I(N__31880));
    CascadeMux I__6288 (
            .O(N__31883),
            .I(N__31877));
    LocalMux I__6287 (
            .O(N__31880),
            .I(N__31874));
    InMux I__6286 (
            .O(N__31877),
            .I(N__31870));
    Span4Mux_v I__6285 (
            .O(N__31874),
            .I(N__31867));
    InMux I__6284 (
            .O(N__31873),
            .I(N__31864));
    LocalMux I__6283 (
            .O(N__31870),
            .I(N__31861));
    Odrv4 I__6282 (
            .O(N__31867),
            .I(\nx.n2203 ));
    LocalMux I__6281 (
            .O(N__31864),
            .I(\nx.n2203 ));
    Odrv12 I__6280 (
            .O(N__31861),
            .I(\nx.n2203 ));
    CascadeMux I__6279 (
            .O(N__31854),
            .I(N__31851));
    InMux I__6278 (
            .O(N__31851),
            .I(N__31848));
    LocalMux I__6277 (
            .O(N__31848),
            .I(\nx.n2270 ));
    CascadeMux I__6276 (
            .O(N__31845),
            .I(\nx.n2302_cascade_ ));
    CascadeMux I__6275 (
            .O(N__31842),
            .I(\nx.n2401_cascade_ ));
    InMux I__6274 (
            .O(N__31839),
            .I(N__31836));
    LocalMux I__6273 (
            .O(N__31836),
            .I(N__31833));
    Odrv4 I__6272 (
            .O(N__31833),
            .I(\nx.n38 ));
    InMux I__6271 (
            .O(N__31830),
            .I(N__31827));
    LocalMux I__6270 (
            .O(N__31827),
            .I(\nx.n37 ));
    CascadeMux I__6269 (
            .O(N__31824),
            .I(\nx.n39_cascade_ ));
    CascadeMux I__6268 (
            .O(N__31821),
            .I(\nx.n2621_cascade_ ));
    CascadeMux I__6267 (
            .O(N__31818),
            .I(N__31815));
    InMux I__6266 (
            .O(N__31815),
            .I(N__31810));
    InMux I__6265 (
            .O(N__31814),
            .I(N__31807));
    InMux I__6264 (
            .O(N__31813),
            .I(N__31804));
    LocalMux I__6263 (
            .O(N__31810),
            .I(N__31801));
    LocalMux I__6262 (
            .O(N__31807),
            .I(\nx.n2707 ));
    LocalMux I__6261 (
            .O(N__31804),
            .I(\nx.n2707 ));
    Odrv4 I__6260 (
            .O(N__31801),
            .I(\nx.n2707 ));
    InMux I__6259 (
            .O(N__31794),
            .I(N__31791));
    LocalMux I__6258 (
            .O(N__31791),
            .I(N__31786));
    InMux I__6257 (
            .O(N__31790),
            .I(N__31783));
    InMux I__6256 (
            .O(N__31789),
            .I(N__31780));
    Span4Mux_v I__6255 (
            .O(N__31786),
            .I(N__31775));
    LocalMux I__6254 (
            .O(N__31783),
            .I(N__31772));
    LocalMux I__6253 (
            .O(N__31780),
            .I(N__31769));
    InMux I__6252 (
            .O(N__31779),
            .I(N__31766));
    InMux I__6251 (
            .O(N__31778),
            .I(N__31763));
    Span4Mux_h I__6250 (
            .O(N__31775),
            .I(N__31760));
    Span4Mux_h I__6249 (
            .O(N__31772),
            .I(N__31755));
    Span4Mux_v I__6248 (
            .O(N__31769),
            .I(N__31755));
    LocalMux I__6247 (
            .O(N__31766),
            .I(\nx.bit_ctr_13 ));
    LocalMux I__6246 (
            .O(N__31763),
            .I(\nx.bit_ctr_13 ));
    Odrv4 I__6245 (
            .O(N__31760),
            .I(\nx.bit_ctr_13 ));
    Odrv4 I__6244 (
            .O(N__31755),
            .I(\nx.bit_ctr_13 ));
    InMux I__6243 (
            .O(N__31746),
            .I(N__31743));
    LocalMux I__6242 (
            .O(N__31743),
            .I(\nx.n2277 ));
    CascadeMux I__6241 (
            .O(N__31740),
            .I(\nx.n2309_cascade_ ));
    CascadeMux I__6240 (
            .O(N__31737),
            .I(\nx.n9697_cascade_ ));
    InMux I__6239 (
            .O(N__31734),
            .I(N__31731));
    LocalMux I__6238 (
            .O(N__31731),
            .I(\nx.n2273 ));
    InMux I__6237 (
            .O(N__31728),
            .I(N__31725));
    LocalMux I__6236 (
            .O(N__31725),
            .I(N__31720));
    InMux I__6235 (
            .O(N__31724),
            .I(N__31717));
    InMux I__6234 (
            .O(N__31723),
            .I(N__31714));
    Span4Mux_h I__6233 (
            .O(N__31720),
            .I(N__31709));
    LocalMux I__6232 (
            .O(N__31717),
            .I(N__31709));
    LocalMux I__6231 (
            .O(N__31714),
            .I(\nx.n2206 ));
    Odrv4 I__6230 (
            .O(N__31709),
            .I(\nx.n2206 ));
    InMux I__6229 (
            .O(N__31704),
            .I(N__31700));
    CascadeMux I__6228 (
            .O(N__31703),
            .I(N__31697));
    LocalMux I__6227 (
            .O(N__31700),
            .I(N__31693));
    InMux I__6226 (
            .O(N__31697),
            .I(N__31690));
    InMux I__6225 (
            .O(N__31696),
            .I(N__31687));
    Span4Mux_h I__6224 (
            .O(N__31693),
            .I(N__31682));
    LocalMux I__6223 (
            .O(N__31690),
            .I(N__31682));
    LocalMux I__6222 (
            .O(N__31687),
            .I(\nx.n2209 ));
    Odrv4 I__6221 (
            .O(N__31682),
            .I(\nx.n2209 ));
    CascadeMux I__6220 (
            .O(N__31677),
            .I(N__31674));
    InMux I__6219 (
            .O(N__31674),
            .I(N__31671));
    LocalMux I__6218 (
            .O(N__31671),
            .I(\nx.n2276 ));
    CascadeMux I__6217 (
            .O(N__31668),
            .I(N__31664));
    InMux I__6216 (
            .O(N__31667),
            .I(N__31661));
    InMux I__6215 (
            .O(N__31664),
            .I(N__31658));
    LocalMux I__6214 (
            .O(N__31661),
            .I(N__31654));
    LocalMux I__6213 (
            .O(N__31658),
            .I(N__31651));
    InMux I__6212 (
            .O(N__31657),
            .I(N__31648));
    Odrv4 I__6211 (
            .O(N__31654),
            .I(\nx.n2695 ));
    Odrv4 I__6210 (
            .O(N__31651),
            .I(\nx.n2695 ));
    LocalMux I__6209 (
            .O(N__31648),
            .I(\nx.n2695 ));
    CascadeMux I__6208 (
            .O(N__31641),
            .I(\nx.n2597_cascade_ ));
    CascadeMux I__6207 (
            .O(N__31638),
            .I(N__31634));
    InMux I__6206 (
            .O(N__31637),
            .I(N__31631));
    InMux I__6205 (
            .O(N__31634),
            .I(N__31628));
    LocalMux I__6204 (
            .O(N__31631),
            .I(N__31625));
    LocalMux I__6203 (
            .O(N__31628),
            .I(N__31622));
    Span4Mux_v I__6202 (
            .O(N__31625),
            .I(N__31619));
    Span4Mux_h I__6201 (
            .O(N__31622),
            .I(N__31616));
    Odrv4 I__6200 (
            .O(N__31619),
            .I(\nx.n2691 ));
    Odrv4 I__6199 (
            .O(N__31616),
            .I(\nx.n2691 ));
    CascadeMux I__6198 (
            .O(N__31611),
            .I(N__31608));
    InMux I__6197 (
            .O(N__31608),
            .I(N__31604));
    CascadeMux I__6196 (
            .O(N__31607),
            .I(N__31601));
    LocalMux I__6195 (
            .O(N__31604),
            .I(N__31598));
    InMux I__6194 (
            .O(N__31601),
            .I(N__31595));
    Span4Mux_v I__6193 (
            .O(N__31598),
            .I(N__31591));
    LocalMux I__6192 (
            .O(N__31595),
            .I(N__31588));
    InMux I__6191 (
            .O(N__31594),
            .I(N__31585));
    Odrv4 I__6190 (
            .O(N__31591),
            .I(\nx.n2690 ));
    Odrv4 I__6189 (
            .O(N__31588),
            .I(\nx.n2690 ));
    LocalMux I__6188 (
            .O(N__31585),
            .I(\nx.n2690 ));
    CascadeMux I__6187 (
            .O(N__31578),
            .I(\nx.n2691_cascade_ ));
    CascadeMux I__6186 (
            .O(N__31575),
            .I(N__31571));
    InMux I__6185 (
            .O(N__31574),
            .I(N__31568));
    InMux I__6184 (
            .O(N__31571),
            .I(N__31565));
    LocalMux I__6183 (
            .O(N__31568),
            .I(N__31562));
    LocalMux I__6182 (
            .O(N__31565),
            .I(N__31559));
    Span4Mux_v I__6181 (
            .O(N__31562),
            .I(N__31555));
    Span4Mux_v I__6180 (
            .O(N__31559),
            .I(N__31552));
    InMux I__6179 (
            .O(N__31558),
            .I(N__31549));
    Odrv4 I__6178 (
            .O(N__31555),
            .I(\nx.n2692 ));
    Odrv4 I__6177 (
            .O(N__31552),
            .I(\nx.n2692 ));
    LocalMux I__6176 (
            .O(N__31549),
            .I(\nx.n2692 ));
    InMux I__6175 (
            .O(N__31542),
            .I(N__31539));
    LocalMux I__6174 (
            .O(N__31539),
            .I(\nx.n36 ));
    CascadeMux I__6173 (
            .O(N__31536),
            .I(N__31533));
    InMux I__6172 (
            .O(N__31533),
            .I(N__31530));
    LocalMux I__6171 (
            .O(N__31530),
            .I(N__31525));
    InMux I__6170 (
            .O(N__31529),
            .I(N__31522));
    InMux I__6169 (
            .O(N__31528),
            .I(N__31519));
    Span4Mux_h I__6168 (
            .O(N__31525),
            .I(N__31516));
    LocalMux I__6167 (
            .O(N__31522),
            .I(\nx.n2700 ));
    LocalMux I__6166 (
            .O(N__31519),
            .I(\nx.n2700 ));
    Odrv4 I__6165 (
            .O(N__31516),
            .I(\nx.n2700 ));
    CascadeMux I__6164 (
            .O(N__31509),
            .I(N__31506));
    InMux I__6163 (
            .O(N__31506),
            .I(N__31502));
    CascadeMux I__6162 (
            .O(N__31505),
            .I(N__31499));
    LocalMux I__6161 (
            .O(N__31502),
            .I(N__31496));
    InMux I__6160 (
            .O(N__31499),
            .I(N__31492));
    Span4Mux_h I__6159 (
            .O(N__31496),
            .I(N__31489));
    InMux I__6158 (
            .O(N__31495),
            .I(N__31486));
    LocalMux I__6157 (
            .O(N__31492),
            .I(\nx.n2688 ));
    Odrv4 I__6156 (
            .O(N__31489),
            .I(\nx.n2688 ));
    LocalMux I__6155 (
            .O(N__31486),
            .I(\nx.n2688 ));
    CascadeMux I__6154 (
            .O(N__31479),
            .I(N__31475));
    CascadeMux I__6153 (
            .O(N__31478),
            .I(N__31472));
    InMux I__6152 (
            .O(N__31475),
            .I(N__31469));
    InMux I__6151 (
            .O(N__31472),
            .I(N__31466));
    LocalMux I__6150 (
            .O(N__31469),
            .I(N__31463));
    LocalMux I__6149 (
            .O(N__31466),
            .I(N__31460));
    Span4Mux_v I__6148 (
            .O(N__31463),
            .I(N__31456));
    Span4Mux_h I__6147 (
            .O(N__31460),
            .I(N__31453));
    InMux I__6146 (
            .O(N__31459),
            .I(N__31450));
    Odrv4 I__6145 (
            .O(N__31456),
            .I(\nx.n2689 ));
    Odrv4 I__6144 (
            .O(N__31453),
            .I(\nx.n2689 ));
    LocalMux I__6143 (
            .O(N__31450),
            .I(\nx.n2689 ));
    CascadeMux I__6142 (
            .O(N__31443),
            .I(\nx.n34_cascade_ ));
    CascadeMux I__6141 (
            .O(N__31440),
            .I(N__31436));
    InMux I__6140 (
            .O(N__31439),
            .I(N__31433));
    InMux I__6139 (
            .O(N__31436),
            .I(N__31429));
    LocalMux I__6138 (
            .O(N__31433),
            .I(N__31426));
    InMux I__6137 (
            .O(N__31432),
            .I(N__31423));
    LocalMux I__6136 (
            .O(N__31429),
            .I(N__31420));
    Odrv4 I__6135 (
            .O(N__31426),
            .I(\nx.n2799 ));
    LocalMux I__6134 (
            .O(N__31423),
            .I(\nx.n2799 ));
    Odrv4 I__6133 (
            .O(N__31420),
            .I(\nx.n2799 ));
    InMux I__6132 (
            .O(N__31413),
            .I(N__31410));
    LocalMux I__6131 (
            .O(N__31410),
            .I(N__31407));
    Span4Mux_v I__6130 (
            .O(N__31407),
            .I(N__31404));
    Odrv4 I__6129 (
            .O(N__31404),
            .I(\nx.n2866 ));
    CascadeMux I__6128 (
            .O(N__31401),
            .I(\nx.n2898_cascade_ ));
    InMux I__6127 (
            .O(N__31398),
            .I(N__31394));
    InMux I__6126 (
            .O(N__31397),
            .I(N__31391));
    LocalMux I__6125 (
            .O(N__31394),
            .I(\nx.n2997 ));
    LocalMux I__6124 (
            .O(N__31391),
            .I(\nx.n2997 ));
    CascadeMux I__6123 (
            .O(N__31386),
            .I(\nx.n2997_cascade_ ));
    InMux I__6122 (
            .O(N__31383),
            .I(N__31380));
    LocalMux I__6121 (
            .O(N__31380),
            .I(N__31377));
    Span4Mux_h I__6120 (
            .O(N__31377),
            .I(N__31374));
    Odrv4 I__6119 (
            .O(N__31374),
            .I(\nx.n45 ));
    InMux I__6118 (
            .O(N__31371),
            .I(N__31366));
    InMux I__6117 (
            .O(N__31370),
            .I(N__31363));
    InMux I__6116 (
            .O(N__31369),
            .I(N__31360));
    LocalMux I__6115 (
            .O(N__31366),
            .I(\nx.n2988 ));
    LocalMux I__6114 (
            .O(N__31363),
            .I(\nx.n2988 ));
    LocalMux I__6113 (
            .O(N__31360),
            .I(\nx.n2988 ));
    InMux I__6112 (
            .O(N__31353),
            .I(N__31350));
    LocalMux I__6111 (
            .O(N__31350),
            .I(N__31347));
    Span4Mux_h I__6110 (
            .O(N__31347),
            .I(N__31344));
    Odrv4 I__6109 (
            .O(N__31344),
            .I(\nx.n2855 ));
    CascadeMux I__6108 (
            .O(N__31341),
            .I(N__31338));
    InMux I__6107 (
            .O(N__31338),
            .I(N__31335));
    LocalMux I__6106 (
            .O(N__31335),
            .I(N__31332));
    Span4Mux_h I__6105 (
            .O(N__31332),
            .I(N__31328));
    InMux I__6104 (
            .O(N__31331),
            .I(N__31325));
    Odrv4 I__6103 (
            .O(N__31328),
            .I(\nx.n2788 ));
    LocalMux I__6102 (
            .O(N__31325),
            .I(\nx.n2788 ));
    InMux I__6101 (
            .O(N__31320),
            .I(N__31317));
    LocalMux I__6100 (
            .O(N__31317),
            .I(N__31314));
    Span4Mux_v I__6099 (
            .O(N__31314),
            .I(N__31311));
    Odrv4 I__6098 (
            .O(N__31311),
            .I(\nx.n2764 ));
    CascadeMux I__6097 (
            .O(N__31308),
            .I(N__31305));
    InMux I__6096 (
            .O(N__31305),
            .I(N__31302));
    LocalMux I__6095 (
            .O(N__31302),
            .I(N__31298));
    CascadeMux I__6094 (
            .O(N__31301),
            .I(N__31295));
    Span4Mux_h I__6093 (
            .O(N__31298),
            .I(N__31291));
    InMux I__6092 (
            .O(N__31295),
            .I(N__31288));
    InMux I__6091 (
            .O(N__31294),
            .I(N__31285));
    Odrv4 I__6090 (
            .O(N__31291),
            .I(\nx.n2697 ));
    LocalMux I__6089 (
            .O(N__31288),
            .I(\nx.n2697 ));
    LocalMux I__6088 (
            .O(N__31285),
            .I(\nx.n2697 ));
    CascadeMux I__6087 (
            .O(N__31278),
            .I(N__31271));
    CascadeMux I__6086 (
            .O(N__31277),
            .I(N__31265));
    CascadeMux I__6085 (
            .O(N__31276),
            .I(N__31262));
    CascadeMux I__6084 (
            .O(N__31275),
            .I(N__31256));
    InMux I__6083 (
            .O(N__31274),
            .I(N__31249));
    InMux I__6082 (
            .O(N__31271),
            .I(N__31244));
    InMux I__6081 (
            .O(N__31270),
            .I(N__31244));
    InMux I__6080 (
            .O(N__31269),
            .I(N__31231));
    InMux I__6079 (
            .O(N__31268),
            .I(N__31231));
    InMux I__6078 (
            .O(N__31265),
            .I(N__31231));
    InMux I__6077 (
            .O(N__31262),
            .I(N__31231));
    InMux I__6076 (
            .O(N__31261),
            .I(N__31231));
    InMux I__6075 (
            .O(N__31260),
            .I(N__31231));
    CascadeMux I__6074 (
            .O(N__31259),
            .I(N__31227));
    InMux I__6073 (
            .O(N__31256),
            .I(N__31223));
    CascadeMux I__6072 (
            .O(N__31255),
            .I(N__31217));
    CascadeMux I__6071 (
            .O(N__31254),
            .I(N__31213));
    CascadeMux I__6070 (
            .O(N__31253),
            .I(N__31209));
    CascadeMux I__6069 (
            .O(N__31252),
            .I(N__31206));
    LocalMux I__6068 (
            .O(N__31249),
            .I(N__31202));
    LocalMux I__6067 (
            .O(N__31244),
            .I(N__31199));
    LocalMux I__6066 (
            .O(N__31231),
            .I(N__31196));
    InMux I__6065 (
            .O(N__31230),
            .I(N__31189));
    InMux I__6064 (
            .O(N__31227),
            .I(N__31189));
    InMux I__6063 (
            .O(N__31226),
            .I(N__31189));
    LocalMux I__6062 (
            .O(N__31223),
            .I(N__31186));
    InMux I__6061 (
            .O(N__31222),
            .I(N__31181));
    InMux I__6060 (
            .O(N__31221),
            .I(N__31181));
    InMux I__6059 (
            .O(N__31220),
            .I(N__31172));
    InMux I__6058 (
            .O(N__31217),
            .I(N__31172));
    InMux I__6057 (
            .O(N__31216),
            .I(N__31172));
    InMux I__6056 (
            .O(N__31213),
            .I(N__31172));
    InMux I__6055 (
            .O(N__31212),
            .I(N__31163));
    InMux I__6054 (
            .O(N__31209),
            .I(N__31163));
    InMux I__6053 (
            .O(N__31206),
            .I(N__31163));
    InMux I__6052 (
            .O(N__31205),
            .I(N__31163));
    Span4Mux_v I__6051 (
            .O(N__31202),
            .I(N__31154));
    Span4Mux_v I__6050 (
            .O(N__31199),
            .I(N__31154));
    Span4Mux_v I__6049 (
            .O(N__31196),
            .I(N__31154));
    LocalMux I__6048 (
            .O(N__31189),
            .I(N__31154));
    Odrv4 I__6047 (
            .O(N__31186),
            .I(\nx.n2720 ));
    LocalMux I__6046 (
            .O(N__31181),
            .I(\nx.n2720 ));
    LocalMux I__6045 (
            .O(N__31172),
            .I(\nx.n2720 ));
    LocalMux I__6044 (
            .O(N__31163),
            .I(\nx.n2720 ));
    Odrv4 I__6043 (
            .O(N__31154),
            .I(\nx.n2720 ));
    CascadeMux I__6042 (
            .O(N__31143),
            .I(N__31140));
    InMux I__6041 (
            .O(N__31140),
            .I(N__31135));
    CascadeMux I__6040 (
            .O(N__31139),
            .I(N__31132));
    InMux I__6039 (
            .O(N__31138),
            .I(N__31129));
    LocalMux I__6038 (
            .O(N__31135),
            .I(N__31126));
    InMux I__6037 (
            .O(N__31132),
            .I(N__31123));
    LocalMux I__6036 (
            .O(N__31129),
            .I(N__31118));
    Span4Mux_h I__6035 (
            .O(N__31126),
            .I(N__31118));
    LocalMux I__6034 (
            .O(N__31123),
            .I(\nx.n2796 ));
    Odrv4 I__6033 (
            .O(N__31118),
            .I(\nx.n2796 ));
    InMux I__6032 (
            .O(N__31113),
            .I(N__31108));
    InMux I__6031 (
            .O(N__31112),
            .I(N__31105));
    InMux I__6030 (
            .O(N__31111),
            .I(N__31102));
    LocalMux I__6029 (
            .O(N__31108),
            .I(N__31099));
    LocalMux I__6028 (
            .O(N__31105),
            .I(\nx.n3000 ));
    LocalMux I__6027 (
            .O(N__31102),
            .I(\nx.n3000 ));
    Odrv4 I__6026 (
            .O(N__31099),
            .I(\nx.n3000 ));
    InMux I__6025 (
            .O(N__31092),
            .I(N__31088));
    InMux I__6024 (
            .O(N__31091),
            .I(N__31085));
    LocalMux I__6023 (
            .O(N__31088),
            .I(\nx.n3001 ));
    LocalMux I__6022 (
            .O(N__31085),
            .I(\nx.n3001 ));
    CascadeMux I__6021 (
            .O(N__31080),
            .I(\nx.n3001_cascade_ ));
    InMux I__6020 (
            .O(N__31077),
            .I(N__31074));
    LocalMux I__6019 (
            .O(N__31074),
            .I(N__31071));
    Odrv4 I__6018 (
            .O(N__31071),
            .I(\nx.n44 ));
    InMux I__6017 (
            .O(N__31068),
            .I(N__31063));
    InMux I__6016 (
            .O(N__31067),
            .I(N__31060));
    InMux I__6015 (
            .O(N__31066),
            .I(N__31057));
    LocalMux I__6014 (
            .O(N__31063),
            .I(\nx.n3003 ));
    LocalMux I__6013 (
            .O(N__31060),
            .I(\nx.n3003 ));
    LocalMux I__6012 (
            .O(N__31057),
            .I(\nx.n3003 ));
    InMux I__6011 (
            .O(N__31050),
            .I(N__31045));
    InMux I__6010 (
            .O(N__31049),
            .I(N__31042));
    InMux I__6009 (
            .O(N__31048),
            .I(N__31039));
    LocalMux I__6008 (
            .O(N__31045),
            .I(\nx.n3005 ));
    LocalMux I__6007 (
            .O(N__31042),
            .I(\nx.n3005 ));
    LocalMux I__6006 (
            .O(N__31039),
            .I(\nx.n3005 ));
    CascadeMux I__6005 (
            .O(N__31032),
            .I(N__31029));
    InMux I__6004 (
            .O(N__31029),
            .I(N__31026));
    LocalMux I__6003 (
            .O(N__31026),
            .I(N__31023));
    Span4Mux_v I__6002 (
            .O(N__31023),
            .I(N__31020));
    Odrv4 I__6001 (
            .O(N__31020),
            .I(\nx.n2863 ));
    CascadeMux I__6000 (
            .O(N__31017),
            .I(\nx.n2895_cascade_ ));
    CascadeMux I__5999 (
            .O(N__31014),
            .I(N__31009));
    InMux I__5998 (
            .O(N__31013),
            .I(N__31006));
    InMux I__5997 (
            .O(N__31012),
            .I(N__31003));
    InMux I__5996 (
            .O(N__31009),
            .I(N__31000));
    LocalMux I__5995 (
            .O(N__31006),
            .I(\nx.n2994 ));
    LocalMux I__5994 (
            .O(N__31003),
            .I(\nx.n2994 ));
    LocalMux I__5993 (
            .O(N__31000),
            .I(\nx.n2994 ));
    CascadeMux I__5992 (
            .O(N__30993),
            .I(\nx.n25_adj_748_cascade_ ));
    InMux I__5991 (
            .O(N__30990),
            .I(N__30987));
    LocalMux I__5990 (
            .O(N__30987),
            .I(\nx.n12785 ));
    InMux I__5989 (
            .O(N__30984),
            .I(N__30981));
    LocalMux I__5988 (
            .O(N__30981),
            .I(\nx.n19_adj_745 ));
    CascadeMux I__5987 (
            .O(N__30978),
            .I(\nx.n12777_cascade_ ));
    InMux I__5986 (
            .O(N__30975),
            .I(N__30972));
    LocalMux I__5985 (
            .O(N__30972),
            .I(\nx.n12779 ));
    CascadeMux I__5984 (
            .O(N__30969),
            .I(\nx.n39_adj_747_cascade_ ));
    InMux I__5983 (
            .O(N__30966),
            .I(N__30963));
    LocalMux I__5982 (
            .O(N__30963),
            .I(\nx.n12789 ));
    InMux I__5981 (
            .O(N__30960),
            .I(N__30957));
    LocalMux I__5980 (
            .O(N__30957),
            .I(N__30954));
    Odrv4 I__5979 (
            .O(N__30954),
            .I(\nx.n12799 ));
    InMux I__5978 (
            .O(N__30951),
            .I(N__30948));
    LocalMux I__5977 (
            .O(N__30948),
            .I(\nx.n29_adj_746 ));
    InMux I__5976 (
            .O(N__30945),
            .I(N__30942));
    LocalMux I__5975 (
            .O(N__30942),
            .I(N__30939));
    Span4Mux_h I__5974 (
            .O(N__30939),
            .I(N__30936));
    Odrv4 I__5973 (
            .O(N__30936),
            .I(\nx.n11_adj_751 ));
    InMux I__5972 (
            .O(N__30933),
            .I(N__30930));
    LocalMux I__5971 (
            .O(N__30930),
            .I(N__30927));
    Odrv4 I__5970 (
            .O(N__30927),
            .I(\nx.n41_adj_752 ));
    InMux I__5969 (
            .O(N__30924),
            .I(N__30921));
    LocalMux I__5968 (
            .O(N__30921),
            .I(N__30916));
    InMux I__5967 (
            .O(N__30920),
            .I(N__30913));
    InMux I__5966 (
            .O(N__30919),
            .I(N__30910));
    Span4Mux_v I__5965 (
            .O(N__30916),
            .I(N__30907));
    LocalMux I__5964 (
            .O(N__30913),
            .I(N__30904));
    LocalMux I__5963 (
            .O(N__30910),
            .I(N__30901));
    Odrv4 I__5962 (
            .O(N__30907),
            .I(\nx.n2989 ));
    Odrv4 I__5961 (
            .O(N__30904),
            .I(\nx.n2989 ));
    Odrv4 I__5960 (
            .O(N__30901),
            .I(\nx.n2989 ));
    CascadeMux I__5959 (
            .O(N__30894),
            .I(N__30891));
    InMux I__5958 (
            .O(N__30891),
            .I(N__30888));
    LocalMux I__5957 (
            .O(N__30888),
            .I(N__30884));
    InMux I__5956 (
            .O(N__30887),
            .I(N__30881));
    Span4Mux_v I__5955 (
            .O(N__30884),
            .I(N__30878));
    LocalMux I__5954 (
            .O(N__30881),
            .I(\nx.n2094 ));
    Odrv4 I__5953 (
            .O(N__30878),
            .I(\nx.n2094 ));
    InMux I__5952 (
            .O(N__30873),
            .I(N__30870));
    LocalMux I__5951 (
            .O(N__30870),
            .I(N__30867));
    Odrv4 I__5950 (
            .O(N__30867),
            .I(\nx.n2161 ));
    InMux I__5949 (
            .O(N__30864),
            .I(bfn_11_31_0_));
    InMux I__5948 (
            .O(N__30861),
            .I(N__30858));
    LocalMux I__5947 (
            .O(N__30858),
            .I(N__30855));
    Span4Mux_v I__5946 (
            .O(N__30855),
            .I(N__30851));
    InMux I__5945 (
            .O(N__30854),
            .I(N__30848));
    Odrv4 I__5944 (
            .O(N__30851),
            .I(\nx.n2093 ));
    LocalMux I__5943 (
            .O(N__30848),
            .I(\nx.n2093 ));
    InMux I__5942 (
            .O(N__30843),
            .I(\nx.n10880 ));
    CascadeMux I__5941 (
            .O(N__30840),
            .I(N__30837));
    InMux I__5940 (
            .O(N__30837),
            .I(N__30834));
    LocalMux I__5939 (
            .O(N__30834),
            .I(N__30830));
    InMux I__5938 (
            .O(N__30833),
            .I(N__30827));
    Span4Mux_h I__5937 (
            .O(N__30830),
            .I(N__30822));
    LocalMux I__5936 (
            .O(N__30827),
            .I(N__30822));
    Odrv4 I__5935 (
            .O(N__30822),
            .I(\nx.n2192 ));
    CascadeMux I__5934 (
            .O(N__30819),
            .I(\nx.n21_adj_750_cascade_ ));
    InMux I__5933 (
            .O(N__30816),
            .I(N__30812));
    InMux I__5932 (
            .O(N__30815),
            .I(N__30808));
    LocalMux I__5931 (
            .O(N__30812),
            .I(N__30805));
    InMux I__5930 (
            .O(N__30811),
            .I(N__30802));
    LocalMux I__5929 (
            .O(N__30808),
            .I(N__30799));
    Span4Mux_v I__5928 (
            .O(N__30805),
            .I(N__30796));
    LocalMux I__5927 (
            .O(N__30802),
            .I(N__30793));
    Span4Mux_v I__5926 (
            .O(N__30799),
            .I(N__30788));
    Span4Mux_v I__5925 (
            .O(N__30796),
            .I(N__30785));
    Span4Mux_v I__5924 (
            .O(N__30793),
            .I(N__30782));
    InMux I__5923 (
            .O(N__30792),
            .I(N__30779));
    InMux I__5922 (
            .O(N__30791),
            .I(N__30776));
    Span4Mux_v I__5921 (
            .O(N__30788),
            .I(N__30771));
    Span4Mux_h I__5920 (
            .O(N__30785),
            .I(N__30771));
    Odrv4 I__5919 (
            .O(N__30782),
            .I(\nx.bit_ctr_3 ));
    LocalMux I__5918 (
            .O(N__30779),
            .I(\nx.bit_ctr_3 ));
    LocalMux I__5917 (
            .O(N__30776),
            .I(\nx.bit_ctr_3 ));
    Odrv4 I__5916 (
            .O(N__30771),
            .I(\nx.bit_ctr_3 ));
    CascadeMux I__5915 (
            .O(N__30762),
            .I(\nx.n12781_cascade_ ));
    InMux I__5914 (
            .O(N__30759),
            .I(N__30756));
    LocalMux I__5913 (
            .O(N__30756),
            .I(N__30753));
    Odrv4 I__5912 (
            .O(N__30753),
            .I(\nx.n12801 ));
    CascadeMux I__5911 (
            .O(N__30750),
            .I(\nx.n27_adj_744_cascade_ ));
    InMux I__5910 (
            .O(N__30747),
            .I(N__30744));
    LocalMux I__5909 (
            .O(N__30744),
            .I(N__30740));
    InMux I__5908 (
            .O(N__30743),
            .I(N__30737));
    Odrv4 I__5907 (
            .O(N__30740),
            .I(\nx.n3209 ));
    LocalMux I__5906 (
            .O(N__30737),
            .I(\nx.n3209 ));
    InMux I__5905 (
            .O(N__30732),
            .I(bfn_11_30_0_));
    InMux I__5904 (
            .O(N__30729),
            .I(\nx.n10872 ));
    CascadeMux I__5903 (
            .O(N__30726),
            .I(N__30723));
    InMux I__5902 (
            .O(N__30723),
            .I(N__30719));
    InMux I__5901 (
            .O(N__30722),
            .I(N__30716));
    LocalMux I__5900 (
            .O(N__30719),
            .I(N__30713));
    LocalMux I__5899 (
            .O(N__30716),
            .I(N__30709));
    Span4Mux_h I__5898 (
            .O(N__30713),
            .I(N__30706));
    InMux I__5897 (
            .O(N__30712),
            .I(N__30703));
    Odrv4 I__5896 (
            .O(N__30709),
            .I(\nx.n2100 ));
    Odrv4 I__5895 (
            .O(N__30706),
            .I(\nx.n2100 ));
    LocalMux I__5894 (
            .O(N__30703),
            .I(\nx.n2100 ));
    CascadeMux I__5893 (
            .O(N__30696),
            .I(N__30693));
    InMux I__5892 (
            .O(N__30693),
            .I(N__30690));
    LocalMux I__5891 (
            .O(N__30690),
            .I(N__30687));
    Odrv4 I__5890 (
            .O(N__30687),
            .I(\nx.n2167 ));
    InMux I__5889 (
            .O(N__30684),
            .I(\nx.n10873 ));
    InMux I__5888 (
            .O(N__30681),
            .I(\nx.n10874 ));
    CascadeMux I__5887 (
            .O(N__30678),
            .I(N__30675));
    InMux I__5886 (
            .O(N__30675),
            .I(N__30672));
    LocalMux I__5885 (
            .O(N__30672),
            .I(N__30667));
    InMux I__5884 (
            .O(N__30671),
            .I(N__30664));
    InMux I__5883 (
            .O(N__30670),
            .I(N__30661));
    Span4Mux_s3_v I__5882 (
            .O(N__30667),
            .I(N__30658));
    LocalMux I__5881 (
            .O(N__30664),
            .I(N__30655));
    LocalMux I__5880 (
            .O(N__30661),
            .I(\nx.n2098 ));
    Odrv4 I__5879 (
            .O(N__30658),
            .I(\nx.n2098 ));
    Odrv4 I__5878 (
            .O(N__30655),
            .I(\nx.n2098 ));
    InMux I__5877 (
            .O(N__30648),
            .I(N__30645));
    LocalMux I__5876 (
            .O(N__30645),
            .I(N__30642));
    Odrv4 I__5875 (
            .O(N__30642),
            .I(\nx.n2165 ));
    InMux I__5874 (
            .O(N__30639),
            .I(\nx.n10875 ));
    CascadeMux I__5873 (
            .O(N__30636),
            .I(N__30632));
    InMux I__5872 (
            .O(N__30635),
            .I(N__30629));
    InMux I__5871 (
            .O(N__30632),
            .I(N__30625));
    LocalMux I__5870 (
            .O(N__30629),
            .I(N__30622));
    InMux I__5869 (
            .O(N__30628),
            .I(N__30619));
    LocalMux I__5868 (
            .O(N__30625),
            .I(\nx.n2097 ));
    Odrv4 I__5867 (
            .O(N__30622),
            .I(\nx.n2097 ));
    LocalMux I__5866 (
            .O(N__30619),
            .I(\nx.n2097 ));
    InMux I__5865 (
            .O(N__30612),
            .I(N__30609));
    LocalMux I__5864 (
            .O(N__30609),
            .I(N__30606));
    Odrv4 I__5863 (
            .O(N__30606),
            .I(\nx.n2164 ));
    InMux I__5862 (
            .O(N__30603),
            .I(\nx.n10876 ));
    CascadeMux I__5861 (
            .O(N__30600),
            .I(N__30597));
    InMux I__5860 (
            .O(N__30597),
            .I(N__30593));
    InMux I__5859 (
            .O(N__30596),
            .I(N__30590));
    LocalMux I__5858 (
            .O(N__30593),
            .I(N__30587));
    LocalMux I__5857 (
            .O(N__30590),
            .I(\nx.n2096 ));
    Odrv4 I__5856 (
            .O(N__30587),
            .I(\nx.n2096 ));
    CascadeMux I__5855 (
            .O(N__30582),
            .I(N__30579));
    InMux I__5854 (
            .O(N__30579),
            .I(N__30576));
    LocalMux I__5853 (
            .O(N__30576),
            .I(\nx.n2163 ));
    InMux I__5852 (
            .O(N__30573),
            .I(\nx.n10877 ));
    CascadeMux I__5851 (
            .O(N__30570),
            .I(N__30566));
    CascadeMux I__5850 (
            .O(N__30569),
            .I(N__30563));
    InMux I__5849 (
            .O(N__30566),
            .I(N__30559));
    InMux I__5848 (
            .O(N__30563),
            .I(N__30556));
    InMux I__5847 (
            .O(N__30562),
            .I(N__30553));
    LocalMux I__5846 (
            .O(N__30559),
            .I(\nx.n2095 ));
    LocalMux I__5845 (
            .O(N__30556),
            .I(\nx.n2095 ));
    LocalMux I__5844 (
            .O(N__30553),
            .I(\nx.n2095 ));
    InMux I__5843 (
            .O(N__30546),
            .I(N__30543));
    LocalMux I__5842 (
            .O(N__30543),
            .I(N__30540));
    Odrv4 I__5841 (
            .O(N__30540),
            .I(\nx.n2162 ));
    InMux I__5840 (
            .O(N__30537),
            .I(\nx.n10878 ));
    CascadeMux I__5839 (
            .O(N__30534),
            .I(N__30529));
    InMux I__5838 (
            .O(N__30533),
            .I(N__30525));
    InMux I__5837 (
            .O(N__30532),
            .I(N__30522));
    InMux I__5836 (
            .O(N__30529),
            .I(N__30519));
    InMux I__5835 (
            .O(N__30528),
            .I(N__30516));
    LocalMux I__5834 (
            .O(N__30525),
            .I(N__30511));
    LocalMux I__5833 (
            .O(N__30522),
            .I(N__30511));
    LocalMux I__5832 (
            .O(N__30519),
            .I(N__30507));
    LocalMux I__5831 (
            .O(N__30516),
            .I(N__30502));
    Span4Mux_v I__5830 (
            .O(N__30511),
            .I(N__30502));
    InMux I__5829 (
            .O(N__30510),
            .I(N__30499));
    Span4Mux_v I__5828 (
            .O(N__30507),
            .I(N__30496));
    Span4Mux_h I__5827 (
            .O(N__30502),
            .I(N__30493));
    LocalMux I__5826 (
            .O(N__30499),
            .I(\nx.bit_ctr_14 ));
    Odrv4 I__5825 (
            .O(N__30496),
            .I(\nx.bit_ctr_14 ));
    Odrv4 I__5824 (
            .O(N__30493),
            .I(\nx.bit_ctr_14 ));
    CascadeMux I__5823 (
            .O(N__30486),
            .I(N__30483));
    InMux I__5822 (
            .O(N__30483),
            .I(N__30480));
    LocalMux I__5821 (
            .O(N__30480),
            .I(N__30477));
    Odrv4 I__5820 (
            .O(N__30477),
            .I(\nx.n2177 ));
    InMux I__5819 (
            .O(N__30474),
            .I(bfn_11_29_0_));
    CascadeMux I__5818 (
            .O(N__30471),
            .I(N__30467));
    InMux I__5817 (
            .O(N__30470),
            .I(N__30464));
    InMux I__5816 (
            .O(N__30467),
            .I(N__30461));
    LocalMux I__5815 (
            .O(N__30464),
            .I(\nx.n2109 ));
    LocalMux I__5814 (
            .O(N__30461),
            .I(\nx.n2109 ));
    InMux I__5813 (
            .O(N__30456),
            .I(N__30453));
    LocalMux I__5812 (
            .O(N__30453),
            .I(\nx.n2176 ));
    InMux I__5811 (
            .O(N__30450),
            .I(\nx.n10864 ));
    CascadeMux I__5810 (
            .O(N__30447),
            .I(N__30443));
    InMux I__5809 (
            .O(N__30446),
            .I(N__30440));
    InMux I__5808 (
            .O(N__30443),
            .I(N__30437));
    LocalMux I__5807 (
            .O(N__30440),
            .I(\nx.n2108 ));
    LocalMux I__5806 (
            .O(N__30437),
            .I(\nx.n2108 ));
    InMux I__5805 (
            .O(N__30432),
            .I(N__30429));
    LocalMux I__5804 (
            .O(N__30429),
            .I(\nx.n2175 ));
    InMux I__5803 (
            .O(N__30426),
            .I(\nx.n10865 ));
    CascadeMux I__5802 (
            .O(N__30423),
            .I(N__30419));
    InMux I__5801 (
            .O(N__30422),
            .I(N__30416));
    InMux I__5800 (
            .O(N__30419),
            .I(N__30413));
    LocalMux I__5799 (
            .O(N__30416),
            .I(\nx.n2107 ));
    LocalMux I__5798 (
            .O(N__30413),
            .I(\nx.n2107 ));
    InMux I__5797 (
            .O(N__30408),
            .I(N__30405));
    LocalMux I__5796 (
            .O(N__30405),
            .I(\nx.n2174 ));
    InMux I__5795 (
            .O(N__30402),
            .I(\nx.n10866 ));
    InMux I__5794 (
            .O(N__30399),
            .I(N__30392));
    InMux I__5793 (
            .O(N__30398),
            .I(N__30392));
    InMux I__5792 (
            .O(N__30397),
            .I(N__30389));
    LocalMux I__5791 (
            .O(N__30392),
            .I(N__30384));
    LocalMux I__5790 (
            .O(N__30389),
            .I(N__30384));
    Odrv4 I__5789 (
            .O(N__30384),
            .I(\nx.n2106 ));
    InMux I__5788 (
            .O(N__30381),
            .I(N__30378));
    LocalMux I__5787 (
            .O(N__30378),
            .I(\nx.n2173 ));
    InMux I__5786 (
            .O(N__30375),
            .I(\nx.n10867 ));
    CascadeMux I__5785 (
            .O(N__30372),
            .I(N__30369));
    InMux I__5784 (
            .O(N__30369),
            .I(N__30366));
    LocalMux I__5783 (
            .O(N__30366),
            .I(N__30362));
    InMux I__5782 (
            .O(N__30365),
            .I(N__30359));
    Odrv4 I__5781 (
            .O(N__30362),
            .I(\nx.n2105 ));
    LocalMux I__5780 (
            .O(N__30359),
            .I(\nx.n2105 ));
    InMux I__5779 (
            .O(N__30354),
            .I(N__30351));
    LocalMux I__5778 (
            .O(N__30351),
            .I(N__30348));
    Odrv4 I__5777 (
            .O(N__30348),
            .I(\nx.n2172 ));
    InMux I__5776 (
            .O(N__30345),
            .I(\nx.n10868 ));
    CascadeMux I__5775 (
            .O(N__30342),
            .I(N__30339));
    InMux I__5774 (
            .O(N__30339),
            .I(N__30334));
    InMux I__5773 (
            .O(N__30338),
            .I(N__30331));
    InMux I__5772 (
            .O(N__30337),
            .I(N__30328));
    LocalMux I__5771 (
            .O(N__30334),
            .I(N__30325));
    LocalMux I__5770 (
            .O(N__30331),
            .I(\nx.n2104 ));
    LocalMux I__5769 (
            .O(N__30328),
            .I(\nx.n2104 ));
    Odrv4 I__5768 (
            .O(N__30325),
            .I(\nx.n2104 ));
    InMux I__5767 (
            .O(N__30318),
            .I(N__30315));
    LocalMux I__5766 (
            .O(N__30315),
            .I(\nx.n2171 ));
    InMux I__5765 (
            .O(N__30312),
            .I(\nx.n10869 ));
    CascadeMux I__5764 (
            .O(N__30309),
            .I(N__30306));
    InMux I__5763 (
            .O(N__30306),
            .I(N__30302));
    InMux I__5762 (
            .O(N__30305),
            .I(N__30299));
    LocalMux I__5761 (
            .O(N__30302),
            .I(N__30296));
    LocalMux I__5760 (
            .O(N__30299),
            .I(\nx.n2103 ));
    Odrv4 I__5759 (
            .O(N__30296),
            .I(\nx.n2103 ));
    InMux I__5758 (
            .O(N__30291),
            .I(N__30288));
    LocalMux I__5757 (
            .O(N__30288),
            .I(\nx.n2170 ));
    InMux I__5756 (
            .O(N__30285),
            .I(\nx.n10870 ));
    CascadeMux I__5755 (
            .O(N__30282),
            .I(N__30278));
    CascadeMux I__5754 (
            .O(N__30281),
            .I(N__30275));
    InMux I__5753 (
            .O(N__30278),
            .I(N__30270));
    InMux I__5752 (
            .O(N__30275),
            .I(N__30270));
    LocalMux I__5751 (
            .O(N__30270),
            .I(N__30267));
    Odrv4 I__5750 (
            .O(N__30267),
            .I(\nx.n2193 ));
    InMux I__5749 (
            .O(N__30264),
            .I(N__30261));
    LocalMux I__5748 (
            .O(N__30261),
            .I(\nx.n2260 ));
    InMux I__5747 (
            .O(N__30258),
            .I(N__30255));
    LocalMux I__5746 (
            .O(N__30255),
            .I(\nx.n29 ));
    InMux I__5745 (
            .O(N__30252),
            .I(N__30249));
    LocalMux I__5744 (
            .O(N__30249),
            .I(N__30246));
    Odrv4 I__5743 (
            .O(N__30246),
            .I(\nx.n28_adj_686 ));
    CascadeMux I__5742 (
            .O(N__30243),
            .I(N__30240));
    InMux I__5741 (
            .O(N__30240),
            .I(N__30237));
    LocalMux I__5740 (
            .O(N__30237),
            .I(\nx.n27_adj_691 ));
    InMux I__5739 (
            .O(N__30234),
            .I(N__30231));
    LocalMux I__5738 (
            .O(N__30231),
            .I(\nx.n30_adj_685 ));
    CascadeMux I__5737 (
            .O(N__30228),
            .I(\nx.n2126_cascade_ ));
    CascadeMux I__5736 (
            .O(N__30225),
            .I(\nx.n2199_cascade_ ));
    CascadeMux I__5735 (
            .O(N__30222),
            .I(\nx.n31_cascade_ ));
    InMux I__5734 (
            .O(N__30219),
            .I(N__30216));
    LocalMux I__5733 (
            .O(N__30216),
            .I(\nx.n28_adj_692 ));
    InMux I__5732 (
            .O(N__30213),
            .I(N__30210));
    LocalMux I__5731 (
            .O(N__30210),
            .I(N__30207));
    Span4Mux_h I__5730 (
            .O(N__30207),
            .I(N__30204));
    Odrv4 I__5729 (
            .O(N__30204),
            .I(\nx.n2264 ));
    InMux I__5728 (
            .O(N__30201),
            .I(\nx.n10893 ));
    InMux I__5727 (
            .O(N__30198),
            .I(\nx.n10894 ));
    InMux I__5726 (
            .O(N__30195),
            .I(\nx.n10895 ));
    InMux I__5725 (
            .O(N__30192),
            .I(bfn_11_27_0_));
    InMux I__5724 (
            .O(N__30189),
            .I(\nx.n10897 ));
    InMux I__5723 (
            .O(N__30186),
            .I(\nx.n10898 ));
    InMux I__5722 (
            .O(N__30183),
            .I(N__30180));
    LocalMux I__5721 (
            .O(N__30180),
            .I(\nx.n2263 ));
    CascadeMux I__5720 (
            .O(N__30177),
            .I(\nx.n2196_cascade_ ));
    InMux I__5719 (
            .O(N__30174),
            .I(\nx.n10884 ));
    InMux I__5718 (
            .O(N__30171),
            .I(\nx.n10885 ));
    InMux I__5717 (
            .O(N__30168),
            .I(\nx.n10886 ));
    InMux I__5716 (
            .O(N__30165),
            .I(\nx.n10887 ));
    InMux I__5715 (
            .O(N__30162),
            .I(bfn_11_26_0_));
    InMux I__5714 (
            .O(N__30159),
            .I(\nx.n10889 ));
    InMux I__5713 (
            .O(N__30156),
            .I(\nx.n10890 ));
    InMux I__5712 (
            .O(N__30153),
            .I(\nx.n10891 ));
    InMux I__5711 (
            .O(N__30150),
            .I(\nx.n10892 ));
    InMux I__5710 (
            .O(N__30147),
            .I(N__30143));
    InMux I__5709 (
            .O(N__30146),
            .I(N__30139));
    LocalMux I__5708 (
            .O(N__30143),
            .I(N__30136));
    InMux I__5707 (
            .O(N__30142),
            .I(N__30133));
    LocalMux I__5706 (
            .O(N__30139),
            .I(N__30129));
    Span4Mux_h I__5705 (
            .O(N__30136),
            .I(N__30124));
    LocalMux I__5704 (
            .O(N__30133),
            .I(N__30124));
    InMux I__5703 (
            .O(N__30132),
            .I(N__30120));
    Span4Mux_h I__5702 (
            .O(N__30129),
            .I(N__30115));
    Span4Mux_v I__5701 (
            .O(N__30124),
            .I(N__30115));
    InMux I__5700 (
            .O(N__30123),
            .I(N__30112));
    LocalMux I__5699 (
            .O(N__30120),
            .I(N__30109));
    Span4Mux_h I__5698 (
            .O(N__30115),
            .I(N__30106));
    LocalMux I__5697 (
            .O(N__30112),
            .I(N__30101));
    Span4Mux_h I__5696 (
            .O(N__30109),
            .I(N__30101));
    Odrv4 I__5695 (
            .O(N__30106),
            .I(\nx.bit_ctr_8 ));
    Odrv4 I__5694 (
            .O(N__30101),
            .I(\nx.bit_ctr_8 ));
    CascadeMux I__5693 (
            .O(N__30096),
            .I(\nx.n2698_cascade_ ));
    InMux I__5692 (
            .O(N__30093),
            .I(N__30090));
    LocalMux I__5691 (
            .O(N__30090),
            .I(\nx.n30 ));
    CascadeMux I__5690 (
            .O(N__30087),
            .I(N__30084));
    InMux I__5689 (
            .O(N__30084),
            .I(N__30080));
    CascadeMux I__5688 (
            .O(N__30083),
            .I(N__30077));
    LocalMux I__5687 (
            .O(N__30080),
            .I(N__30074));
    InMux I__5686 (
            .O(N__30077),
            .I(N__30071));
    Odrv4 I__5685 (
            .O(N__30074),
            .I(\nx.n2693 ));
    LocalMux I__5684 (
            .O(N__30071),
            .I(\nx.n2693 ));
    CascadeMux I__5683 (
            .O(N__30066),
            .I(N__30063));
    InMux I__5682 (
            .O(N__30063),
            .I(N__30059));
    CascadeMux I__5681 (
            .O(N__30062),
            .I(N__30056));
    LocalMux I__5680 (
            .O(N__30059),
            .I(N__30052));
    InMux I__5679 (
            .O(N__30056),
            .I(N__30049));
    InMux I__5678 (
            .O(N__30055),
            .I(N__30046));
    Odrv4 I__5677 (
            .O(N__30052),
            .I(\nx.n2694 ));
    LocalMux I__5676 (
            .O(N__30049),
            .I(\nx.n2694 ));
    LocalMux I__5675 (
            .O(N__30046),
            .I(\nx.n2694 ));
    CascadeMux I__5674 (
            .O(N__30039),
            .I(\nx.n2693_cascade_ ));
    CascadeMux I__5673 (
            .O(N__30036),
            .I(N__30032));
    InMux I__5672 (
            .O(N__30035),
            .I(N__30028));
    InMux I__5671 (
            .O(N__30032),
            .I(N__30025));
    InMux I__5670 (
            .O(N__30031),
            .I(N__30022));
    LocalMux I__5669 (
            .O(N__30028),
            .I(\nx.n2696 ));
    LocalMux I__5668 (
            .O(N__30025),
            .I(\nx.n2696 ));
    LocalMux I__5667 (
            .O(N__30022),
            .I(\nx.n2696 ));
    InMux I__5666 (
            .O(N__30015),
            .I(N__30012));
    LocalMux I__5665 (
            .O(N__30012),
            .I(\nx.n37_adj_677 ));
    CascadeMux I__5664 (
            .O(N__30009),
            .I(N__30006));
    InMux I__5663 (
            .O(N__30006),
            .I(N__30003));
    LocalMux I__5662 (
            .O(N__30003),
            .I(N__30000));
    Span4Mux_h I__5661 (
            .O(N__30000),
            .I(N__29996));
    CascadeMux I__5660 (
            .O(N__29999),
            .I(N__29992));
    Span4Mux_v I__5659 (
            .O(N__29996),
            .I(N__29989));
    InMux I__5658 (
            .O(N__29995),
            .I(N__29986));
    InMux I__5657 (
            .O(N__29992),
            .I(N__29983));
    Odrv4 I__5656 (
            .O(N__29989),
            .I(\nx.n2709 ));
    LocalMux I__5655 (
            .O(N__29986),
            .I(\nx.n2709 ));
    LocalMux I__5654 (
            .O(N__29983),
            .I(\nx.n2709 ));
    InMux I__5653 (
            .O(N__29976),
            .I(bfn_11_25_0_));
    InMux I__5652 (
            .O(N__29973),
            .I(\nx.n10881 ));
    InMux I__5651 (
            .O(N__29970),
            .I(\nx.n10882 ));
    InMux I__5650 (
            .O(N__29967),
            .I(\nx.n10883 ));
    CascadeMux I__5649 (
            .O(N__29964),
            .I(\nx.n2706_cascade_ ));
    InMux I__5648 (
            .O(N__29961),
            .I(N__29958));
    LocalMux I__5647 (
            .O(N__29958),
            .I(\nx.n40_adj_687 ));
    InMux I__5646 (
            .O(N__29955),
            .I(N__29952));
    LocalMux I__5645 (
            .O(N__29952),
            .I(N__29949));
    Odrv4 I__5644 (
            .O(N__29949),
            .I(\nx.n2755 ));
    CascadeMux I__5643 (
            .O(N__29946),
            .I(N__29943));
    InMux I__5642 (
            .O(N__29943),
            .I(N__29939));
    InMux I__5641 (
            .O(N__29942),
            .I(N__29935));
    LocalMux I__5640 (
            .O(N__29939),
            .I(N__29932));
    InMux I__5639 (
            .O(N__29938),
            .I(N__29929));
    LocalMux I__5638 (
            .O(N__29935),
            .I(\nx.n2787 ));
    Odrv4 I__5637 (
            .O(N__29932),
            .I(\nx.n2787 ));
    LocalMux I__5636 (
            .O(N__29929),
            .I(\nx.n2787 ));
    CascadeMux I__5635 (
            .O(N__29922),
            .I(N__29918));
    InMux I__5634 (
            .O(N__29921),
            .I(N__29915));
    InMux I__5633 (
            .O(N__29918),
            .I(N__29912));
    LocalMux I__5632 (
            .O(N__29915),
            .I(\nx.n2699 ));
    LocalMux I__5631 (
            .O(N__29912),
            .I(\nx.n2699 ));
    InMux I__5630 (
            .O(N__29907),
            .I(N__29904));
    LocalMux I__5629 (
            .O(N__29904),
            .I(\nx.n2766 ));
    CascadeMux I__5628 (
            .O(N__29901),
            .I(\nx.n2699_cascade_ ));
    CascadeMux I__5627 (
            .O(N__29898),
            .I(N__29895));
    InMux I__5626 (
            .O(N__29895),
            .I(N__29891));
    CascadeMux I__5625 (
            .O(N__29894),
            .I(N__29888));
    LocalMux I__5624 (
            .O(N__29891),
            .I(N__29885));
    InMux I__5623 (
            .O(N__29888),
            .I(N__29882));
    Odrv4 I__5622 (
            .O(N__29885),
            .I(\nx.n2701 ));
    LocalMux I__5621 (
            .O(N__29882),
            .I(\nx.n2701 ));
    CascadeMux I__5620 (
            .O(N__29877),
            .I(\nx.n2701_cascade_ ));
    CascadeMux I__5619 (
            .O(N__29874),
            .I(N__29871));
    InMux I__5618 (
            .O(N__29871),
            .I(N__29868));
    LocalMux I__5617 (
            .O(N__29868),
            .I(N__29865));
    Odrv4 I__5616 (
            .O(N__29865),
            .I(\nx.n42_adj_683 ));
    CascadeMux I__5615 (
            .O(N__29862),
            .I(N__29859));
    InMux I__5614 (
            .O(N__29859),
            .I(N__29855));
    CascadeMux I__5613 (
            .O(N__29858),
            .I(N__29852));
    LocalMux I__5612 (
            .O(N__29855),
            .I(N__29849));
    InMux I__5611 (
            .O(N__29852),
            .I(N__29846));
    Odrv4 I__5610 (
            .O(N__29849),
            .I(\nx.n2698 ));
    LocalMux I__5609 (
            .O(N__29846),
            .I(\nx.n2698 ));
    InMux I__5608 (
            .O(N__29841),
            .I(N__29838));
    LocalMux I__5607 (
            .O(N__29838),
            .I(N__29835));
    Odrv4 I__5606 (
            .O(N__29835),
            .I(\nx.n2765 ));
    InMux I__5605 (
            .O(N__29832),
            .I(N__29829));
    LocalMux I__5604 (
            .O(N__29829),
            .I(\nx.n41_adj_688 ));
    InMux I__5603 (
            .O(N__29826),
            .I(N__29823));
    LocalMux I__5602 (
            .O(N__29823),
            .I(N__29820));
    Odrv4 I__5601 (
            .O(N__29820),
            .I(\nx.n2767 ));
    CascadeMux I__5600 (
            .O(N__29817),
            .I(N__29814));
    InMux I__5599 (
            .O(N__29814),
            .I(N__29811));
    LocalMux I__5598 (
            .O(N__29811),
            .I(N__29808));
    Span4Mux_h I__5597 (
            .O(N__29808),
            .I(N__29805));
    Odrv4 I__5596 (
            .O(N__29805),
            .I(\nx.n2854 ));
    CascadeMux I__5595 (
            .O(N__29802),
            .I(\nx.n2886_cascade_ ));
    InMux I__5594 (
            .O(N__29799),
            .I(N__29794));
    InMux I__5593 (
            .O(N__29798),
            .I(N__29789));
    InMux I__5592 (
            .O(N__29797),
            .I(N__29789));
    LocalMux I__5591 (
            .O(N__29794),
            .I(\nx.n2985 ));
    LocalMux I__5590 (
            .O(N__29789),
            .I(\nx.n2985 ));
    CascadeMux I__5589 (
            .O(N__29784),
            .I(N__29781));
    InMux I__5588 (
            .O(N__29781),
            .I(N__29778));
    LocalMux I__5587 (
            .O(N__29778),
            .I(\nx.n2774 ));
    CascadeMux I__5586 (
            .O(N__29775),
            .I(N__29770));
    CascadeMux I__5585 (
            .O(N__29774),
            .I(N__29767));
    InMux I__5584 (
            .O(N__29773),
            .I(N__29764));
    InMux I__5583 (
            .O(N__29770),
            .I(N__29761));
    InMux I__5582 (
            .O(N__29767),
            .I(N__29758));
    LocalMux I__5581 (
            .O(N__29764),
            .I(\nx.n2800 ));
    LocalMux I__5580 (
            .O(N__29761),
            .I(\nx.n2800 ));
    LocalMux I__5579 (
            .O(N__29758),
            .I(\nx.n2800 ));
    InMux I__5578 (
            .O(N__29751),
            .I(N__29748));
    LocalMux I__5577 (
            .O(N__29748),
            .I(N__29745));
    Odrv4 I__5576 (
            .O(N__29745),
            .I(\nx.n2867 ));
    CascadeMux I__5575 (
            .O(N__29742),
            .I(N__29738));
    InMux I__5574 (
            .O(N__29741),
            .I(N__29735));
    InMux I__5573 (
            .O(N__29738),
            .I(N__29732));
    LocalMux I__5572 (
            .O(N__29735),
            .I(\nx.n2706 ));
    LocalMux I__5571 (
            .O(N__29732),
            .I(\nx.n2706 ));
    InMux I__5570 (
            .O(N__29727),
            .I(\nx.n11074 ));
    InMux I__5569 (
            .O(N__29724),
            .I(N__29720));
    InMux I__5568 (
            .O(N__29723),
            .I(N__29717));
    LocalMux I__5567 (
            .O(N__29720),
            .I(\nx.n2987 ));
    LocalMux I__5566 (
            .O(N__29717),
            .I(\nx.n2987 ));
    InMux I__5565 (
            .O(N__29712),
            .I(\nx.n11075 ));
    InMux I__5564 (
            .O(N__29709),
            .I(bfn_11_21_0_));
    InMux I__5563 (
            .O(N__29706),
            .I(\nx.n11077 ));
    CascadeMux I__5562 (
            .O(N__29703),
            .I(N__29698));
    CascadeMux I__5561 (
            .O(N__29702),
            .I(N__29695));
    CascadeMux I__5560 (
            .O(N__29701),
            .I(N__29692));
    InMux I__5559 (
            .O(N__29698),
            .I(N__29666));
    InMux I__5558 (
            .O(N__29695),
            .I(N__29661));
    InMux I__5557 (
            .O(N__29692),
            .I(N__29661));
    CascadeMux I__5556 (
            .O(N__29691),
            .I(N__29658));
    CascadeMux I__5555 (
            .O(N__29690),
            .I(N__29655));
    CascadeMux I__5554 (
            .O(N__29689),
            .I(N__29652));
    CascadeMux I__5553 (
            .O(N__29688),
            .I(N__29649));
    CascadeMux I__5552 (
            .O(N__29687),
            .I(N__29646));
    CascadeMux I__5551 (
            .O(N__29686),
            .I(N__29643));
    CascadeMux I__5550 (
            .O(N__29685),
            .I(N__29640));
    CascadeMux I__5549 (
            .O(N__29684),
            .I(N__29637));
    CascadeMux I__5548 (
            .O(N__29683),
            .I(N__29634));
    CascadeMux I__5547 (
            .O(N__29682),
            .I(N__29631));
    CascadeMux I__5546 (
            .O(N__29681),
            .I(N__29628));
    CascadeMux I__5545 (
            .O(N__29680),
            .I(N__29625));
    CascadeMux I__5544 (
            .O(N__29679),
            .I(N__29622));
    CascadeMux I__5543 (
            .O(N__29678),
            .I(N__29619));
    CascadeMux I__5542 (
            .O(N__29677),
            .I(N__29616));
    CascadeMux I__5541 (
            .O(N__29676),
            .I(N__29613));
    CascadeMux I__5540 (
            .O(N__29675),
            .I(N__29610));
    CascadeMux I__5539 (
            .O(N__29674),
            .I(N__29607));
    CascadeMux I__5538 (
            .O(N__29673),
            .I(N__29604));
    CascadeMux I__5537 (
            .O(N__29672),
            .I(N__29601));
    CascadeMux I__5536 (
            .O(N__29671),
            .I(N__29598));
    CascadeMux I__5535 (
            .O(N__29670),
            .I(N__29595));
    InMux I__5534 (
            .O(N__29669),
            .I(N__29592));
    LocalMux I__5533 (
            .O(N__29666),
            .I(N__29587));
    LocalMux I__5532 (
            .O(N__29661),
            .I(N__29587));
    InMux I__5531 (
            .O(N__29658),
            .I(N__29578));
    InMux I__5530 (
            .O(N__29655),
            .I(N__29578));
    InMux I__5529 (
            .O(N__29652),
            .I(N__29578));
    InMux I__5528 (
            .O(N__29649),
            .I(N__29578));
    InMux I__5527 (
            .O(N__29646),
            .I(N__29569));
    InMux I__5526 (
            .O(N__29643),
            .I(N__29569));
    InMux I__5525 (
            .O(N__29640),
            .I(N__29569));
    InMux I__5524 (
            .O(N__29637),
            .I(N__29569));
    InMux I__5523 (
            .O(N__29634),
            .I(N__29560));
    InMux I__5522 (
            .O(N__29631),
            .I(N__29560));
    InMux I__5521 (
            .O(N__29628),
            .I(N__29560));
    InMux I__5520 (
            .O(N__29625),
            .I(N__29560));
    InMux I__5519 (
            .O(N__29622),
            .I(N__29551));
    InMux I__5518 (
            .O(N__29619),
            .I(N__29551));
    InMux I__5517 (
            .O(N__29616),
            .I(N__29551));
    InMux I__5516 (
            .O(N__29613),
            .I(N__29551));
    InMux I__5515 (
            .O(N__29610),
            .I(N__29544));
    InMux I__5514 (
            .O(N__29607),
            .I(N__29544));
    InMux I__5513 (
            .O(N__29604),
            .I(N__29544));
    InMux I__5512 (
            .O(N__29601),
            .I(N__29537));
    InMux I__5511 (
            .O(N__29598),
            .I(N__29537));
    InMux I__5510 (
            .O(N__29595),
            .I(N__29537));
    LocalMux I__5509 (
            .O(N__29592),
            .I(N__29534));
    Odrv4 I__5508 (
            .O(N__29587),
            .I(\nx.n3017 ));
    LocalMux I__5507 (
            .O(N__29578),
            .I(\nx.n3017 ));
    LocalMux I__5506 (
            .O(N__29569),
            .I(\nx.n3017 ));
    LocalMux I__5505 (
            .O(N__29560),
            .I(\nx.n3017 ));
    LocalMux I__5504 (
            .O(N__29551),
            .I(\nx.n3017 ));
    LocalMux I__5503 (
            .O(N__29544),
            .I(\nx.n3017 ));
    LocalMux I__5502 (
            .O(N__29537),
            .I(\nx.n3017 ));
    Odrv4 I__5501 (
            .O(N__29534),
            .I(\nx.n3017 ));
    InMux I__5500 (
            .O(N__29517),
            .I(\nx.n11078 ));
    InMux I__5499 (
            .O(N__29514),
            .I(N__29511));
    LocalMux I__5498 (
            .O(N__29511),
            .I(N__29508));
    Odrv4 I__5497 (
            .O(N__29508),
            .I(\nx.n40_adj_670 ));
    InMux I__5496 (
            .O(N__29505),
            .I(N__29501));
    InMux I__5495 (
            .O(N__29504),
            .I(N__29498));
    LocalMux I__5494 (
            .O(N__29501),
            .I(N__29492));
    LocalMux I__5493 (
            .O(N__29498),
            .I(N__29492));
    InMux I__5492 (
            .O(N__29497),
            .I(N__29489));
    Odrv4 I__5491 (
            .O(N__29492),
            .I(\nx.n2996 ));
    LocalMux I__5490 (
            .O(N__29489),
            .I(\nx.n2996 ));
    InMux I__5489 (
            .O(N__29484),
            .I(N__29481));
    LocalMux I__5488 (
            .O(N__29481),
            .I(\nx.n41_adj_736 ));
    InMux I__5487 (
            .O(N__29478),
            .I(N__29473));
    InMux I__5486 (
            .O(N__29477),
            .I(N__29470));
    InMux I__5485 (
            .O(N__29476),
            .I(N__29467));
    LocalMux I__5484 (
            .O(N__29473),
            .I(N__29462));
    LocalMux I__5483 (
            .O(N__29470),
            .I(N__29462));
    LocalMux I__5482 (
            .O(N__29467),
            .I(N__29459));
    Span4Mux_v I__5481 (
            .O(N__29462),
            .I(N__29454));
    Span4Mux_h I__5480 (
            .O(N__29459),
            .I(N__29454));
    Odrv4 I__5479 (
            .O(N__29454),
            .I(\nx.n2998 ));
    InMux I__5478 (
            .O(N__29451),
            .I(\nx.n11065 ));
    InMux I__5477 (
            .O(N__29448),
            .I(\nx.n11066 ));
    InMux I__5476 (
            .O(N__29445),
            .I(\nx.n11067 ));
    InMux I__5475 (
            .O(N__29442),
            .I(bfn_11_20_0_));
    InMux I__5474 (
            .O(N__29439),
            .I(\nx.n11069 ));
    InMux I__5473 (
            .O(N__29436),
            .I(\nx.n11070 ));
    InMux I__5472 (
            .O(N__29433),
            .I(\nx.n11071 ));
    InMux I__5471 (
            .O(N__29430),
            .I(\nx.n11072 ));
    InMux I__5470 (
            .O(N__29427),
            .I(\nx.n11073 ));
    InMux I__5469 (
            .O(N__29424),
            .I(\nx.n11056 ));
    InMux I__5468 (
            .O(N__29421),
            .I(\nx.n11057 ));
    InMux I__5467 (
            .O(N__29418),
            .I(\nx.n11058 ));
    InMux I__5466 (
            .O(N__29415),
            .I(\nx.n11059 ));
    InMux I__5465 (
            .O(N__29412),
            .I(bfn_11_19_0_));
    InMux I__5464 (
            .O(N__29409),
            .I(\nx.n11061 ));
    InMux I__5463 (
            .O(N__29406),
            .I(\nx.n11062 ));
    InMux I__5462 (
            .O(N__29403),
            .I(\nx.n11063 ));
    InMux I__5461 (
            .O(N__29400),
            .I(\nx.n11064 ));
    CascadeMux I__5460 (
            .O(N__29397),
            .I(\nx.n42_adj_739_cascade_ ));
    CascadeMux I__5459 (
            .O(N__29394),
            .I(\nx.n32_adj_740_cascade_ ));
    InMux I__5458 (
            .O(N__29391),
            .I(N__29388));
    LocalMux I__5457 (
            .O(N__29388),
            .I(N__29385));
    Span4Mux_h I__5456 (
            .O(N__29385),
            .I(N__29382));
    Odrv4 I__5455 (
            .O(N__29382),
            .I(\nx.n44_adj_741 ));
    InMux I__5454 (
            .O(N__29379),
            .I(N__29376));
    LocalMux I__5453 (
            .O(N__29376),
            .I(\nx.n50_adj_742 ));
    InMux I__5452 (
            .O(N__29373),
            .I(N__29370));
    LocalMux I__5451 (
            .O(N__29370),
            .I(N__29367));
    Span4Mux_v I__5450 (
            .O(N__29367),
            .I(N__29364));
    Span4Mux_h I__5449 (
            .O(N__29364),
            .I(N__29361));
    Odrv4 I__5448 (
            .O(N__29361),
            .I(\nx.n47 ));
    CascadeMux I__5447 (
            .O(N__29358),
            .I(\nx.n49_cascade_ ));
    InMux I__5446 (
            .O(N__29355),
            .I(N__29352));
    LocalMux I__5445 (
            .O(N__29352),
            .I(\nx.n48 ));
    CascadeMux I__5444 (
            .O(N__29349),
            .I(\nx.n3116_cascade_ ));
    InMux I__5443 (
            .O(N__29346),
            .I(N__29342));
    InMux I__5442 (
            .O(N__29345),
            .I(N__29339));
    LocalMux I__5441 (
            .O(N__29342),
            .I(N__29333));
    LocalMux I__5440 (
            .O(N__29339),
            .I(N__29333));
    InMux I__5439 (
            .O(N__29338),
            .I(N__29330));
    Span4Mux_v I__5438 (
            .O(N__29333),
            .I(N__29325));
    LocalMux I__5437 (
            .O(N__29330),
            .I(N__29322));
    InMux I__5436 (
            .O(N__29329),
            .I(N__29319));
    InMux I__5435 (
            .O(N__29328),
            .I(N__29316));
    Span4Mux_h I__5434 (
            .O(N__29325),
            .I(N__29313));
    Span4Mux_h I__5433 (
            .O(N__29322),
            .I(N__29310));
    LocalMux I__5432 (
            .O(N__29319),
            .I(\nx.bit_ctr_5 ));
    LocalMux I__5431 (
            .O(N__29316),
            .I(\nx.bit_ctr_5 ));
    Odrv4 I__5430 (
            .O(N__29313),
            .I(\nx.bit_ctr_5 ));
    Odrv4 I__5429 (
            .O(N__29310),
            .I(\nx.bit_ctr_5 ));
    InMux I__5428 (
            .O(N__29301),
            .I(bfn_11_18_0_));
    InMux I__5427 (
            .O(N__29298),
            .I(N__29294));
    InMux I__5426 (
            .O(N__29297),
            .I(N__29291));
    LocalMux I__5425 (
            .O(N__29294),
            .I(N__29286));
    LocalMux I__5424 (
            .O(N__29291),
            .I(N__29286));
    Span4Mux_h I__5423 (
            .O(N__29286),
            .I(N__29283));
    Span4Mux_h I__5422 (
            .O(N__29283),
            .I(N__29280));
    Odrv4 I__5421 (
            .O(N__29280),
            .I(\nx.n3009 ));
    CascadeMux I__5420 (
            .O(N__29277),
            .I(N__29273));
    CascadeMux I__5419 (
            .O(N__29276),
            .I(N__29270));
    InMux I__5418 (
            .O(N__29273),
            .I(N__29267));
    InMux I__5417 (
            .O(N__29270),
            .I(N__29264));
    LocalMux I__5416 (
            .O(N__29267),
            .I(N__29259));
    LocalMux I__5415 (
            .O(N__29264),
            .I(N__29259));
    Span4Mux_h I__5414 (
            .O(N__29259),
            .I(N__29256));
    Odrv4 I__5413 (
            .O(N__29256),
            .I(\nx.n13600 ));
    InMux I__5412 (
            .O(N__29253),
            .I(\nx.n11053 ));
    InMux I__5411 (
            .O(N__29250),
            .I(N__29245));
    InMux I__5410 (
            .O(N__29249),
            .I(N__29242));
    InMux I__5409 (
            .O(N__29248),
            .I(N__29239));
    LocalMux I__5408 (
            .O(N__29245),
            .I(\nx.n3008 ));
    LocalMux I__5407 (
            .O(N__29242),
            .I(\nx.n3008 ));
    LocalMux I__5406 (
            .O(N__29239),
            .I(\nx.n3008 ));
    InMux I__5405 (
            .O(N__29232),
            .I(\nx.n11054 ));
    InMux I__5404 (
            .O(N__29229),
            .I(N__29224));
    InMux I__5403 (
            .O(N__29228),
            .I(N__29221));
    InMux I__5402 (
            .O(N__29227),
            .I(N__29218));
    LocalMux I__5401 (
            .O(N__29224),
            .I(\nx.n3007 ));
    LocalMux I__5400 (
            .O(N__29221),
            .I(\nx.n3007 ));
    LocalMux I__5399 (
            .O(N__29218),
            .I(\nx.n3007 ));
    InMux I__5398 (
            .O(N__29211),
            .I(\nx.n11055 ));
    CascadeMux I__5397 (
            .O(N__29208),
            .I(\nx.n2193_cascade_ ));
    InMux I__5396 (
            .O(N__29205),
            .I(N__29201));
    CascadeMux I__5395 (
            .O(N__29204),
            .I(N__29197));
    LocalMux I__5394 (
            .O(N__29201),
            .I(N__29194));
    InMux I__5393 (
            .O(N__29200),
            .I(N__29191));
    InMux I__5392 (
            .O(N__29197),
            .I(N__29188));
    Span4Mux_v I__5391 (
            .O(N__29194),
            .I(N__29181));
    LocalMux I__5390 (
            .O(N__29191),
            .I(N__29181));
    LocalMux I__5389 (
            .O(N__29188),
            .I(N__29181));
    Span4Mux_h I__5388 (
            .O(N__29181),
            .I(N__29178));
    Odrv4 I__5387 (
            .O(N__29178),
            .I(\nx.n2009 ));
    CascadeMux I__5386 (
            .O(N__29175),
            .I(N__29172));
    InMux I__5385 (
            .O(N__29172),
            .I(N__29169));
    LocalMux I__5384 (
            .O(N__29169),
            .I(N__29166));
    Span4Mux_v I__5383 (
            .O(N__29166),
            .I(N__29163));
    Odrv4 I__5382 (
            .O(N__29163),
            .I(\nx.n2076 ));
    CascadeMux I__5381 (
            .O(N__29160),
            .I(\nx.n2108_cascade_ ));
    CascadeMux I__5380 (
            .O(N__29157),
            .I(N__29154));
    InMux I__5379 (
            .O(N__29154),
            .I(N__29150));
    InMux I__5378 (
            .O(N__29153),
            .I(N__29147));
    LocalMux I__5377 (
            .O(N__29150),
            .I(N__29144));
    LocalMux I__5376 (
            .O(N__29147),
            .I(N__29140));
    Span4Mux_h I__5375 (
            .O(N__29144),
            .I(N__29137));
    InMux I__5374 (
            .O(N__29143),
            .I(N__29134));
    Odrv4 I__5373 (
            .O(N__29140),
            .I(\nx.n1996 ));
    Odrv4 I__5372 (
            .O(N__29137),
            .I(\nx.n1996 ));
    LocalMux I__5371 (
            .O(N__29134),
            .I(\nx.n1996 ));
    CascadeMux I__5370 (
            .O(N__29127),
            .I(N__29117));
    CascadeMux I__5369 (
            .O(N__29126),
            .I(N__29113));
    CascadeMux I__5368 (
            .O(N__29125),
            .I(N__29108));
    CascadeMux I__5367 (
            .O(N__29124),
            .I(N__29102));
    CascadeMux I__5366 (
            .O(N__29123),
            .I(N__29099));
    CascadeMux I__5365 (
            .O(N__29122),
            .I(N__29096));
    InMux I__5364 (
            .O(N__29121),
            .I(N__29089));
    InMux I__5363 (
            .O(N__29120),
            .I(N__29089));
    InMux I__5362 (
            .O(N__29117),
            .I(N__29084));
    InMux I__5361 (
            .O(N__29116),
            .I(N__29084));
    InMux I__5360 (
            .O(N__29113),
            .I(N__29075));
    InMux I__5359 (
            .O(N__29112),
            .I(N__29075));
    InMux I__5358 (
            .O(N__29111),
            .I(N__29075));
    InMux I__5357 (
            .O(N__29108),
            .I(N__29075));
    InMux I__5356 (
            .O(N__29107),
            .I(N__29068));
    InMux I__5355 (
            .O(N__29106),
            .I(N__29068));
    InMux I__5354 (
            .O(N__29105),
            .I(N__29068));
    InMux I__5353 (
            .O(N__29102),
            .I(N__29057));
    InMux I__5352 (
            .O(N__29099),
            .I(N__29057));
    InMux I__5351 (
            .O(N__29096),
            .I(N__29057));
    InMux I__5350 (
            .O(N__29095),
            .I(N__29057));
    InMux I__5349 (
            .O(N__29094),
            .I(N__29057));
    LocalMux I__5348 (
            .O(N__29089),
            .I(N__29048));
    LocalMux I__5347 (
            .O(N__29084),
            .I(N__29048));
    LocalMux I__5346 (
            .O(N__29075),
            .I(N__29048));
    LocalMux I__5345 (
            .O(N__29068),
            .I(N__29048));
    LocalMux I__5344 (
            .O(N__29057),
            .I(\nx.n2027 ));
    Odrv4 I__5343 (
            .O(N__29048),
            .I(\nx.n2027 ));
    InMux I__5342 (
            .O(N__29043),
            .I(N__29040));
    LocalMux I__5341 (
            .O(N__29040),
            .I(N__29037));
    Odrv4 I__5340 (
            .O(N__29037),
            .I(\nx.n2063 ));
    InMux I__5339 (
            .O(N__29034),
            .I(N__29031));
    LocalMux I__5338 (
            .O(N__29031),
            .I(N__29028));
    Odrv4 I__5337 (
            .O(N__29028),
            .I(\nx.n2075 ));
    CascadeMux I__5336 (
            .O(N__29025),
            .I(N__29022));
    InMux I__5335 (
            .O(N__29022),
            .I(N__29017));
    InMux I__5334 (
            .O(N__29021),
            .I(N__29014));
    CascadeMux I__5333 (
            .O(N__29020),
            .I(N__29011));
    LocalMux I__5332 (
            .O(N__29017),
            .I(N__29008));
    LocalMux I__5331 (
            .O(N__29014),
            .I(N__29005));
    InMux I__5330 (
            .O(N__29011),
            .I(N__29002));
    Span4Mux_v I__5329 (
            .O(N__29008),
            .I(N__28995));
    Span4Mux_h I__5328 (
            .O(N__29005),
            .I(N__28995));
    LocalMux I__5327 (
            .O(N__29002),
            .I(N__28995));
    Odrv4 I__5326 (
            .O(N__28995),
            .I(\nx.n2008 ));
    CascadeMux I__5325 (
            .O(N__28992),
            .I(\nx.n2107_cascade_ ));
    InMux I__5324 (
            .O(N__28989),
            .I(N__28986));
    LocalMux I__5323 (
            .O(N__28986),
            .I(\nx.n24_adj_684 ));
    InMux I__5322 (
            .O(N__28983),
            .I(N__28979));
    CascadeMux I__5321 (
            .O(N__28982),
            .I(N__28976));
    LocalMux I__5320 (
            .O(N__28979),
            .I(N__28973));
    InMux I__5319 (
            .O(N__28976),
            .I(N__28970));
    Span4Mux_v I__5318 (
            .O(N__28973),
            .I(N__28965));
    LocalMux I__5317 (
            .O(N__28970),
            .I(N__28965));
    Span4Mux_h I__5316 (
            .O(N__28965),
            .I(N__28961));
    InMux I__5315 (
            .O(N__28964),
            .I(N__28958));
    Odrv4 I__5314 (
            .O(N__28961),
            .I(\nx.n1997 ));
    LocalMux I__5313 (
            .O(N__28958),
            .I(\nx.n1997 ));
    CascadeMux I__5312 (
            .O(N__28953),
            .I(N__28950));
    InMux I__5311 (
            .O(N__28950),
            .I(N__28947));
    LocalMux I__5310 (
            .O(N__28947),
            .I(\nx.n2064 ));
    CascadeMux I__5309 (
            .O(N__28944),
            .I(\nx.n2096_cascade_ ));
    InMux I__5308 (
            .O(N__28941),
            .I(N__28938));
    LocalMux I__5307 (
            .O(N__28938),
            .I(N__28933));
    InMux I__5306 (
            .O(N__28937),
            .I(N__28930));
    InMux I__5305 (
            .O(N__28936),
            .I(N__28926));
    Span4Mux_v I__5304 (
            .O(N__28933),
            .I(N__28921));
    LocalMux I__5303 (
            .O(N__28930),
            .I(N__28921));
    InMux I__5302 (
            .O(N__28929),
            .I(N__28918));
    LocalMux I__5301 (
            .O(N__28926),
            .I(N__28914));
    Span4Mux_v I__5300 (
            .O(N__28921),
            .I(N__28909));
    LocalMux I__5299 (
            .O(N__28918),
            .I(N__28909));
    InMux I__5298 (
            .O(N__28917),
            .I(N__28906));
    Span4Mux_h I__5297 (
            .O(N__28914),
            .I(N__28903));
    Span4Mux_h I__5296 (
            .O(N__28909),
            .I(N__28900));
    LocalMux I__5295 (
            .O(N__28906),
            .I(\nx.bit_ctr_15 ));
    Odrv4 I__5294 (
            .O(N__28903),
            .I(\nx.bit_ctr_15 ));
    Odrv4 I__5293 (
            .O(N__28900),
            .I(\nx.bit_ctr_15 ));
    InMux I__5292 (
            .O(N__28893),
            .I(N__28890));
    LocalMux I__5291 (
            .O(N__28890),
            .I(N__28887));
    Span4Mux_v I__5290 (
            .O(N__28887),
            .I(N__28884));
    Odrv4 I__5289 (
            .O(N__28884),
            .I(\nx.n2077 ));
    CascadeMux I__5288 (
            .O(N__28881),
            .I(\nx.n2109_cascade_ ));
    CascadeMux I__5287 (
            .O(N__28878),
            .I(\nx.n2202_cascade_ ));
    InMux I__5286 (
            .O(N__28875),
            .I(N__28872));
    LocalMux I__5285 (
            .O(N__28872),
            .I(\nx.n18_adj_682 ));
    CascadeMux I__5284 (
            .O(N__28869),
            .I(N__28864));
    InMux I__5283 (
            .O(N__28868),
            .I(N__28859));
    InMux I__5282 (
            .O(N__28867),
            .I(N__28859));
    InMux I__5281 (
            .O(N__28864),
            .I(N__28856));
    LocalMux I__5280 (
            .O(N__28859),
            .I(N__28851));
    LocalMux I__5279 (
            .O(N__28856),
            .I(N__28851));
    Odrv4 I__5278 (
            .O(N__28851),
            .I(\nx.n2007 ));
    CascadeMux I__5277 (
            .O(N__28848),
            .I(N__28844));
    CascadeMux I__5276 (
            .O(N__28847),
            .I(N__28840));
    InMux I__5275 (
            .O(N__28844),
            .I(N__28837));
    InMux I__5274 (
            .O(N__28843),
            .I(N__28832));
    InMux I__5273 (
            .O(N__28840),
            .I(N__28832));
    LocalMux I__5272 (
            .O(N__28837),
            .I(N__28827));
    LocalMux I__5271 (
            .O(N__28832),
            .I(N__28827));
    Span4Mux_h I__5270 (
            .O(N__28827),
            .I(N__28824));
    Odrv4 I__5269 (
            .O(N__28824),
            .I(\nx.n2003 ));
    CascadeMux I__5268 (
            .O(N__28821),
            .I(N__28816));
    InMux I__5267 (
            .O(N__28820),
            .I(N__28813));
    InMux I__5266 (
            .O(N__28819),
            .I(N__28810));
    InMux I__5265 (
            .O(N__28816),
            .I(N__28807));
    LocalMux I__5264 (
            .O(N__28813),
            .I(N__28804));
    LocalMux I__5263 (
            .O(N__28810),
            .I(\nx.n2000 ));
    LocalMux I__5262 (
            .O(N__28807),
            .I(\nx.n2000 ));
    Odrv4 I__5261 (
            .O(N__28804),
            .I(\nx.n2000 ));
    InMux I__5260 (
            .O(N__28797),
            .I(N__28794));
    LocalMux I__5259 (
            .O(N__28794),
            .I(\nx.n27 ));
    InMux I__5258 (
            .O(N__28791),
            .I(N__28786));
    CascadeMux I__5257 (
            .O(N__28790),
            .I(N__28783));
    CascadeMux I__5256 (
            .O(N__28789),
            .I(N__28780));
    LocalMux I__5255 (
            .O(N__28786),
            .I(N__28777));
    InMux I__5254 (
            .O(N__28783),
            .I(N__28774));
    InMux I__5253 (
            .O(N__28780),
            .I(N__28771));
    Odrv4 I__5252 (
            .O(N__28777),
            .I(\nx.n2004 ));
    LocalMux I__5251 (
            .O(N__28774),
            .I(\nx.n2004 ));
    LocalMux I__5250 (
            .O(N__28771),
            .I(\nx.n2004 ));
    InMux I__5249 (
            .O(N__28764),
            .I(N__28761));
    LocalMux I__5248 (
            .O(N__28761),
            .I(\nx.n2071 ));
    CascadeMux I__5247 (
            .O(N__28758),
            .I(\nx.n2103_cascade_ ));
    CascadeMux I__5246 (
            .O(N__28755),
            .I(N__28751));
    InMux I__5245 (
            .O(N__28754),
            .I(N__28748));
    InMux I__5244 (
            .O(N__28751),
            .I(N__28745));
    LocalMux I__5243 (
            .O(N__28748),
            .I(N__28741));
    LocalMux I__5242 (
            .O(N__28745),
            .I(N__28738));
    InMux I__5241 (
            .O(N__28744),
            .I(N__28735));
    Odrv4 I__5240 (
            .O(N__28741),
            .I(\nx.n1998 ));
    Odrv4 I__5239 (
            .O(N__28738),
            .I(\nx.n1998 ));
    LocalMux I__5238 (
            .O(N__28735),
            .I(\nx.n1998 ));
    InMux I__5237 (
            .O(N__28728),
            .I(N__28725));
    LocalMux I__5236 (
            .O(N__28725),
            .I(\nx.n2065 ));
    InMux I__5235 (
            .O(N__28722),
            .I(N__28719));
    LocalMux I__5234 (
            .O(N__28719),
            .I(\nx.n2073 ));
    CascadeMux I__5233 (
            .O(N__28716),
            .I(N__28713));
    InMux I__5232 (
            .O(N__28713),
            .I(N__28708));
    InMux I__5231 (
            .O(N__28712),
            .I(N__28705));
    CascadeMux I__5230 (
            .O(N__28711),
            .I(N__28702));
    LocalMux I__5229 (
            .O(N__28708),
            .I(N__28699));
    LocalMux I__5228 (
            .O(N__28705),
            .I(N__28696));
    InMux I__5227 (
            .O(N__28702),
            .I(N__28693));
    Span4Mux_v I__5226 (
            .O(N__28699),
            .I(N__28686));
    Span4Mux_h I__5225 (
            .O(N__28696),
            .I(N__28686));
    LocalMux I__5224 (
            .O(N__28693),
            .I(N__28686));
    Odrv4 I__5223 (
            .O(N__28686),
            .I(\nx.n2006 ));
    CascadeMux I__5222 (
            .O(N__28683),
            .I(\nx.n2105_cascade_ ));
    InMux I__5221 (
            .O(N__28680),
            .I(N__28676));
    CascadeMux I__5220 (
            .O(N__28679),
            .I(N__28673));
    LocalMux I__5219 (
            .O(N__28676),
            .I(N__28669));
    InMux I__5218 (
            .O(N__28673),
            .I(N__28666));
    InMux I__5217 (
            .O(N__28672),
            .I(N__28663));
    Span4Mux_v I__5216 (
            .O(N__28669),
            .I(N__28656));
    LocalMux I__5215 (
            .O(N__28666),
            .I(N__28656));
    LocalMux I__5214 (
            .O(N__28663),
            .I(N__28656));
    Odrv4 I__5213 (
            .O(N__28656),
            .I(\nx.n2005 ));
    CascadeMux I__5212 (
            .O(N__28653),
            .I(N__28650));
    InMux I__5211 (
            .O(N__28650),
            .I(N__28647));
    LocalMux I__5210 (
            .O(N__28647),
            .I(\nx.n2072 ));
    CascadeMux I__5209 (
            .O(N__28644),
            .I(N__28640));
    InMux I__5208 (
            .O(N__28643),
            .I(N__28637));
    InMux I__5207 (
            .O(N__28640),
            .I(N__28633));
    LocalMux I__5206 (
            .O(N__28637),
            .I(N__28630));
    InMux I__5205 (
            .O(N__28636),
            .I(N__28627));
    LocalMux I__5204 (
            .O(N__28633),
            .I(N__28624));
    Odrv4 I__5203 (
            .O(N__28630),
            .I(\nx.n2002 ));
    LocalMux I__5202 (
            .O(N__28627),
            .I(\nx.n2002 ));
    Odrv4 I__5201 (
            .O(N__28624),
            .I(\nx.n2002 ));
    InMux I__5200 (
            .O(N__28617),
            .I(N__28614));
    LocalMux I__5199 (
            .O(N__28614),
            .I(\nx.n2069 ));
    InMux I__5198 (
            .O(N__28611),
            .I(\nx.n11003 ));
    CascadeMux I__5197 (
            .O(N__28608),
            .I(N__28604));
    InMux I__5196 (
            .O(N__28607),
            .I(N__28601));
    InMux I__5195 (
            .O(N__28604),
            .I(N__28598));
    LocalMux I__5194 (
            .O(N__28601),
            .I(N__28595));
    LocalMux I__5193 (
            .O(N__28598),
            .I(\nx.n2786 ));
    Odrv12 I__5192 (
            .O(N__28595),
            .I(\nx.n2786 ));
    CascadeMux I__5191 (
            .O(N__28590),
            .I(N__28587));
    InMux I__5190 (
            .O(N__28587),
            .I(N__28584));
    LocalMux I__5189 (
            .O(N__28584),
            .I(\nx.n2070 ));
    CascadeMux I__5188 (
            .O(N__28581),
            .I(\nx.n9709_cascade_ ));
    InMux I__5187 (
            .O(N__28578),
            .I(N__28575));
    LocalMux I__5186 (
            .O(N__28575),
            .I(N__28572));
    Span4Mux_h I__5185 (
            .O(N__28572),
            .I(N__28569));
    Odrv4 I__5184 (
            .O(N__28569),
            .I(\nx.n25 ));
    CascadeMux I__5183 (
            .O(N__28566),
            .I(\nx.n26_adj_681_cascade_ ));
    CascadeMux I__5182 (
            .O(N__28563),
            .I(\nx.n2027_cascade_ ));
    InMux I__5181 (
            .O(N__28560),
            .I(N__28557));
    LocalMux I__5180 (
            .O(N__28557),
            .I(\nx.n2074 ));
    CascadeMux I__5179 (
            .O(N__28554),
            .I(N__28550));
    InMux I__5178 (
            .O(N__28553),
            .I(N__28547));
    InMux I__5177 (
            .O(N__28550),
            .I(N__28544));
    LocalMux I__5176 (
            .O(N__28547),
            .I(N__28541));
    LocalMux I__5175 (
            .O(N__28544),
            .I(\nx.n2001 ));
    Odrv4 I__5174 (
            .O(N__28541),
            .I(\nx.n2001 ));
    InMux I__5173 (
            .O(N__28536),
            .I(N__28533));
    LocalMux I__5172 (
            .O(N__28533),
            .I(\nx.n28_adj_680 ));
    CascadeMux I__5171 (
            .O(N__28530),
            .I(N__28527));
    InMux I__5170 (
            .O(N__28527),
            .I(N__28524));
    LocalMux I__5169 (
            .O(N__28524),
            .I(N__28519));
    InMux I__5168 (
            .O(N__28523),
            .I(N__28514));
    InMux I__5167 (
            .O(N__28522),
            .I(N__28514));
    Odrv4 I__5166 (
            .O(N__28519),
            .I(\nx.n1999 ));
    LocalMux I__5165 (
            .O(N__28514),
            .I(\nx.n1999 ));
    CascadeMux I__5164 (
            .O(N__28509),
            .I(N__28506));
    InMux I__5163 (
            .O(N__28506),
            .I(N__28503));
    LocalMux I__5162 (
            .O(N__28503),
            .I(\nx.n2066 ));
    InMux I__5161 (
            .O(N__28500),
            .I(N__28497));
    LocalMux I__5160 (
            .O(N__28497),
            .I(N__28494));
    Odrv4 I__5159 (
            .O(N__28494),
            .I(\nx.n2763 ));
    InMux I__5158 (
            .O(N__28491),
            .I(\nx.n10994 ));
    CascadeMux I__5157 (
            .O(N__28488),
            .I(N__28485));
    InMux I__5156 (
            .O(N__28485),
            .I(N__28482));
    LocalMux I__5155 (
            .O(N__28482),
            .I(\nx.n2762 ));
    InMux I__5154 (
            .O(N__28479),
            .I(\nx.n10995 ));
    InMux I__5153 (
            .O(N__28476),
            .I(N__28473));
    LocalMux I__5152 (
            .O(N__28473),
            .I(\nx.n2761 ));
    InMux I__5151 (
            .O(N__28470),
            .I(bfn_10_25_0_));
    InMux I__5150 (
            .O(N__28467),
            .I(N__28464));
    LocalMux I__5149 (
            .O(N__28464),
            .I(\nx.n2760 ));
    InMux I__5148 (
            .O(N__28461),
            .I(\nx.n10997 ));
    InMux I__5147 (
            .O(N__28458),
            .I(N__28455));
    LocalMux I__5146 (
            .O(N__28455),
            .I(N__28452));
    Span4Mux_v I__5145 (
            .O(N__28452),
            .I(N__28449));
    Odrv4 I__5144 (
            .O(N__28449),
            .I(\nx.n2759 ));
    InMux I__5143 (
            .O(N__28446),
            .I(\nx.n10998 ));
    InMux I__5142 (
            .O(N__28443),
            .I(N__28440));
    LocalMux I__5141 (
            .O(N__28440),
            .I(\nx.n2758 ));
    InMux I__5140 (
            .O(N__28437),
            .I(\nx.n10999 ));
    InMux I__5139 (
            .O(N__28434),
            .I(N__28431));
    LocalMux I__5138 (
            .O(N__28431),
            .I(\nx.n2757 ));
    InMux I__5137 (
            .O(N__28428),
            .I(\nx.n11000 ));
    InMux I__5136 (
            .O(N__28425),
            .I(N__28422));
    LocalMux I__5135 (
            .O(N__28422),
            .I(N__28419));
    Odrv4 I__5134 (
            .O(N__28419),
            .I(\nx.n2756 ));
    InMux I__5133 (
            .O(N__28416),
            .I(\nx.n11001 ));
    InMux I__5132 (
            .O(N__28413),
            .I(\nx.n11002 ));
    InMux I__5131 (
            .O(N__28410),
            .I(\nx.n10985 ));
    InMux I__5130 (
            .O(N__28407),
            .I(N__28404));
    LocalMux I__5129 (
            .O(N__28404),
            .I(N__28401));
    Odrv12 I__5128 (
            .O(N__28401),
            .I(\nx.n2771 ));
    InMux I__5127 (
            .O(N__28398),
            .I(\nx.n10986 ));
    CascadeMux I__5126 (
            .O(N__28395),
            .I(N__28392));
    InMux I__5125 (
            .O(N__28392),
            .I(N__28389));
    LocalMux I__5124 (
            .O(N__28389),
            .I(N__28386));
    Odrv12 I__5123 (
            .O(N__28386),
            .I(\nx.n2770 ));
    InMux I__5122 (
            .O(N__28383),
            .I(\nx.n10987 ));
    InMux I__5121 (
            .O(N__28380),
            .I(N__28377));
    LocalMux I__5120 (
            .O(N__28377),
            .I(\nx.n2769 ));
    InMux I__5119 (
            .O(N__28374),
            .I(bfn_10_24_0_));
    InMux I__5118 (
            .O(N__28371),
            .I(N__28368));
    LocalMux I__5117 (
            .O(N__28368),
            .I(N__28365));
    Odrv4 I__5116 (
            .O(N__28365),
            .I(\nx.n2768 ));
    InMux I__5115 (
            .O(N__28362),
            .I(\nx.n10989 ));
    InMux I__5114 (
            .O(N__28359),
            .I(\nx.n10990 ));
    InMux I__5113 (
            .O(N__28356),
            .I(\nx.n10991 ));
    InMux I__5112 (
            .O(N__28353),
            .I(\nx.n10992 ));
    InMux I__5111 (
            .O(N__28350),
            .I(\nx.n10993 ));
    CascadeMux I__5110 (
            .O(N__28347),
            .I(\nx.n2788_cascade_ ));
    CascadeMux I__5109 (
            .O(N__28344),
            .I(N__28341));
    InMux I__5108 (
            .O(N__28341),
            .I(N__28337));
    CascadeMux I__5107 (
            .O(N__28340),
            .I(N__28333));
    LocalMux I__5106 (
            .O(N__28337),
            .I(N__28330));
    InMux I__5105 (
            .O(N__28336),
            .I(N__28327));
    InMux I__5104 (
            .O(N__28333),
            .I(N__28324));
    Span4Mux_h I__5103 (
            .O(N__28330),
            .I(N__28319));
    LocalMux I__5102 (
            .O(N__28327),
            .I(N__28319));
    LocalMux I__5101 (
            .O(N__28324),
            .I(\nx.n2789 ));
    Odrv4 I__5100 (
            .O(N__28319),
            .I(\nx.n2789 ));
    CascadeMux I__5099 (
            .O(N__28314),
            .I(\nx.n26_adj_706_cascade_ ));
    InMux I__5098 (
            .O(N__28311),
            .I(N__28308));
    LocalMux I__5097 (
            .O(N__28308),
            .I(N__28305));
    Odrv4 I__5096 (
            .O(N__28305),
            .I(\nx.n38_adj_713 ));
    InMux I__5095 (
            .O(N__28302),
            .I(N__28299));
    LocalMux I__5094 (
            .O(N__28299),
            .I(N__28296));
    Odrv4 I__5093 (
            .O(N__28296),
            .I(\nx.n43_adj_735 ));
    InMux I__5092 (
            .O(N__28293),
            .I(N__28290));
    LocalMux I__5091 (
            .O(N__28290),
            .I(N__28287));
    Span4Mux_v I__5090 (
            .O(N__28287),
            .I(N__28284));
    Odrv4 I__5089 (
            .O(N__28284),
            .I(\nx.n2777 ));
    InMux I__5088 (
            .O(N__28281),
            .I(bfn_10_23_0_));
    InMux I__5087 (
            .O(N__28278),
            .I(N__28275));
    LocalMux I__5086 (
            .O(N__28275),
            .I(N__28272));
    Span4Mux_v I__5085 (
            .O(N__28272),
            .I(N__28269));
    Odrv4 I__5084 (
            .O(N__28269),
            .I(\nx.n2776 ));
    InMux I__5083 (
            .O(N__28266),
            .I(\nx.n10981 ));
    InMux I__5082 (
            .O(N__28263),
            .I(N__28260));
    LocalMux I__5081 (
            .O(N__28260),
            .I(N__28257));
    Odrv4 I__5080 (
            .O(N__28257),
            .I(\nx.n2775 ));
    InMux I__5079 (
            .O(N__28254),
            .I(\nx.n10982 ));
    InMux I__5078 (
            .O(N__28251),
            .I(\nx.n10983 ));
    InMux I__5077 (
            .O(N__28248),
            .I(N__28245));
    LocalMux I__5076 (
            .O(N__28245),
            .I(\nx.n2773 ));
    InMux I__5075 (
            .O(N__28242),
            .I(\nx.n10984 ));
    InMux I__5074 (
            .O(N__28239),
            .I(N__28236));
    LocalMux I__5073 (
            .O(N__28236),
            .I(\nx.n2772 ));
    InMux I__5072 (
            .O(N__28233),
            .I(N__28230));
    LocalMux I__5071 (
            .O(N__28230),
            .I(N__28226));
    InMux I__5070 (
            .O(N__28229),
            .I(N__28223));
    Odrv4 I__5069 (
            .O(N__28226),
            .I(\nx.n2809 ));
    LocalMux I__5068 (
            .O(N__28223),
            .I(\nx.n2809 ));
    CascadeMux I__5067 (
            .O(N__28218),
            .I(\nx.n2809_cascade_ ));
    InMux I__5066 (
            .O(N__28215),
            .I(N__28210));
    InMux I__5065 (
            .O(N__28214),
            .I(N__28207));
    InMux I__5064 (
            .O(N__28213),
            .I(N__28202));
    LocalMux I__5063 (
            .O(N__28210),
            .I(N__28199));
    LocalMux I__5062 (
            .O(N__28207),
            .I(N__28196));
    InMux I__5061 (
            .O(N__28206),
            .I(N__28193));
    InMux I__5060 (
            .O(N__28205),
            .I(N__28190));
    LocalMux I__5059 (
            .O(N__28202),
            .I(N__28187));
    Span4Mux_v I__5058 (
            .O(N__28199),
            .I(N__28180));
    Span4Mux_h I__5057 (
            .O(N__28196),
            .I(N__28180));
    LocalMux I__5056 (
            .O(N__28193),
            .I(N__28180));
    LocalMux I__5055 (
            .O(N__28190),
            .I(N__28175));
    Span4Mux_v I__5054 (
            .O(N__28187),
            .I(N__28175));
    Span4Mux_h I__5053 (
            .O(N__28180),
            .I(N__28172));
    Odrv4 I__5052 (
            .O(N__28175),
            .I(\nx.bit_ctr_7 ));
    Odrv4 I__5051 (
            .O(N__28172),
            .I(\nx.bit_ctr_7 ));
    InMux I__5050 (
            .O(N__28167),
            .I(N__28164));
    LocalMux I__5049 (
            .O(N__28164),
            .I(\nx.n30_adj_704 ));
    CascadeMux I__5048 (
            .O(N__28161),
            .I(N__28157));
    InMux I__5047 (
            .O(N__28160),
            .I(N__28154));
    InMux I__5046 (
            .O(N__28157),
            .I(N__28151));
    LocalMux I__5045 (
            .O(N__28154),
            .I(\nx.n2802 ));
    LocalMux I__5044 (
            .O(N__28151),
            .I(\nx.n2802 ));
    InMux I__5043 (
            .O(N__28146),
            .I(N__28143));
    LocalMux I__5042 (
            .O(N__28143),
            .I(\nx.n2869 ));
    CascadeMux I__5041 (
            .O(N__28140),
            .I(\nx.n2802_cascade_ ));
    InMux I__5040 (
            .O(N__28137),
            .I(N__28133));
    CascadeMux I__5039 (
            .O(N__28136),
            .I(N__28130));
    LocalMux I__5038 (
            .O(N__28133),
            .I(N__28126));
    InMux I__5037 (
            .O(N__28130),
            .I(N__28123));
    InMux I__5036 (
            .O(N__28129),
            .I(N__28120));
    Odrv4 I__5035 (
            .O(N__28126),
            .I(\nx.n2795 ));
    LocalMux I__5034 (
            .O(N__28123),
            .I(\nx.n2795 ));
    LocalMux I__5033 (
            .O(N__28120),
            .I(\nx.n2795 ));
    CascadeMux I__5032 (
            .O(N__28113),
            .I(\nx.n2720_cascade_ ));
    InMux I__5031 (
            .O(N__28110),
            .I(N__28103));
    InMux I__5030 (
            .O(N__28109),
            .I(N__28103));
    CascadeMux I__5029 (
            .O(N__28108),
            .I(N__28100));
    LocalMux I__5028 (
            .O(N__28103),
            .I(N__28097));
    InMux I__5027 (
            .O(N__28100),
            .I(N__28094));
    Span4Mux_h I__5026 (
            .O(N__28097),
            .I(N__28091));
    LocalMux I__5025 (
            .O(N__28094),
            .I(N__28088));
    Odrv4 I__5024 (
            .O(N__28091),
            .I(\nx.n2801 ));
    Odrv4 I__5023 (
            .O(N__28088),
            .I(\nx.n2801 ));
    CascadeMux I__5022 (
            .O(N__28083),
            .I(N__28078));
    InMux I__5021 (
            .O(N__28082),
            .I(N__28075));
    InMux I__5020 (
            .O(N__28081),
            .I(N__28072));
    InMux I__5019 (
            .O(N__28078),
            .I(N__28069));
    LocalMux I__5018 (
            .O(N__28075),
            .I(\nx.n2808 ));
    LocalMux I__5017 (
            .O(N__28072),
            .I(\nx.n2808 ));
    LocalMux I__5016 (
            .O(N__28069),
            .I(\nx.n2808 ));
    CascadeMux I__5015 (
            .O(N__28062),
            .I(\nx.n40_adj_705_cascade_ ));
    CascadeMux I__5014 (
            .O(N__28059),
            .I(\nx.n44_adj_721_cascade_ ));
    InMux I__5013 (
            .O(N__28056),
            .I(N__28053));
    LocalMux I__5012 (
            .O(N__28053),
            .I(N__28050));
    Odrv4 I__5011 (
            .O(N__28050),
            .I(\nx.n2862 ));
    CascadeMux I__5010 (
            .O(N__28047),
            .I(\nx.n2819_cascade_ ));
    InMux I__5009 (
            .O(N__28044),
            .I(N__28041));
    LocalMux I__5008 (
            .O(N__28041),
            .I(\nx.n2874 ));
    InMux I__5007 (
            .O(N__28038),
            .I(N__28035));
    LocalMux I__5006 (
            .O(N__28035),
            .I(\nx.n42_adj_730 ));
    CascadeMux I__5005 (
            .O(N__28032),
            .I(N__28028));
    CascadeMux I__5004 (
            .O(N__28031),
            .I(N__28024));
    InMux I__5003 (
            .O(N__28028),
            .I(N__28019));
    InMux I__5002 (
            .O(N__28027),
            .I(N__28019));
    InMux I__5001 (
            .O(N__28024),
            .I(N__28016));
    LocalMux I__5000 (
            .O(N__28019),
            .I(\nx.n2807 ));
    LocalMux I__4999 (
            .O(N__28016),
            .I(\nx.n2807 ));
    CascadeMux I__4998 (
            .O(N__28011),
            .I(\nx.n2987_cascade_ ));
    CascadeMux I__4997 (
            .O(N__28008),
            .I(\nx.n41_cascade_ ));
    InMux I__4996 (
            .O(N__28005),
            .I(N__28002));
    LocalMux I__4995 (
            .O(N__28002),
            .I(\nx.n39_adj_671 ));
    CascadeMux I__4994 (
            .O(N__27999),
            .I(\nx.n50_cascade_ ));
    InMux I__4993 (
            .O(N__27996),
            .I(N__27993));
    LocalMux I__4992 (
            .O(N__27993),
            .I(N__27990));
    Odrv4 I__4991 (
            .O(N__27990),
            .I(\nx.n2877 ));
    InMux I__4990 (
            .O(N__27987),
            .I(N__27984));
    LocalMux I__4989 (
            .O(N__27984),
            .I(N__27981));
    Span4Mux_v I__4988 (
            .O(N__27981),
            .I(N__27978));
    Odrv4 I__4987 (
            .O(N__27978),
            .I(\nx.n2857 ));
    InMux I__4986 (
            .O(N__27975),
            .I(N__27971));
    CascadeMux I__4985 (
            .O(N__27974),
            .I(N__27967));
    LocalMux I__4984 (
            .O(N__27971),
            .I(N__27964));
    CascadeMux I__4983 (
            .O(N__27970),
            .I(N__27961));
    InMux I__4982 (
            .O(N__27967),
            .I(N__27958));
    Span4Mux_h I__4981 (
            .O(N__27964),
            .I(N__27955));
    InMux I__4980 (
            .O(N__27961),
            .I(N__27952));
    LocalMux I__4979 (
            .O(N__27958),
            .I(N__27949));
    Odrv4 I__4978 (
            .O(N__27955),
            .I(\nx.n2790 ));
    LocalMux I__4977 (
            .O(N__27952),
            .I(\nx.n2790 ));
    Odrv12 I__4976 (
            .O(N__27949),
            .I(\nx.n2790 ));
    CascadeMux I__4975 (
            .O(N__27942),
            .I(\nx.n2889_cascade_ ));
    InMux I__4974 (
            .O(N__27939),
            .I(N__27936));
    LocalMux I__4973 (
            .O(N__27936),
            .I(N__27933));
    Odrv4 I__4972 (
            .O(N__27933),
            .I(\nx.n2868 ));
    CascadeMux I__4971 (
            .O(N__27930),
            .I(\nx.n12811_cascade_ ));
    CascadeMux I__4970 (
            .O(N__27927),
            .I(\nx.n12813_cascade_ ));
    InMux I__4969 (
            .O(N__27924),
            .I(N__27921));
    LocalMux I__4968 (
            .O(N__27921),
            .I(\nx.n12815 ));
    InMux I__4967 (
            .O(N__27918),
            .I(N__27915));
    LocalMux I__4966 (
            .O(N__27915),
            .I(\nx.n43_adj_753 ));
    CascadeMux I__4965 (
            .O(N__27912),
            .I(\nx.n46_cascade_ ));
    CascadeMux I__4964 (
            .O(N__27909),
            .I(\nx.n13_adj_743_cascade_ ));
    InMux I__4963 (
            .O(N__27906),
            .I(N__27903));
    LocalMux I__4962 (
            .O(N__27903),
            .I(\nx.n12775 ));
    CascadeMux I__4961 (
            .O(N__27900),
            .I(\nx.n12787_cascade_ ));
    InMux I__4960 (
            .O(N__27897),
            .I(N__27894));
    LocalMux I__4959 (
            .O(N__27894),
            .I(\nx.n12803 ));
    InMux I__4958 (
            .O(N__27891),
            .I(N__27888));
    LocalMux I__4957 (
            .O(N__27888),
            .I(\nx.n35_adj_738 ));
    InMux I__4956 (
            .O(N__27885),
            .I(N__27879));
    InMux I__4955 (
            .O(N__27884),
            .I(N__27879));
    LocalMux I__4954 (
            .O(N__27879),
            .I(N__27875));
    InMux I__4953 (
            .O(N__27878),
            .I(N__27872));
    Odrv4 I__4952 (
            .O(N__27875),
            .I(blink_counter_21));
    LocalMux I__4951 (
            .O(N__27872),
            .I(blink_counter_21));
    InMux I__4950 (
            .O(N__27867),
            .I(n10664));
    InMux I__4949 (
            .O(N__27864),
            .I(N__27858));
    InMux I__4948 (
            .O(N__27863),
            .I(N__27858));
    LocalMux I__4947 (
            .O(N__27858),
            .I(N__27854));
    InMux I__4946 (
            .O(N__27857),
            .I(N__27851));
    Odrv12 I__4945 (
            .O(N__27854),
            .I(blink_counter_22));
    LocalMux I__4944 (
            .O(N__27851),
            .I(blink_counter_22));
    InMux I__4943 (
            .O(N__27846),
            .I(n10665));
    CascadeMux I__4942 (
            .O(N__27843),
            .I(N__27839));
    InMux I__4941 (
            .O(N__27842),
            .I(N__27834));
    InMux I__4940 (
            .O(N__27839),
            .I(N__27834));
    LocalMux I__4939 (
            .O(N__27834),
            .I(N__27830));
    InMux I__4938 (
            .O(N__27833),
            .I(N__27827));
    Odrv4 I__4937 (
            .O(N__27830),
            .I(blink_counter_23));
    LocalMux I__4936 (
            .O(N__27827),
            .I(blink_counter_23));
    InMux I__4935 (
            .O(N__27822),
            .I(n10666));
    CascadeMux I__4934 (
            .O(N__27819),
            .I(N__27816));
    InMux I__4933 (
            .O(N__27816),
            .I(N__27810));
    InMux I__4932 (
            .O(N__27815),
            .I(N__27810));
    LocalMux I__4931 (
            .O(N__27810),
            .I(N__27807));
    Span4Mux_v I__4930 (
            .O(N__27807),
            .I(N__27803));
    InMux I__4929 (
            .O(N__27806),
            .I(N__27800));
    Odrv4 I__4928 (
            .O(N__27803),
            .I(blink_counter_24));
    LocalMux I__4927 (
            .O(N__27800),
            .I(blink_counter_24));
    InMux I__4926 (
            .O(N__27795),
            .I(bfn_9_32_0_));
    InMux I__4925 (
            .O(N__27792),
            .I(n10668));
    InMux I__4924 (
            .O(N__27789),
            .I(N__27786));
    LocalMux I__4923 (
            .O(N__27786),
            .I(N__27783));
    Span4Mux_v I__4922 (
            .O(N__27783),
            .I(N__27779));
    InMux I__4921 (
            .O(N__27782),
            .I(N__27776));
    Odrv4 I__4920 (
            .O(N__27779),
            .I(blink_counter_25));
    LocalMux I__4919 (
            .O(N__27776),
            .I(blink_counter_25));
    CascadeMux I__4918 (
            .O(N__27771),
            .I(\nx.n45_adj_754_cascade_ ));
    CascadeMux I__4917 (
            .O(N__27768),
            .I(\nx.n12809_cascade_ ));
    InMux I__4916 (
            .O(N__27765),
            .I(N__27762));
    LocalMux I__4915 (
            .O(N__27762),
            .I(n13));
    InMux I__4914 (
            .O(N__27759),
            .I(n10656));
    InMux I__4913 (
            .O(N__27756),
            .I(N__27753));
    LocalMux I__4912 (
            .O(N__27753),
            .I(n12));
    InMux I__4911 (
            .O(N__27750),
            .I(n10657));
    InMux I__4910 (
            .O(N__27747),
            .I(N__27744));
    LocalMux I__4909 (
            .O(N__27744),
            .I(n11));
    InMux I__4908 (
            .O(N__27741),
            .I(n10658));
    InMux I__4907 (
            .O(N__27738),
            .I(N__27735));
    LocalMux I__4906 (
            .O(N__27735),
            .I(n10_adj_806));
    InMux I__4905 (
            .O(N__27732),
            .I(bfn_9_31_0_));
    InMux I__4904 (
            .O(N__27729),
            .I(N__27726));
    LocalMux I__4903 (
            .O(N__27726),
            .I(n9_adj_807));
    InMux I__4902 (
            .O(N__27723),
            .I(n10660));
    InMux I__4901 (
            .O(N__27720),
            .I(N__27717));
    LocalMux I__4900 (
            .O(N__27717),
            .I(n8));
    InMux I__4899 (
            .O(N__27714),
            .I(n10661));
    InMux I__4898 (
            .O(N__27711),
            .I(N__27708));
    LocalMux I__4897 (
            .O(N__27708),
            .I(n7_adj_808));
    InMux I__4896 (
            .O(N__27705),
            .I(n10662));
    InMux I__4895 (
            .O(N__27702),
            .I(N__27699));
    LocalMux I__4894 (
            .O(N__27699),
            .I(n6_adj_809));
    InMux I__4893 (
            .O(N__27696),
            .I(n10663));
    InMux I__4892 (
            .O(N__27693),
            .I(N__27690));
    LocalMux I__4891 (
            .O(N__27690),
            .I(n21));
    InMux I__4890 (
            .O(N__27687),
            .I(n10648));
    InMux I__4889 (
            .O(N__27684),
            .I(N__27681));
    LocalMux I__4888 (
            .O(N__27681),
            .I(n20));
    InMux I__4887 (
            .O(N__27678),
            .I(n10649));
    InMux I__4886 (
            .O(N__27675),
            .I(N__27672));
    LocalMux I__4885 (
            .O(N__27672),
            .I(n19_adj_800));
    InMux I__4884 (
            .O(N__27669),
            .I(n10650));
    InMux I__4883 (
            .O(N__27666),
            .I(N__27663));
    LocalMux I__4882 (
            .O(N__27663),
            .I(n18));
    InMux I__4881 (
            .O(N__27660),
            .I(bfn_9_30_0_));
    InMux I__4880 (
            .O(N__27657),
            .I(N__27654));
    LocalMux I__4879 (
            .O(N__27654),
            .I(n17));
    InMux I__4878 (
            .O(N__27651),
            .I(n10652));
    InMux I__4877 (
            .O(N__27648),
            .I(N__27645));
    LocalMux I__4876 (
            .O(N__27645),
            .I(n16));
    InMux I__4875 (
            .O(N__27642),
            .I(n10653));
    InMux I__4874 (
            .O(N__27639),
            .I(N__27636));
    LocalMux I__4873 (
            .O(N__27636),
            .I(n15));
    InMux I__4872 (
            .O(N__27633),
            .I(n10654));
    InMux I__4871 (
            .O(N__27630),
            .I(N__27627));
    LocalMux I__4870 (
            .O(N__27627),
            .I(n14_adj_802));
    InMux I__4869 (
            .O(N__27624),
            .I(n10655));
    InMux I__4868 (
            .O(N__27621),
            .I(N__27618));
    LocalMux I__4867 (
            .O(N__27618),
            .I(N__27615));
    Odrv4 I__4866 (
            .O(N__27615),
            .I(\nx.n1969 ));
    CascadeMux I__4865 (
            .O(N__27612),
            .I(N__27609));
    InMux I__4864 (
            .O(N__27609),
            .I(N__27606));
    LocalMux I__4863 (
            .O(N__27606),
            .I(N__27602));
    CascadeMux I__4862 (
            .O(N__27605),
            .I(N__27598));
    Span4Mux_h I__4861 (
            .O(N__27602),
            .I(N__27595));
    InMux I__4860 (
            .O(N__27601),
            .I(N__27592));
    InMux I__4859 (
            .O(N__27598),
            .I(N__27589));
    Odrv4 I__4858 (
            .O(N__27595),
            .I(\nx.n1902 ));
    LocalMux I__4857 (
            .O(N__27592),
            .I(\nx.n1902 ));
    LocalMux I__4856 (
            .O(N__27589),
            .I(\nx.n1902 ));
    CascadeMux I__4855 (
            .O(N__27582),
            .I(N__27577));
    CascadeMux I__4854 (
            .O(N__27581),
            .I(N__27573));
    CascadeMux I__4853 (
            .O(N__27580),
            .I(N__27569));
    InMux I__4852 (
            .O(N__27577),
            .I(N__27558));
    InMux I__4851 (
            .O(N__27576),
            .I(N__27558));
    InMux I__4850 (
            .O(N__27573),
            .I(N__27558));
    InMux I__4849 (
            .O(N__27572),
            .I(N__27558));
    InMux I__4848 (
            .O(N__27569),
            .I(N__27553));
    InMux I__4847 (
            .O(N__27568),
            .I(N__27553));
    CascadeMux I__4846 (
            .O(N__27567),
            .I(N__27547));
    LocalMux I__4845 (
            .O(N__27558),
            .I(N__27540));
    LocalMux I__4844 (
            .O(N__27553),
            .I(N__27537));
    InMux I__4843 (
            .O(N__27552),
            .I(N__27534));
    InMux I__4842 (
            .O(N__27551),
            .I(N__27525));
    InMux I__4841 (
            .O(N__27550),
            .I(N__27525));
    InMux I__4840 (
            .O(N__27547),
            .I(N__27525));
    InMux I__4839 (
            .O(N__27546),
            .I(N__27525));
    CascadeMux I__4838 (
            .O(N__27545),
            .I(N__27522));
    CascadeMux I__4837 (
            .O(N__27544),
            .I(N__27519));
    InMux I__4836 (
            .O(N__27543),
            .I(N__27515));
    Span4Mux_v I__4835 (
            .O(N__27540),
            .I(N__27510));
    Span4Mux_v I__4834 (
            .O(N__27537),
            .I(N__27510));
    LocalMux I__4833 (
            .O(N__27534),
            .I(N__27505));
    LocalMux I__4832 (
            .O(N__27525),
            .I(N__27505));
    InMux I__4831 (
            .O(N__27522),
            .I(N__27498));
    InMux I__4830 (
            .O(N__27519),
            .I(N__27498));
    InMux I__4829 (
            .O(N__27518),
            .I(N__27498));
    LocalMux I__4828 (
            .O(N__27515),
            .I(\nx.n1928 ));
    Odrv4 I__4827 (
            .O(N__27510),
            .I(\nx.n1928 ));
    Odrv4 I__4826 (
            .O(N__27505),
            .I(\nx.n1928 ));
    LocalMux I__4825 (
            .O(N__27498),
            .I(\nx.n1928 ));
    InMux I__4824 (
            .O(N__27489),
            .I(N__27486));
    LocalMux I__4823 (
            .O(N__27486),
            .I(\nx.n2068 ));
    CascadeMux I__4822 (
            .O(N__27483),
            .I(\nx.n2001_cascade_ ));
    InMux I__4821 (
            .O(N__27480),
            .I(N__27477));
    LocalMux I__4820 (
            .O(N__27477),
            .I(\nx.n2067 ));
    CascadeMux I__4819 (
            .O(N__27474),
            .I(\nx.n2099_cascade_ ));
    InMux I__4818 (
            .O(N__27471),
            .I(N__27468));
    LocalMux I__4817 (
            .O(N__27468),
            .I(n26_adj_798));
    InMux I__4816 (
            .O(N__27465),
            .I(bfn_9_29_0_));
    InMux I__4815 (
            .O(N__27462),
            .I(N__27459));
    LocalMux I__4814 (
            .O(N__27459),
            .I(n25));
    InMux I__4813 (
            .O(N__27456),
            .I(n10644));
    InMux I__4812 (
            .O(N__27453),
            .I(N__27450));
    LocalMux I__4811 (
            .O(N__27450),
            .I(n24));
    InMux I__4810 (
            .O(N__27447),
            .I(n10645));
    InMux I__4809 (
            .O(N__27444),
            .I(N__27441));
    LocalMux I__4808 (
            .O(N__27441),
            .I(n23));
    InMux I__4807 (
            .O(N__27438),
            .I(n10646));
    InMux I__4806 (
            .O(N__27435),
            .I(N__27432));
    LocalMux I__4805 (
            .O(N__27432),
            .I(n22_adj_799));
    InMux I__4804 (
            .O(N__27429),
            .I(n10647));
    InMux I__4803 (
            .O(N__27426),
            .I(\nx.n10858 ));
    InMux I__4802 (
            .O(N__27423),
            .I(\nx.n10859 ));
    InMux I__4801 (
            .O(N__27420),
            .I(\nx.n10860 ));
    InMux I__4800 (
            .O(N__27417),
            .I(\nx.n10861 ));
    InMux I__4799 (
            .O(N__27414),
            .I(\nx.n10862 ));
    InMux I__4798 (
            .O(N__27411),
            .I(N__27408));
    LocalMux I__4797 (
            .O(N__27408),
            .I(N__27404));
    InMux I__4796 (
            .O(N__27407),
            .I(N__27401));
    Odrv4 I__4795 (
            .O(N__27404),
            .I(\nx.n1994 ));
    LocalMux I__4794 (
            .O(N__27401),
            .I(\nx.n1994 ));
    InMux I__4793 (
            .O(N__27396),
            .I(bfn_9_28_0_));
    CascadeMux I__4792 (
            .O(N__27393),
            .I(N__27389));
    CascadeMux I__4791 (
            .O(N__27392),
            .I(N__27386));
    InMux I__4790 (
            .O(N__27389),
            .I(N__27383));
    InMux I__4789 (
            .O(N__27386),
            .I(N__27380));
    LocalMux I__4788 (
            .O(N__27383),
            .I(N__27375));
    LocalMux I__4787 (
            .O(N__27380),
            .I(N__27375));
    Span4Mux_v I__4786 (
            .O(N__27375),
            .I(N__27372));
    Span4Mux_h I__4785 (
            .O(N__27372),
            .I(N__27369));
    Odrv4 I__4784 (
            .O(N__27369),
            .I(\nx.n1995 ));
    InMux I__4783 (
            .O(N__27366),
            .I(N__27363));
    LocalMux I__4782 (
            .O(N__27363),
            .I(\nx.n2062 ));
    CascadeMux I__4781 (
            .O(N__27360),
            .I(\nx.n2094_cascade_ ));
    InMux I__4780 (
            .O(N__27357),
            .I(N__27352));
    CascadeMux I__4779 (
            .O(N__27356),
            .I(N__27349));
    InMux I__4778 (
            .O(N__27355),
            .I(N__27346));
    LocalMux I__4777 (
            .O(N__27352),
            .I(N__27343));
    InMux I__4776 (
            .O(N__27349),
            .I(N__27340));
    LocalMux I__4775 (
            .O(N__27346),
            .I(N__27337));
    Odrv4 I__4774 (
            .O(N__27343),
            .I(\nx.n1901 ));
    LocalMux I__4773 (
            .O(N__27340),
            .I(\nx.n1901 ));
    Odrv4 I__4772 (
            .O(N__27337),
            .I(\nx.n1901 ));
    InMux I__4771 (
            .O(N__27330),
            .I(N__27327));
    LocalMux I__4770 (
            .O(N__27327),
            .I(N__27324));
    Odrv4 I__4769 (
            .O(N__27324),
            .I(\nx.n1968 ));
    InMux I__4768 (
            .O(N__27321),
            .I(\nx.n10849 ));
    InMux I__4767 (
            .O(N__27318),
            .I(\nx.n10850 ));
    InMux I__4766 (
            .O(N__27315),
            .I(\nx.n10851 ));
    InMux I__4765 (
            .O(N__27312),
            .I(\nx.n10852 ));
    InMux I__4764 (
            .O(N__27309),
            .I(\nx.n10853 ));
    InMux I__4763 (
            .O(N__27306),
            .I(\nx.n10854 ));
    InMux I__4762 (
            .O(N__27303),
            .I(bfn_9_27_0_));
    InMux I__4761 (
            .O(N__27300),
            .I(\nx.n10856 ));
    InMux I__4760 (
            .O(N__27297),
            .I(\nx.n10857 ));
    InMux I__4759 (
            .O(N__27294),
            .I(N__27290));
    InMux I__4758 (
            .O(N__27293),
            .I(N__27286));
    LocalMux I__4757 (
            .O(N__27290),
            .I(N__27283));
    InMux I__4756 (
            .O(N__27289),
            .I(N__27280));
    LocalMux I__4755 (
            .O(N__27286),
            .I(N__27275));
    Span4Mux_v I__4754 (
            .O(N__27283),
            .I(N__27275));
    LocalMux I__4753 (
            .O(N__27280),
            .I(N__27272));
    Span4Mux_v I__4752 (
            .O(N__27275),
            .I(N__27267));
    Span4Mux_h I__4751 (
            .O(N__27272),
            .I(N__27264));
    InMux I__4750 (
            .O(N__27271),
            .I(N__27261));
    InMux I__4749 (
            .O(N__27270),
            .I(N__27258));
    Span4Mux_h I__4748 (
            .O(N__27267),
            .I(N__27255));
    Span4Mux_v I__4747 (
            .O(N__27264),
            .I(N__27252));
    LocalMux I__4746 (
            .O(N__27261),
            .I(neopxl_color_5));
    LocalMux I__4745 (
            .O(N__27258),
            .I(neopxl_color_5));
    Odrv4 I__4744 (
            .O(N__27255),
            .I(neopxl_color_5));
    Odrv4 I__4743 (
            .O(N__27252),
            .I(neopxl_color_5));
    SRMux I__4742 (
            .O(N__27243),
            .I(N__27240));
    LocalMux I__4741 (
            .O(N__27240),
            .I(N__27237));
    Span4Mux_v I__4740 (
            .O(N__27237),
            .I(N__27234));
    Sp12to4 I__4739 (
            .O(N__27234),
            .I(N__27231));
    Odrv12 I__4738 (
            .O(N__27231),
            .I(n22));
    InMux I__4737 (
            .O(N__27228),
            .I(N__27225));
    LocalMux I__4736 (
            .O(N__27225),
            .I(N__27222));
    Span4Mux_h I__4735 (
            .O(N__27222),
            .I(N__27219));
    Odrv4 I__4734 (
            .O(N__27219),
            .I(\nx.n1966 ));
    InMux I__4733 (
            .O(N__27216),
            .I(N__27213));
    LocalMux I__4732 (
            .O(N__27213),
            .I(N__27209));
    CascadeMux I__4731 (
            .O(N__27212),
            .I(N__27206));
    Span4Mux_h I__4730 (
            .O(N__27209),
            .I(N__27202));
    InMux I__4729 (
            .O(N__27206),
            .I(N__27199));
    InMux I__4728 (
            .O(N__27205),
            .I(N__27196));
    Odrv4 I__4727 (
            .O(N__27202),
            .I(\nx.n1899 ));
    LocalMux I__4726 (
            .O(N__27199),
            .I(\nx.n1899 ));
    LocalMux I__4725 (
            .O(N__27196),
            .I(\nx.n1899 ));
    InMux I__4724 (
            .O(N__27189),
            .I(N__27186));
    LocalMux I__4723 (
            .O(N__27186),
            .I(N__27183));
    Span4Mux_h I__4722 (
            .O(N__27183),
            .I(N__27180));
    Odrv4 I__4721 (
            .O(N__27180),
            .I(\nx.n1967 ));
    CascadeMux I__4720 (
            .O(N__27177),
            .I(N__27174));
    InMux I__4719 (
            .O(N__27174),
            .I(N__27171));
    LocalMux I__4718 (
            .O(N__27171),
            .I(N__27167));
    CascadeMux I__4717 (
            .O(N__27170),
            .I(N__27164));
    Span4Mux_h I__4716 (
            .O(N__27167),
            .I(N__27160));
    InMux I__4715 (
            .O(N__27164),
            .I(N__27157));
    InMux I__4714 (
            .O(N__27163),
            .I(N__27154));
    Odrv4 I__4713 (
            .O(N__27160),
            .I(\nx.n1900 ));
    LocalMux I__4712 (
            .O(N__27157),
            .I(\nx.n1900 ));
    LocalMux I__4711 (
            .O(N__27154),
            .I(\nx.n1900 ));
    InMux I__4710 (
            .O(N__27147),
            .I(N__27144));
    LocalMux I__4709 (
            .O(N__27144),
            .I(N__27141));
    Span4Mux_h I__4708 (
            .O(N__27141),
            .I(N__27138));
    Odrv4 I__4707 (
            .O(N__27138),
            .I(\nx.n1970 ));
    InMux I__4706 (
            .O(N__27135),
            .I(N__27132));
    LocalMux I__4705 (
            .O(N__27132),
            .I(N__27128));
    CascadeMux I__4704 (
            .O(N__27131),
            .I(N__27124));
    Span4Mux_h I__4703 (
            .O(N__27128),
            .I(N__27121));
    InMux I__4702 (
            .O(N__27127),
            .I(N__27118));
    InMux I__4701 (
            .O(N__27124),
            .I(N__27115));
    Odrv4 I__4700 (
            .O(N__27121),
            .I(\nx.n1903 ));
    LocalMux I__4699 (
            .O(N__27118),
            .I(\nx.n1903 ));
    LocalMux I__4698 (
            .O(N__27115),
            .I(\nx.n1903 ));
    InMux I__4697 (
            .O(N__27108),
            .I(N__27105));
    LocalMux I__4696 (
            .O(N__27105),
            .I(N__27102));
    Span4Mux_h I__4695 (
            .O(N__27102),
            .I(N__27099));
    Odrv4 I__4694 (
            .O(N__27099),
            .I(\nx.n1972 ));
    CascadeMux I__4693 (
            .O(N__27096),
            .I(N__27093));
    InMux I__4692 (
            .O(N__27093),
            .I(N__27090));
    LocalMux I__4691 (
            .O(N__27090),
            .I(N__27085));
    CascadeMux I__4690 (
            .O(N__27089),
            .I(N__27082));
    CascadeMux I__4689 (
            .O(N__27088),
            .I(N__27079));
    Span4Mux_h I__4688 (
            .O(N__27085),
            .I(N__27076));
    InMux I__4687 (
            .O(N__27082),
            .I(N__27073));
    InMux I__4686 (
            .O(N__27079),
            .I(N__27070));
    Odrv4 I__4685 (
            .O(N__27076),
            .I(\nx.n1905 ));
    LocalMux I__4684 (
            .O(N__27073),
            .I(\nx.n1905 ));
    LocalMux I__4683 (
            .O(N__27070),
            .I(\nx.n1905 ));
    InMux I__4682 (
            .O(N__27063),
            .I(bfn_9_26_0_));
    InMux I__4681 (
            .O(N__27060),
            .I(\nx.n10848 ));
    InMux I__4680 (
            .O(N__27057),
            .I(\nx.n11025 ));
    InMux I__4679 (
            .O(N__27054),
            .I(\nx.n11026 ));
    InMux I__4678 (
            .O(N__27051),
            .I(bfn_9_24_0_));
    CascadeMux I__4677 (
            .O(N__27048),
            .I(N__27043));
    InMux I__4676 (
            .O(N__27047),
            .I(N__27038));
    InMux I__4675 (
            .O(N__27046),
            .I(N__27038));
    InMux I__4674 (
            .O(N__27043),
            .I(N__27035));
    LocalMux I__4673 (
            .O(N__27038),
            .I(N__27032));
    LocalMux I__4672 (
            .O(N__27035),
            .I(\nx.n2792 ));
    Odrv12 I__4671 (
            .O(N__27032),
            .I(\nx.n2792 ));
    InMux I__4670 (
            .O(N__27027),
            .I(N__27024));
    LocalMux I__4669 (
            .O(N__27024),
            .I(N__27021));
    Span12Mux_v I__4668 (
            .O(N__27021),
            .I(N__27018));
    Odrv12 I__4667 (
            .O(N__27018),
            .I(neopxl_color_prev_5));
    InMux I__4666 (
            .O(N__27015),
            .I(\nx.n11016 ));
    InMux I__4665 (
            .O(N__27012),
            .I(\nx.n11017 ));
    InMux I__4664 (
            .O(N__27009),
            .I(\nx.n11018 ));
    InMux I__4663 (
            .O(N__27006),
            .I(bfn_9_23_0_));
    InMux I__4662 (
            .O(N__27003),
            .I(\nx.n11020 ));
    InMux I__4661 (
            .O(N__27000),
            .I(N__26997));
    LocalMux I__4660 (
            .O(N__26997),
            .I(N__26994));
    Odrv4 I__4659 (
            .O(N__26994),
            .I(\nx.n2859 ));
    InMux I__4658 (
            .O(N__26991),
            .I(\nx.n11021 ));
    CascadeMux I__4657 (
            .O(N__26988),
            .I(N__26985));
    InMux I__4656 (
            .O(N__26985),
            .I(N__26982));
    LocalMux I__4655 (
            .O(N__26982),
            .I(N__26978));
    InMux I__4654 (
            .O(N__26981),
            .I(N__26975));
    Odrv4 I__4653 (
            .O(N__26978),
            .I(\nx.n2791 ));
    LocalMux I__4652 (
            .O(N__26975),
            .I(\nx.n2791 ));
    InMux I__4651 (
            .O(N__26970),
            .I(N__26967));
    LocalMux I__4650 (
            .O(N__26967),
            .I(N__26964));
    Odrv4 I__4649 (
            .O(N__26964),
            .I(\nx.n2858 ));
    InMux I__4648 (
            .O(N__26961),
            .I(\nx.n11022 ));
    InMux I__4647 (
            .O(N__26958),
            .I(\nx.n11023 ));
    InMux I__4646 (
            .O(N__26955),
            .I(N__26952));
    LocalMux I__4645 (
            .O(N__26952),
            .I(N__26949));
    Odrv4 I__4644 (
            .O(N__26949),
            .I(\nx.n2856 ));
    InMux I__4643 (
            .O(N__26946),
            .I(\nx.n11024 ));
    InMux I__4642 (
            .O(N__26943),
            .I(\nx.n11007 ));
    InMux I__4641 (
            .O(N__26940),
            .I(\nx.n11008 ));
    InMux I__4640 (
            .O(N__26937),
            .I(\nx.n11009 ));
    InMux I__4639 (
            .O(N__26934),
            .I(\nx.n11010 ));
    InMux I__4638 (
            .O(N__26931),
            .I(bfn_9_22_0_));
    InMux I__4637 (
            .O(N__26928),
            .I(\nx.n11012 ));
    InMux I__4636 (
            .O(N__26925),
            .I(\nx.n11013 ));
    InMux I__4635 (
            .O(N__26922),
            .I(\nx.n11014 ));
    InMux I__4634 (
            .O(N__26919),
            .I(\nx.n11015 ));
    CascadeMux I__4633 (
            .O(N__26916),
            .I(\nx.n2791_cascade_ ));
    InMux I__4632 (
            .O(N__26913),
            .I(bfn_9_21_0_));
    CascadeMux I__4631 (
            .O(N__26910),
            .I(N__26907));
    InMux I__4630 (
            .O(N__26907),
            .I(N__26904));
    LocalMux I__4629 (
            .O(N__26904),
            .I(N__26901));
    Odrv4 I__4628 (
            .O(N__26901),
            .I(\nx.n2876 ));
    InMux I__4627 (
            .O(N__26898),
            .I(\nx.n11004 ));
    InMux I__4626 (
            .O(N__26895),
            .I(N__26892));
    LocalMux I__4625 (
            .O(N__26892),
            .I(N__26889));
    Odrv4 I__4624 (
            .O(N__26889),
            .I(\nx.n2875 ));
    InMux I__4623 (
            .O(N__26886),
            .I(\nx.n11005 ));
    InMux I__4622 (
            .O(N__26883),
            .I(\nx.n11006 ));
    InMux I__4621 (
            .O(N__26880),
            .I(N__26877));
    LocalMux I__4620 (
            .O(N__26877),
            .I(N__26874));
    Span4Mux_h I__4619 (
            .O(N__26874),
            .I(N__26871));
    Span4Mux_v I__4618 (
            .O(N__26871),
            .I(N__26867));
    InMux I__4617 (
            .O(N__26870),
            .I(N__26864));
    Odrv4 I__4616 (
            .O(N__26867),
            .I(\nx.bit_ctr_2 ));
    LocalMux I__4615 (
            .O(N__26864),
            .I(\nx.bit_ctr_2 ));
    InMux I__4614 (
            .O(N__26859),
            .I(N__26856));
    LocalMux I__4613 (
            .O(N__26856),
            .I(N__26850));
    InMux I__4612 (
            .O(N__26855),
            .I(N__26847));
    InMux I__4611 (
            .O(N__26854),
            .I(N__26844));
    InMux I__4610 (
            .O(N__26853),
            .I(N__26841));
    Span4Mux_v I__4609 (
            .O(N__26850),
            .I(N__26838));
    LocalMux I__4608 (
            .O(N__26847),
            .I(N__26831));
    LocalMux I__4607 (
            .O(N__26844),
            .I(N__26831));
    LocalMux I__4606 (
            .O(N__26841),
            .I(N__26831));
    Span4Mux_h I__4605 (
            .O(N__26838),
            .I(N__26826));
    Span4Mux_v I__4604 (
            .O(N__26831),
            .I(N__26826));
    Odrv4 I__4603 (
            .O(N__26826),
            .I(state_3_N_448_1));
    CascadeMux I__4602 (
            .O(N__26823),
            .I(N__26820));
    InMux I__4601 (
            .O(N__26820),
            .I(N__26817));
    LocalMux I__4600 (
            .O(N__26817),
            .I(\nx.color_bit_N_642_4 ));
    InMux I__4599 (
            .O(N__26814),
            .I(N__26811));
    LocalMux I__4598 (
            .O(N__26811),
            .I(N__26808));
    Odrv4 I__4597 (
            .O(N__26808),
            .I(\nx.n13622 ));
    CascadeMux I__4596 (
            .O(N__26805),
            .I(N__26791));
    CascadeMux I__4595 (
            .O(N__26804),
            .I(N__26788));
    InMux I__4594 (
            .O(N__26803),
            .I(N__26781));
    InMux I__4593 (
            .O(N__26802),
            .I(N__26781));
    InMux I__4592 (
            .O(N__26801),
            .I(N__26781));
    InMux I__4591 (
            .O(N__26800),
            .I(N__26778));
    InMux I__4590 (
            .O(N__26799),
            .I(N__26772));
    InMux I__4589 (
            .O(N__26798),
            .I(N__26772));
    CascadeMux I__4588 (
            .O(N__26797),
            .I(N__26769));
    InMux I__4587 (
            .O(N__26796),
            .I(N__26760));
    InMux I__4586 (
            .O(N__26795),
            .I(N__26760));
    InMux I__4585 (
            .O(N__26794),
            .I(N__26760));
    InMux I__4584 (
            .O(N__26791),
            .I(N__26760));
    InMux I__4583 (
            .O(N__26788),
            .I(N__26757));
    LocalMux I__4582 (
            .O(N__26781),
            .I(N__26754));
    LocalMux I__4581 (
            .O(N__26778),
            .I(N__26751));
    InMux I__4580 (
            .O(N__26777),
            .I(N__26748));
    LocalMux I__4579 (
            .O(N__26772),
            .I(N__26745));
    InMux I__4578 (
            .O(N__26769),
            .I(N__26742));
    LocalMux I__4577 (
            .O(N__26760),
            .I(N__26737));
    LocalMux I__4576 (
            .O(N__26757),
            .I(N__26737));
    Span4Mux_v I__4575 (
            .O(N__26754),
            .I(N__26732));
    Span4Mux_h I__4574 (
            .O(N__26751),
            .I(N__26732));
    LocalMux I__4573 (
            .O(N__26748),
            .I(N__26725));
    Span4Mux_v I__4572 (
            .O(N__26745),
            .I(N__26725));
    LocalMux I__4571 (
            .O(N__26742),
            .I(N__26725));
    Span4Mux_h I__4570 (
            .O(N__26737),
            .I(N__26720));
    Span4Mux_h I__4569 (
            .O(N__26732),
            .I(N__26720));
    Odrv4 I__4568 (
            .O(N__26725),
            .I(state_0_adj_792));
    Odrv4 I__4567 (
            .O(N__26720),
            .I(state_0_adj_792));
    CEMux I__4566 (
            .O(N__26715),
            .I(N__26712));
    LocalMux I__4565 (
            .O(N__26712),
            .I(N__26709));
    Span4Mux_h I__4564 (
            .O(N__26709),
            .I(N__26705));
    InMux I__4563 (
            .O(N__26708),
            .I(N__26702));
    Odrv4 I__4562 (
            .O(N__26705),
            .I(n7671));
    LocalMux I__4561 (
            .O(N__26702),
            .I(n7671));
    SRMux I__4560 (
            .O(N__26697),
            .I(N__26694));
    LocalMux I__4559 (
            .O(N__26694),
            .I(N__26691));
    Odrv4 I__4558 (
            .O(N__26691),
            .I(\nx.n7983 ));
    CascadeMux I__4557 (
            .O(N__26688),
            .I(N__26685));
    InMux I__4556 (
            .O(N__26685),
            .I(N__26682));
    LocalMux I__4555 (
            .O(N__26682),
            .I(\nx.n12817 ));
    CascadeMux I__4554 (
            .O(N__26679),
            .I(\nx.n12819_cascade_ ));
    InMux I__4553 (
            .O(N__26676),
            .I(N__26673));
    LocalMux I__4552 (
            .O(N__26673),
            .I(\nx.n12821 ));
    CascadeMux I__4551 (
            .O(N__26670),
            .I(\nx.n3009_cascade_ ));
    InMux I__4550 (
            .O(N__26667),
            .I(N__26664));
    LocalMux I__4549 (
            .O(N__26664),
            .I(N__26661));
    Odrv12 I__4548 (
            .O(N__26661),
            .I(\nx.n1971 ));
    CascadeMux I__4547 (
            .O(N__26658),
            .I(N__26655));
    InMux I__4546 (
            .O(N__26655),
            .I(N__26650));
    CascadeMux I__4545 (
            .O(N__26654),
            .I(N__26647));
    InMux I__4544 (
            .O(N__26653),
            .I(N__26644));
    LocalMux I__4543 (
            .O(N__26650),
            .I(N__26641));
    InMux I__4542 (
            .O(N__26647),
            .I(N__26638));
    LocalMux I__4541 (
            .O(N__26644),
            .I(N__26635));
    Odrv4 I__4540 (
            .O(N__26641),
            .I(\nx.n1904 ));
    LocalMux I__4539 (
            .O(N__26638),
            .I(\nx.n1904 ));
    Odrv4 I__4538 (
            .O(N__26635),
            .I(\nx.n1904 ));
    InMux I__4537 (
            .O(N__26628),
            .I(N__26625));
    LocalMux I__4536 (
            .O(N__26625),
            .I(n13360));
    CascadeMux I__4535 (
            .O(N__26622),
            .I(n13361_cascade_));
    IoInMux I__4534 (
            .O(N__26619),
            .I(N__26616));
    LocalMux I__4533 (
            .O(N__26616),
            .I(N__26613));
    Span12Mux_s1_v I__4532 (
            .O(N__26613),
            .I(N__26610));
    Odrv12 I__4531 (
            .O(N__26610),
            .I(LED_c));
    InMux I__4530 (
            .O(N__26607),
            .I(N__26600));
    InMux I__4529 (
            .O(N__26606),
            .I(N__26600));
    InMux I__4528 (
            .O(N__26605),
            .I(N__26597));
    LocalMux I__4527 (
            .O(N__26600),
            .I(N__26593));
    LocalMux I__4526 (
            .O(N__26597),
            .I(N__26590));
    InMux I__4525 (
            .O(N__26596),
            .I(N__26587));
    Span12Mux_s8_h I__4524 (
            .O(N__26593),
            .I(N__26584));
    Span4Mux_h I__4523 (
            .O(N__26590),
            .I(N__26581));
    LocalMux I__4522 (
            .O(N__26587),
            .I(neopxl_color_12));
    Odrv12 I__4521 (
            .O(N__26584),
            .I(neopxl_color_12));
    Odrv4 I__4520 (
            .O(N__26581),
            .I(neopxl_color_12));
    InMux I__4519 (
            .O(N__26574),
            .I(N__26571));
    LocalMux I__4518 (
            .O(N__26571),
            .I(\nx.n59 ));
    CascadeMux I__4517 (
            .O(N__26568),
            .I(\nx.n61_cascade_ ));
    InMux I__4516 (
            .O(N__26565),
            .I(N__26561));
    InMux I__4515 (
            .O(N__26564),
            .I(N__26558));
    LocalMux I__4514 (
            .O(N__26561),
            .I(N__26555));
    LocalMux I__4513 (
            .O(N__26558),
            .I(\nx.n11153 ));
    Odrv4 I__4512 (
            .O(N__26555),
            .I(\nx.n11153 ));
    InMux I__4511 (
            .O(N__26550),
            .I(\nx.n10845 ));
    InMux I__4510 (
            .O(N__26547),
            .I(\nx.n10846 ));
    CascadeMux I__4509 (
            .O(N__26544),
            .I(N__26540));
    InMux I__4508 (
            .O(N__26543),
            .I(N__26537));
    InMux I__4507 (
            .O(N__26540),
            .I(N__26534));
    LocalMux I__4506 (
            .O(N__26537),
            .I(N__26531));
    LocalMux I__4505 (
            .O(N__26534),
            .I(\nx.n1895 ));
    Odrv4 I__4504 (
            .O(N__26531),
            .I(\nx.n1895 ));
    InMux I__4503 (
            .O(N__26526),
            .I(\nx.n10847 ));
    InMux I__4502 (
            .O(N__26523),
            .I(N__26520));
    LocalMux I__4501 (
            .O(N__26520),
            .I(N__26517));
    Odrv4 I__4500 (
            .O(N__26517),
            .I(\nx.n24 ));
    CascadeMux I__4499 (
            .O(N__26514),
            .I(N__26511));
    InMux I__4498 (
            .O(N__26511),
            .I(N__26508));
    LocalMux I__4497 (
            .O(N__26508),
            .I(\nx.n1963 ));
    CascadeMux I__4496 (
            .O(N__26505),
            .I(N__26501));
    CascadeMux I__4495 (
            .O(N__26504),
            .I(N__26497));
    InMux I__4494 (
            .O(N__26501),
            .I(N__26494));
    InMux I__4493 (
            .O(N__26500),
            .I(N__26491));
    InMux I__4492 (
            .O(N__26497),
            .I(N__26488));
    LocalMux I__4491 (
            .O(N__26494),
            .I(N__26485));
    LocalMux I__4490 (
            .O(N__26491),
            .I(\nx.n1896 ));
    LocalMux I__4489 (
            .O(N__26488),
            .I(\nx.n1896 ));
    Odrv4 I__4488 (
            .O(N__26485),
            .I(\nx.n1896 ));
    CascadeMux I__4487 (
            .O(N__26478),
            .I(\nx.n1995_cascade_ ));
    InMux I__4486 (
            .O(N__26475),
            .I(N__26472));
    LocalMux I__4485 (
            .O(N__26472),
            .I(\nx.n1965 ));
    CascadeMux I__4484 (
            .O(N__26469),
            .I(N__26464));
    CascadeMux I__4483 (
            .O(N__26468),
            .I(N__26461));
    CascadeMux I__4482 (
            .O(N__26467),
            .I(N__26458));
    InMux I__4481 (
            .O(N__26464),
            .I(N__26455));
    InMux I__4480 (
            .O(N__26461),
            .I(N__26452));
    InMux I__4479 (
            .O(N__26458),
            .I(N__26449));
    LocalMux I__4478 (
            .O(N__26455),
            .I(\nx.n1898 ));
    LocalMux I__4477 (
            .O(N__26452),
            .I(\nx.n1898 ));
    LocalMux I__4476 (
            .O(N__26449),
            .I(\nx.n1898 ));
    InMux I__4475 (
            .O(N__26442),
            .I(N__26439));
    LocalMux I__4474 (
            .O(N__26439),
            .I(\nx.n1964 ));
    CascadeMux I__4473 (
            .O(N__26436),
            .I(N__26433));
    InMux I__4472 (
            .O(N__26433),
            .I(N__26428));
    InMux I__4471 (
            .O(N__26432),
            .I(N__26423));
    InMux I__4470 (
            .O(N__26431),
            .I(N__26423));
    LocalMux I__4469 (
            .O(N__26428),
            .I(\nx.n1897 ));
    LocalMux I__4468 (
            .O(N__26423),
            .I(\nx.n1897 ));
    CascadeMux I__4467 (
            .O(N__26418),
            .I(N__26413));
    InMux I__4466 (
            .O(N__26417),
            .I(N__26408));
    InMux I__4465 (
            .O(N__26416),
            .I(N__26408));
    InMux I__4464 (
            .O(N__26413),
            .I(N__26405));
    LocalMux I__4463 (
            .O(N__26408),
            .I(\nx.n1906 ));
    LocalMux I__4462 (
            .O(N__26405),
            .I(\nx.n1906 ));
    InMux I__4461 (
            .O(N__26400),
            .I(N__26397));
    LocalMux I__4460 (
            .O(N__26397),
            .I(\nx.n1973 ));
    InMux I__4459 (
            .O(N__26394),
            .I(\nx.n10836 ));
    InMux I__4458 (
            .O(N__26391),
            .I(\nx.n10837 ));
    InMux I__4457 (
            .O(N__26388),
            .I(\nx.n10838 ));
    InMux I__4456 (
            .O(N__26385),
            .I(\nx.n10839 ));
    InMux I__4455 (
            .O(N__26382),
            .I(bfn_7_28_0_));
    InMux I__4454 (
            .O(N__26379),
            .I(\nx.n10841 ));
    InMux I__4453 (
            .O(N__26376),
            .I(\nx.n10842 ));
    InMux I__4452 (
            .O(N__26373),
            .I(\nx.n10843 ));
    InMux I__4451 (
            .O(N__26370),
            .I(\nx.n10844 ));
    CascadeMux I__4450 (
            .O(N__26367),
            .I(\nx.n28_adj_679_cascade_ ));
    InMux I__4449 (
            .O(N__26364),
            .I(N__26361));
    LocalMux I__4448 (
            .O(N__26361),
            .I(\nx.n16_adj_678 ));
    CascadeMux I__4447 (
            .O(N__26358),
            .I(\nx.n1928_cascade_ ));
    InMux I__4446 (
            .O(N__26355),
            .I(N__26350));
    InMux I__4445 (
            .O(N__26354),
            .I(N__26345));
    InMux I__4444 (
            .O(N__26353),
            .I(N__26342));
    LocalMux I__4443 (
            .O(N__26350),
            .I(N__26339));
    InMux I__4442 (
            .O(N__26349),
            .I(N__26334));
    InMux I__4441 (
            .O(N__26348),
            .I(N__26334));
    LocalMux I__4440 (
            .O(N__26345),
            .I(\nx.bit_ctr_16 ));
    LocalMux I__4439 (
            .O(N__26342),
            .I(\nx.bit_ctr_16 ));
    Odrv4 I__4438 (
            .O(N__26339),
            .I(\nx.bit_ctr_16 ));
    LocalMux I__4437 (
            .O(N__26334),
            .I(\nx.bit_ctr_16 ));
    InMux I__4436 (
            .O(N__26325),
            .I(N__26322));
    LocalMux I__4435 (
            .O(N__26322),
            .I(N__26319));
    Odrv4 I__4434 (
            .O(N__26319),
            .I(\nx.n1977 ));
    InMux I__4433 (
            .O(N__26316),
            .I(bfn_7_27_0_));
    CascadeMux I__4432 (
            .O(N__26313),
            .I(N__26310));
    InMux I__4431 (
            .O(N__26310),
            .I(N__26305));
    CascadeMux I__4430 (
            .O(N__26309),
            .I(N__26302));
    InMux I__4429 (
            .O(N__26308),
            .I(N__26299));
    LocalMux I__4428 (
            .O(N__26305),
            .I(N__26296));
    InMux I__4427 (
            .O(N__26302),
            .I(N__26293));
    LocalMux I__4426 (
            .O(N__26299),
            .I(\nx.n1909 ));
    Odrv4 I__4425 (
            .O(N__26296),
            .I(\nx.n1909 ));
    LocalMux I__4424 (
            .O(N__26293),
            .I(\nx.n1909 ));
    InMux I__4423 (
            .O(N__26286),
            .I(N__26283));
    LocalMux I__4422 (
            .O(N__26283),
            .I(\nx.n1976 ));
    InMux I__4421 (
            .O(N__26280),
            .I(\nx.n10833 ));
    CascadeMux I__4420 (
            .O(N__26277),
            .I(N__26272));
    InMux I__4419 (
            .O(N__26276),
            .I(N__26267));
    InMux I__4418 (
            .O(N__26275),
            .I(N__26267));
    InMux I__4417 (
            .O(N__26272),
            .I(N__26264));
    LocalMux I__4416 (
            .O(N__26267),
            .I(\nx.n1908 ));
    LocalMux I__4415 (
            .O(N__26264),
            .I(\nx.n1908 ));
    InMux I__4414 (
            .O(N__26259),
            .I(N__26256));
    LocalMux I__4413 (
            .O(N__26256),
            .I(\nx.n1975 ));
    InMux I__4412 (
            .O(N__26253),
            .I(\nx.n10834 ));
    CascadeMux I__4411 (
            .O(N__26250),
            .I(N__26245));
    InMux I__4410 (
            .O(N__26249),
            .I(N__26240));
    InMux I__4409 (
            .O(N__26248),
            .I(N__26240));
    InMux I__4408 (
            .O(N__26245),
            .I(N__26237));
    LocalMux I__4407 (
            .O(N__26240),
            .I(\nx.n1907 ));
    LocalMux I__4406 (
            .O(N__26237),
            .I(\nx.n1907 ));
    CascadeMux I__4405 (
            .O(N__26232),
            .I(N__26229));
    InMux I__4404 (
            .O(N__26229),
            .I(N__26226));
    LocalMux I__4403 (
            .O(N__26226),
            .I(\nx.n1974 ));
    InMux I__4402 (
            .O(N__26223),
            .I(\nx.n10835 ));
    CascadeMux I__4401 (
            .O(N__26220),
            .I(N__26216));
    InMux I__4400 (
            .O(N__26219),
            .I(N__26213));
    InMux I__4399 (
            .O(N__26216),
            .I(N__26210));
    LocalMux I__4398 (
            .O(N__26213),
            .I(N__26204));
    LocalMux I__4397 (
            .O(N__26210),
            .I(N__26201));
    InMux I__4396 (
            .O(N__26209),
            .I(N__26198));
    InMux I__4395 (
            .O(N__26208),
            .I(N__26195));
    InMux I__4394 (
            .O(N__26207),
            .I(N__26192));
    Span4Mux_v I__4393 (
            .O(N__26204),
            .I(N__26187));
    Span4Mux_v I__4392 (
            .O(N__26201),
            .I(N__26187));
    LocalMux I__4391 (
            .O(N__26198),
            .I(N__26182));
    LocalMux I__4390 (
            .O(N__26195),
            .I(N__26182));
    LocalMux I__4389 (
            .O(N__26192),
            .I(neopxl_color_6));
    Odrv4 I__4388 (
            .O(N__26187),
            .I(neopxl_color_6));
    Odrv12 I__4387 (
            .O(N__26182),
            .I(neopxl_color_6));
    CascadeMux I__4386 (
            .O(N__26175),
            .I(N__26171));
    InMux I__4385 (
            .O(N__26174),
            .I(N__26167));
    InMux I__4384 (
            .O(N__26171),
            .I(N__26162));
    InMux I__4383 (
            .O(N__26170),
            .I(N__26162));
    LocalMux I__4382 (
            .O(N__26167),
            .I(N__26156));
    LocalMux I__4381 (
            .O(N__26162),
            .I(N__26156));
    InMux I__4380 (
            .O(N__26161),
            .I(N__26152));
    Span4Mux_v I__4379 (
            .O(N__26156),
            .I(N__26149));
    InMux I__4378 (
            .O(N__26155),
            .I(N__26146));
    LocalMux I__4377 (
            .O(N__26152),
            .I(\nx.bit_ctr_0 ));
    Odrv4 I__4376 (
            .O(N__26149),
            .I(\nx.bit_ctr_0 ));
    LocalMux I__4375 (
            .O(N__26146),
            .I(\nx.bit_ctr_0 ));
    InMux I__4374 (
            .O(N__26139),
            .I(N__26136));
    LocalMux I__4373 (
            .O(N__26136),
            .I(N__26133));
    Odrv12 I__4372 (
            .O(N__26133),
            .I(\nx.n13373 ));
    InMux I__4371 (
            .O(N__26130),
            .I(N__26123));
    InMux I__4370 (
            .O(N__26129),
            .I(N__26114));
    InMux I__4369 (
            .O(N__26128),
            .I(N__26114));
    InMux I__4368 (
            .O(N__26127),
            .I(N__26114));
    InMux I__4367 (
            .O(N__26126),
            .I(N__26114));
    LocalMux I__4366 (
            .O(N__26123),
            .I(neopxl_color_7));
    LocalMux I__4365 (
            .O(N__26114),
            .I(neopxl_color_7));
    SRMux I__4364 (
            .O(N__26109),
            .I(N__26106));
    LocalMux I__4363 (
            .O(N__26106),
            .I(N__26103));
    Odrv12 I__4362 (
            .O(N__26103),
            .I(n22_adj_793));
    CascadeMux I__4361 (
            .O(N__26100),
            .I(\nx.n26_cascade_ ));
    InMux I__4360 (
            .O(N__26097),
            .I(N__26094));
    LocalMux I__4359 (
            .O(N__26094),
            .I(\nx.n20 ));
    CascadeMux I__4358 (
            .O(N__26091),
            .I(\nx.n11912_cascade_ ));
    InMux I__4357 (
            .O(N__26088),
            .I(N__26085));
    LocalMux I__4356 (
            .O(N__26085),
            .I(\nx.n58 ));
    CascadeMux I__4355 (
            .O(N__26082),
            .I(N__26078));
    InMux I__4354 (
            .O(N__26081),
            .I(N__26075));
    InMux I__4353 (
            .O(N__26078),
            .I(N__26070));
    LocalMux I__4352 (
            .O(N__26075),
            .I(N__26065));
    InMux I__4351 (
            .O(N__26074),
            .I(N__26060));
    InMux I__4350 (
            .O(N__26073),
            .I(N__26060));
    LocalMux I__4349 (
            .O(N__26070),
            .I(N__26057));
    InMux I__4348 (
            .O(N__26069),
            .I(N__26054));
    InMux I__4347 (
            .O(N__26068),
            .I(N__26051));
    Span4Mux_h I__4346 (
            .O(N__26065),
            .I(N__26046));
    LocalMux I__4345 (
            .O(N__26060),
            .I(N__26046));
    Sp12to4 I__4344 (
            .O(N__26057),
            .I(N__26041));
    LocalMux I__4343 (
            .O(N__26054),
            .I(N__26041));
    LocalMux I__4342 (
            .O(N__26051),
            .I(\nx.bit_ctr_29 ));
    Odrv4 I__4341 (
            .O(N__26046),
            .I(\nx.bit_ctr_29 ));
    Odrv12 I__4340 (
            .O(N__26041),
            .I(\nx.bit_ctr_29 ));
    CascadeMux I__4339 (
            .O(N__26034),
            .I(N__26030));
    CascadeMux I__4338 (
            .O(N__26033),
            .I(N__26026));
    InMux I__4337 (
            .O(N__26030),
            .I(N__26022));
    InMux I__4336 (
            .O(N__26029),
            .I(N__26017));
    InMux I__4335 (
            .O(N__26026),
            .I(N__26017));
    InMux I__4334 (
            .O(N__26025),
            .I(N__26013));
    LocalMux I__4333 (
            .O(N__26022),
            .I(N__26010));
    LocalMux I__4332 (
            .O(N__26017),
            .I(N__26007));
    InMux I__4331 (
            .O(N__26016),
            .I(N__26004));
    LocalMux I__4330 (
            .O(N__26013),
            .I(N__26001));
    Span4Mux_h I__4329 (
            .O(N__26010),
            .I(N__25996));
    Span4Mux_h I__4328 (
            .O(N__26007),
            .I(N__25996));
    LocalMux I__4327 (
            .O(N__26004),
            .I(\nx.bit_ctr_30 ));
    Odrv12 I__4326 (
            .O(N__26001),
            .I(\nx.bit_ctr_30 ));
    Odrv4 I__4325 (
            .O(N__25996),
            .I(\nx.bit_ctr_30 ));
    CascadeMux I__4324 (
            .O(N__25989),
            .I(N__25986));
    InMux I__4323 (
            .O(N__25986),
            .I(N__25979));
    InMux I__4322 (
            .O(N__25985),
            .I(N__25979));
    CascadeMux I__4321 (
            .O(N__25984),
            .I(N__25975));
    LocalMux I__4320 (
            .O(N__25979),
            .I(N__25971));
    InMux I__4319 (
            .O(N__25978),
            .I(N__25968));
    InMux I__4318 (
            .O(N__25975),
            .I(N__25965));
    InMux I__4317 (
            .O(N__25974),
            .I(N__25962));
    Span4Mux_h I__4316 (
            .O(N__25971),
            .I(N__25959));
    LocalMux I__4315 (
            .O(N__25968),
            .I(N__25954));
    LocalMux I__4314 (
            .O(N__25965),
            .I(N__25954));
    LocalMux I__4313 (
            .O(N__25962),
            .I(\nx.bit_ctr_31 ));
    Odrv4 I__4312 (
            .O(N__25959),
            .I(\nx.bit_ctr_31 ));
    Odrv12 I__4311 (
            .O(N__25954),
            .I(\nx.bit_ctr_31 ));
    InMux I__4310 (
            .O(N__25947),
            .I(N__25944));
    LocalMux I__4309 (
            .O(N__25944),
            .I(\nx.n9803 ));
    InMux I__4308 (
            .O(N__25941),
            .I(N__25935));
    InMux I__4307 (
            .O(N__25940),
            .I(N__25928));
    InMux I__4306 (
            .O(N__25939),
            .I(N__25928));
    InMux I__4305 (
            .O(N__25938),
            .I(N__25928));
    LocalMux I__4304 (
            .O(N__25935),
            .I(N__25922));
    LocalMux I__4303 (
            .O(N__25928),
            .I(N__25919));
    InMux I__4302 (
            .O(N__25927),
            .I(N__25914));
    InMux I__4301 (
            .O(N__25926),
            .I(N__25914));
    InMux I__4300 (
            .O(N__25925),
            .I(N__25911));
    Span4Mux_v I__4299 (
            .O(N__25922),
            .I(N__25904));
    Span4Mux_v I__4298 (
            .O(N__25919),
            .I(N__25904));
    LocalMux I__4297 (
            .O(N__25914),
            .I(N__25904));
    LocalMux I__4296 (
            .O(N__25911),
            .I(\nx.bit_ctr_27 ));
    Odrv4 I__4295 (
            .O(N__25904),
            .I(\nx.bit_ctr_27 ));
    InMux I__4294 (
            .O(N__25899),
            .I(N__25890));
    InMux I__4293 (
            .O(N__25898),
            .I(N__25885));
    InMux I__4292 (
            .O(N__25897),
            .I(N__25885));
    InMux I__4291 (
            .O(N__25896),
            .I(N__25878));
    InMux I__4290 (
            .O(N__25895),
            .I(N__25878));
    InMux I__4289 (
            .O(N__25894),
            .I(N__25878));
    InMux I__4288 (
            .O(N__25893),
            .I(N__25875));
    LocalMux I__4287 (
            .O(N__25890),
            .I(N__25872));
    LocalMux I__4286 (
            .O(N__25885),
            .I(N__25869));
    LocalMux I__4285 (
            .O(N__25878),
            .I(N__25866));
    LocalMux I__4284 (
            .O(N__25875),
            .I(\nx.bit_ctr_28 ));
    Odrv4 I__4283 (
            .O(N__25872),
            .I(\nx.bit_ctr_28 ));
    Odrv12 I__4282 (
            .O(N__25869),
            .I(\nx.bit_ctr_28 ));
    Odrv4 I__4281 (
            .O(N__25866),
            .I(\nx.bit_ctr_28 ));
    CascadeMux I__4280 (
            .O(N__25857),
            .I(N__25852));
    CascadeMux I__4279 (
            .O(N__25856),
            .I(N__25849));
    CascadeMux I__4278 (
            .O(N__25855),
            .I(N__25846));
    InMux I__4277 (
            .O(N__25852),
            .I(N__25843));
    InMux I__4276 (
            .O(N__25849),
            .I(N__25840));
    InMux I__4275 (
            .O(N__25846),
            .I(N__25837));
    LocalMux I__4274 (
            .O(N__25843),
            .I(\nx.n11912 ));
    LocalMux I__4273 (
            .O(N__25840),
            .I(\nx.n11912 ));
    LocalMux I__4272 (
            .O(N__25837),
            .I(\nx.n11912 ));
    InMux I__4271 (
            .O(N__25830),
            .I(N__25824));
    InMux I__4270 (
            .O(N__25829),
            .I(N__25819));
    InMux I__4269 (
            .O(N__25828),
            .I(N__25819));
    InMux I__4268 (
            .O(N__25827),
            .I(N__25816));
    LocalMux I__4267 (
            .O(N__25824),
            .I(\nx.n708 ));
    LocalMux I__4266 (
            .O(N__25819),
            .I(\nx.n708 ));
    LocalMux I__4265 (
            .O(N__25816),
            .I(\nx.n708 ));
    CascadeMux I__4264 (
            .O(N__25809),
            .I(N__25804));
    InMux I__4263 (
            .O(N__25808),
            .I(N__25801));
    InMux I__4262 (
            .O(N__25807),
            .I(N__25796));
    InMux I__4261 (
            .O(N__25804),
            .I(N__25796));
    LocalMux I__4260 (
            .O(N__25801),
            .I(N__25791));
    LocalMux I__4259 (
            .O(N__25796),
            .I(N__25791));
    Odrv4 I__4258 (
            .O(N__25791),
            .I(\nx.n5703 ));
    InMux I__4257 (
            .O(N__25788),
            .I(N__25785));
    LocalMux I__4256 (
            .O(N__25785),
            .I(N__25782));
    Span4Mux_v I__4255 (
            .O(N__25782),
            .I(N__25779));
    Odrv4 I__4254 (
            .O(N__25779),
            .I(n10_adj_846));
    InMux I__4253 (
            .O(N__25776),
            .I(N__25773));
    LocalMux I__4252 (
            .O(N__25773),
            .I(neopxl_color_prev_7));
    CascadeMux I__4251 (
            .O(N__25770),
            .I(N__25766));
    InMux I__4250 (
            .O(N__25769),
            .I(N__25761));
    InMux I__4249 (
            .O(N__25766),
            .I(N__25761));
    LocalMux I__4248 (
            .O(N__25761),
            .I(N__25758));
    Span4Mux_h I__4247 (
            .O(N__25758),
            .I(N__25753));
    InMux I__4246 (
            .O(N__25757),
            .I(N__25750));
    InMux I__4245 (
            .O(N__25756),
            .I(N__25747));
    Span4Mux_v I__4244 (
            .O(N__25753),
            .I(N__25744));
    LocalMux I__4243 (
            .O(N__25750),
            .I(neopxl_color_15));
    LocalMux I__4242 (
            .O(N__25747),
            .I(neopxl_color_15));
    Odrv4 I__4241 (
            .O(N__25744),
            .I(neopxl_color_15));
    InMux I__4240 (
            .O(N__25737),
            .I(N__25734));
    LocalMux I__4239 (
            .O(N__25734),
            .I(neopxl_color_prev_15));
    CascadeMux I__4238 (
            .O(N__25731),
            .I(N__25727));
    CascadeMux I__4237 (
            .O(N__25730),
            .I(N__25724));
    InMux I__4236 (
            .O(N__25727),
            .I(N__25721));
    InMux I__4235 (
            .O(N__25724),
            .I(N__25718));
    LocalMux I__4234 (
            .O(N__25721),
            .I(\nx.n7497 ));
    LocalMux I__4233 (
            .O(N__25718),
            .I(\nx.n7497 ));
    InMux I__4232 (
            .O(N__25713),
            .I(N__25710));
    LocalMux I__4231 (
            .O(N__25710),
            .I(\nx.n976 ));
    InMux I__4230 (
            .O(N__25707),
            .I(\nx.n10738 ));
    CascadeMux I__4229 (
            .O(N__25704),
            .I(N__25701));
    InMux I__4228 (
            .O(N__25701),
            .I(N__25698));
    LocalMux I__4227 (
            .O(N__25698),
            .I(\nx.n7899 ));
    CascadeMux I__4226 (
            .O(N__25695),
            .I(N__25691));
    InMux I__4225 (
            .O(N__25694),
            .I(N__25688));
    InMux I__4224 (
            .O(N__25691),
            .I(N__25685));
    LocalMux I__4223 (
            .O(N__25688),
            .I(\nx.n975 ));
    LocalMux I__4222 (
            .O(N__25685),
            .I(\nx.n975 ));
    InMux I__4221 (
            .O(N__25680),
            .I(\nx.n10739 ));
    InMux I__4220 (
            .O(N__25677),
            .I(N__25671));
    InMux I__4219 (
            .O(N__25676),
            .I(N__25671));
    LocalMux I__4218 (
            .O(N__25671),
            .I(\nx.n974 ));
    InMux I__4217 (
            .O(N__25668),
            .I(\nx.n10740 ));
    CascadeMux I__4216 (
            .O(N__25665),
            .I(N__25661));
    CascadeMux I__4215 (
            .O(N__25664),
            .I(N__25658));
    InMux I__4214 (
            .O(N__25661),
            .I(N__25654));
    InMux I__4213 (
            .O(N__25658),
            .I(N__25651));
    InMux I__4212 (
            .O(N__25657),
            .I(N__25648));
    LocalMux I__4211 (
            .O(N__25654),
            .I(\nx.n906 ));
    LocalMux I__4210 (
            .O(N__25651),
            .I(\nx.n906 ));
    LocalMux I__4209 (
            .O(N__25648),
            .I(\nx.n906 ));
    InMux I__4208 (
            .O(N__25641),
            .I(N__25638));
    LocalMux I__4207 (
            .O(N__25638),
            .I(\nx.n973 ));
    InMux I__4206 (
            .O(N__25635),
            .I(\nx.n10741 ));
    InMux I__4205 (
            .O(N__25632),
            .I(N__25629));
    LocalMux I__4204 (
            .O(N__25629),
            .I(\nx.n13594 ));
    CascadeMux I__4203 (
            .O(N__25626),
            .I(N__25623));
    InMux I__4202 (
            .O(N__25623),
            .I(N__25620));
    LocalMux I__4201 (
            .O(N__25620),
            .I(\nx.n905 ));
    InMux I__4200 (
            .O(N__25617),
            .I(\nx.n10742 ));
    InMux I__4199 (
            .O(N__25614),
            .I(N__25611));
    LocalMux I__4198 (
            .O(N__25611),
            .I(N__25607));
    InMux I__4197 (
            .O(N__25610),
            .I(N__25604));
    Odrv4 I__4196 (
            .O(N__25607),
            .I(\nx.n4 ));
    LocalMux I__4195 (
            .O(N__25604),
            .I(\nx.n4 ));
    CascadeMux I__4194 (
            .O(N__25599),
            .I(N__25596));
    InMux I__4193 (
            .O(N__25596),
            .I(N__25589));
    InMux I__4192 (
            .O(N__25595),
            .I(N__25589));
    InMux I__4191 (
            .O(N__25594),
            .I(N__25586));
    LocalMux I__4190 (
            .O(N__25589),
            .I(\nx.n807 ));
    LocalMux I__4189 (
            .O(N__25586),
            .I(\nx.n807 ));
    CascadeMux I__4188 (
            .O(N__25581),
            .I(N__25576));
    InMux I__4187 (
            .O(N__25580),
            .I(N__25571));
    InMux I__4186 (
            .O(N__25579),
            .I(N__25571));
    InMux I__4185 (
            .O(N__25576),
            .I(N__25568));
    LocalMux I__4184 (
            .O(N__25571),
            .I(\nx.n11866 ));
    LocalMux I__4183 (
            .O(N__25568),
            .I(\nx.n11866 ));
    InMux I__4182 (
            .O(N__25563),
            .I(N__25554));
    InMux I__4181 (
            .O(N__25562),
            .I(N__25554));
    InMux I__4180 (
            .O(N__25561),
            .I(N__25551));
    InMux I__4179 (
            .O(N__25560),
            .I(N__25546));
    InMux I__4178 (
            .O(N__25559),
            .I(N__25546));
    LocalMux I__4177 (
            .O(N__25554),
            .I(\nx.n838 ));
    LocalMux I__4176 (
            .O(N__25551),
            .I(\nx.n838 ));
    LocalMux I__4175 (
            .O(N__25546),
            .I(\nx.n838 ));
    CascadeMux I__4174 (
            .O(N__25539),
            .I(N__25536));
    InMux I__4173 (
            .O(N__25536),
            .I(N__25532));
    InMux I__4172 (
            .O(N__25535),
            .I(N__25529));
    LocalMux I__4171 (
            .O(N__25532),
            .I(\nx.n11868 ));
    LocalMux I__4170 (
            .O(N__25529),
            .I(\nx.n11868 ));
    InMux I__4169 (
            .O(N__25524),
            .I(N__25519));
    InMux I__4168 (
            .O(N__25523),
            .I(N__25516));
    InMux I__4167 (
            .O(N__25522),
            .I(N__25511));
    LocalMux I__4166 (
            .O(N__25519),
            .I(N__25506));
    LocalMux I__4165 (
            .O(N__25516),
            .I(N__25506));
    InMux I__4164 (
            .O(N__25515),
            .I(N__25503));
    InMux I__4163 (
            .O(N__25514),
            .I(N__25500));
    LocalMux I__4162 (
            .O(N__25511),
            .I(N__25497));
    Span4Mux_v I__4161 (
            .O(N__25506),
            .I(N__25494));
    LocalMux I__4160 (
            .O(N__25503),
            .I(N__25491));
    LocalMux I__4159 (
            .O(N__25500),
            .I(\nx.bit_ctr_17 ));
    Odrv4 I__4158 (
            .O(N__25497),
            .I(\nx.bit_ctr_17 ));
    Odrv4 I__4157 (
            .O(N__25494),
            .I(\nx.bit_ctr_17 ));
    Odrv12 I__4156 (
            .O(N__25491),
            .I(\nx.bit_ctr_17 ));
    InMux I__4155 (
            .O(N__25482),
            .I(N__25478));
    CascadeMux I__4154 (
            .O(N__25481),
            .I(N__25473));
    LocalMux I__4153 (
            .O(N__25478),
            .I(N__25470));
    InMux I__4152 (
            .O(N__25477),
            .I(N__25467));
    InMux I__4151 (
            .O(N__25476),
            .I(N__25464));
    InMux I__4150 (
            .O(N__25473),
            .I(N__25460));
    Span4Mux_v I__4149 (
            .O(N__25470),
            .I(N__25455));
    LocalMux I__4148 (
            .O(N__25467),
            .I(N__25455));
    LocalMux I__4147 (
            .O(N__25464),
            .I(N__25452));
    InMux I__4146 (
            .O(N__25463),
            .I(N__25449));
    LocalMux I__4145 (
            .O(N__25460),
            .I(N__25446));
    Span4Mux_h I__4144 (
            .O(N__25455),
            .I(N__25441));
    Span4Mux_h I__4143 (
            .O(N__25452),
            .I(N__25441));
    LocalMux I__4142 (
            .O(N__25449),
            .I(\nx.bit_ctr_22 ));
    Odrv4 I__4141 (
            .O(N__25446),
            .I(\nx.bit_ctr_22 ));
    Odrv4 I__4140 (
            .O(N__25441),
            .I(\nx.bit_ctr_22 ));
    InMux I__4139 (
            .O(N__25434),
            .I(N__25431));
    LocalMux I__4138 (
            .O(N__25431),
            .I(N__25428));
    Span4Mux_h I__4137 (
            .O(N__25428),
            .I(N__25425));
    Odrv4 I__4136 (
            .O(N__25425),
            .I(\nx.n44_adj_782 ));
    InMux I__4135 (
            .O(N__25422),
            .I(N__25419));
    LocalMux I__4134 (
            .O(N__25419),
            .I(\nx.n11941 ));
    CascadeMux I__4133 (
            .O(N__25416),
            .I(N__25412));
    CascadeMux I__4132 (
            .O(N__25415),
            .I(N__25408));
    InMux I__4131 (
            .O(N__25412),
            .I(N__25403));
    InMux I__4130 (
            .O(N__25411),
            .I(N__25403));
    InMux I__4129 (
            .O(N__25408),
            .I(N__25400));
    LocalMux I__4128 (
            .O(N__25403),
            .I(\nx.n1008 ));
    LocalMux I__4127 (
            .O(N__25400),
            .I(\nx.n1008 ));
    CascadeMux I__4126 (
            .O(N__25395),
            .I(N__25391));
    InMux I__4125 (
            .O(N__25394),
            .I(N__25388));
    InMux I__4124 (
            .O(N__25391),
            .I(N__25385));
    LocalMux I__4123 (
            .O(N__25388),
            .I(\nx.n1006 ));
    LocalMux I__4122 (
            .O(N__25385),
            .I(\nx.n1006 ));
    CascadeMux I__4121 (
            .O(N__25380),
            .I(\nx.n12837_cascade_ ));
    CascadeMux I__4120 (
            .O(N__25377),
            .I(\nx.n905_cascade_ ));
    InMux I__4119 (
            .O(N__25374),
            .I(N__25371));
    LocalMux I__4118 (
            .O(N__25371),
            .I(\nx.n12839 ));
    CascadeMux I__4117 (
            .O(N__25368),
            .I(N__25362));
    CascadeMux I__4116 (
            .O(N__25367),
            .I(N__25359));
    InMux I__4115 (
            .O(N__25366),
            .I(N__25352));
    InMux I__4114 (
            .O(N__25365),
            .I(N__25352));
    InMux I__4113 (
            .O(N__25362),
            .I(N__25345));
    InMux I__4112 (
            .O(N__25359),
            .I(N__25345));
    InMux I__4111 (
            .O(N__25358),
            .I(N__25345));
    InMux I__4110 (
            .O(N__25357),
            .I(N__25342));
    LocalMux I__4109 (
            .O(N__25352),
            .I(\nx.n11174 ));
    LocalMux I__4108 (
            .O(N__25345),
            .I(\nx.n11174 ));
    LocalMux I__4107 (
            .O(N__25342),
            .I(\nx.n11174 ));
    CascadeMux I__4106 (
            .O(N__25335),
            .I(\nx.n11174_cascade_ ));
    CascadeMux I__4105 (
            .O(N__25332),
            .I(N__25329));
    InMux I__4104 (
            .O(N__25329),
            .I(N__25323));
    InMux I__4103 (
            .O(N__25328),
            .I(N__25320));
    InMux I__4102 (
            .O(N__25327),
            .I(N__25317));
    InMux I__4101 (
            .O(N__25326),
            .I(N__25314));
    LocalMux I__4100 (
            .O(N__25323),
            .I(N__25310));
    LocalMux I__4099 (
            .O(N__25320),
            .I(N__25307));
    LocalMux I__4098 (
            .O(N__25317),
            .I(N__25302));
    LocalMux I__4097 (
            .O(N__25314),
            .I(N__25302));
    InMux I__4096 (
            .O(N__25313),
            .I(N__25299));
    Span4Mux_h I__4095 (
            .O(N__25310),
            .I(N__25296));
    Span4Mux_v I__4094 (
            .O(N__25307),
            .I(N__25291));
    Span4Mux_h I__4093 (
            .O(N__25302),
            .I(N__25291));
    LocalMux I__4092 (
            .O(N__25299),
            .I(\nx.bit_ctr_26 ));
    Odrv4 I__4091 (
            .O(N__25296),
            .I(\nx.bit_ctr_26 ));
    Odrv4 I__4090 (
            .O(N__25291),
            .I(\nx.bit_ctr_26 ));
    CascadeMux I__4089 (
            .O(N__25284),
            .I(N__25281));
    InMux I__4088 (
            .O(N__25281),
            .I(N__25278));
    LocalMux I__4087 (
            .O(N__25278),
            .I(N__25275));
    Odrv4 I__4086 (
            .O(N__25275),
            .I(\nx.n977 ));
    InMux I__4085 (
            .O(N__25272),
            .I(bfn_7_22_0_));
    InMux I__4084 (
            .O(N__25269),
            .I(N__25265));
    CascadeMux I__4083 (
            .O(N__25268),
            .I(N__25262));
    LocalMux I__4082 (
            .O(N__25265),
            .I(N__25259));
    InMux I__4081 (
            .O(N__25262),
            .I(N__25255));
    Span4Mux_h I__4080 (
            .O(N__25259),
            .I(N__25252));
    InMux I__4079 (
            .O(N__25258),
            .I(N__25249));
    LocalMux I__4078 (
            .O(N__25255),
            .I(N__25246));
    Odrv4 I__4077 (
            .O(N__25252),
            .I(timer_28));
    LocalMux I__4076 (
            .O(N__25249),
            .I(timer_28));
    Odrv4 I__4075 (
            .O(N__25246),
            .I(timer_28));
    InMux I__4074 (
            .O(N__25239),
            .I(N__25221));
    InMux I__4073 (
            .O(N__25238),
            .I(N__25213));
    InMux I__4072 (
            .O(N__25237),
            .I(N__25208));
    InMux I__4071 (
            .O(N__25236),
            .I(N__25208));
    InMux I__4070 (
            .O(N__25235),
            .I(N__25201));
    InMux I__4069 (
            .O(N__25234),
            .I(N__25201));
    InMux I__4068 (
            .O(N__25233),
            .I(N__25201));
    InMux I__4067 (
            .O(N__25232),
            .I(N__25194));
    InMux I__4066 (
            .O(N__25231),
            .I(N__25194));
    InMux I__4065 (
            .O(N__25230),
            .I(N__25194));
    InMux I__4064 (
            .O(N__25229),
            .I(N__25185));
    InMux I__4063 (
            .O(N__25228),
            .I(N__25185));
    InMux I__4062 (
            .O(N__25227),
            .I(N__25185));
    InMux I__4061 (
            .O(N__25226),
            .I(N__25185));
    InMux I__4060 (
            .O(N__25225),
            .I(N__25180));
    InMux I__4059 (
            .O(N__25224),
            .I(N__25180));
    LocalMux I__4058 (
            .O(N__25221),
            .I(N__25173));
    InMux I__4057 (
            .O(N__25220),
            .I(N__25170));
    InMux I__4056 (
            .O(N__25219),
            .I(N__25167));
    InMux I__4055 (
            .O(N__25218),
            .I(N__25158));
    InMux I__4054 (
            .O(N__25217),
            .I(N__25158));
    InMux I__4053 (
            .O(N__25216),
            .I(N__25158));
    LocalMux I__4052 (
            .O(N__25213),
            .I(N__25152));
    LocalMux I__4051 (
            .O(N__25208),
            .I(N__25143));
    LocalMux I__4050 (
            .O(N__25201),
            .I(N__25143));
    LocalMux I__4049 (
            .O(N__25194),
            .I(N__25143));
    LocalMux I__4048 (
            .O(N__25185),
            .I(N__25143));
    LocalMux I__4047 (
            .O(N__25180),
            .I(N__25140));
    InMux I__4046 (
            .O(N__25179),
            .I(N__25131));
    InMux I__4045 (
            .O(N__25178),
            .I(N__25131));
    InMux I__4044 (
            .O(N__25177),
            .I(N__25131));
    InMux I__4043 (
            .O(N__25176),
            .I(N__25131));
    Span4Mux_s3_h I__4042 (
            .O(N__25173),
            .I(N__25126));
    LocalMux I__4041 (
            .O(N__25170),
            .I(N__25126));
    LocalMux I__4040 (
            .O(N__25167),
            .I(N__25123));
    InMux I__4039 (
            .O(N__25166),
            .I(N__25118));
    InMux I__4038 (
            .O(N__25165),
            .I(N__25118));
    LocalMux I__4037 (
            .O(N__25158),
            .I(N__25113));
    InMux I__4036 (
            .O(N__25157),
            .I(N__25110));
    InMux I__4035 (
            .O(N__25156),
            .I(N__25107));
    InMux I__4034 (
            .O(N__25155),
            .I(N__25104));
    Span4Mux_v I__4033 (
            .O(N__25152),
            .I(N__25095));
    Span4Mux_v I__4032 (
            .O(N__25143),
            .I(N__25095));
    Span4Mux_s1_h I__4031 (
            .O(N__25140),
            .I(N__25095));
    LocalMux I__4030 (
            .O(N__25131),
            .I(N__25095));
    Span4Mux_v I__4029 (
            .O(N__25126),
            .I(N__25088));
    Span4Mux_h I__4028 (
            .O(N__25123),
            .I(N__25088));
    LocalMux I__4027 (
            .O(N__25118),
            .I(N__25088));
    InMux I__4026 (
            .O(N__25117),
            .I(N__25083));
    InMux I__4025 (
            .O(N__25116),
            .I(N__25083));
    Odrv12 I__4024 (
            .O(N__25113),
            .I(n11353));
    LocalMux I__4023 (
            .O(N__25110),
            .I(n11353));
    LocalMux I__4022 (
            .O(N__25107),
            .I(n11353));
    LocalMux I__4021 (
            .O(N__25104),
            .I(n11353));
    Odrv4 I__4020 (
            .O(N__25095),
            .I(n11353));
    Odrv4 I__4019 (
            .O(N__25088),
            .I(n11353));
    LocalMux I__4018 (
            .O(N__25083),
            .I(n11353));
    InMux I__4017 (
            .O(N__25068),
            .I(N__25064));
    InMux I__4016 (
            .O(N__25067),
            .I(N__25061));
    LocalMux I__4015 (
            .O(N__25064),
            .I(N__25058));
    LocalMux I__4014 (
            .O(N__25061),
            .I(neo_pixel_transmitter_t0_28));
    Odrv4 I__4013 (
            .O(N__25058),
            .I(neo_pixel_transmitter_t0_28));
    InMux I__4012 (
            .O(N__25053),
            .I(N__25050));
    LocalMux I__4011 (
            .O(N__25050),
            .I(n9_adj_847));
    SRMux I__4010 (
            .O(N__25047),
            .I(N__25044));
    LocalMux I__4009 (
            .O(N__25044),
            .I(N__25041));
    Span4Mux_v I__4008 (
            .O(N__25041),
            .I(N__25038));
    Span4Mux_h I__4007 (
            .O(N__25038),
            .I(N__25035));
    Odrv4 I__4006 (
            .O(N__25035),
            .I(current_pin_7__N_153));
    InMux I__4005 (
            .O(N__25032),
            .I(N__25029));
    LocalMux I__4004 (
            .O(N__25029),
            .I(neopxl_color_prev_14));
    CascadeMux I__4003 (
            .O(N__25026),
            .I(N__25020));
    InMux I__4002 (
            .O(N__25025),
            .I(N__25017));
    InMux I__4001 (
            .O(N__25024),
            .I(N__25010));
    InMux I__4000 (
            .O(N__25023),
            .I(N__25010));
    InMux I__3999 (
            .O(N__25020),
            .I(N__25010));
    LocalMux I__3998 (
            .O(N__25017),
            .I(N__25007));
    LocalMux I__3997 (
            .O(N__25010),
            .I(neopxl_color_13));
    Odrv4 I__3996 (
            .O(N__25007),
            .I(neopxl_color_13));
    InMux I__3995 (
            .O(N__25002),
            .I(N__24999));
    LocalMux I__3994 (
            .O(N__24999),
            .I(neopxl_color_prev_13));
    InMux I__3993 (
            .O(N__24996),
            .I(N__24993));
    LocalMux I__3992 (
            .O(N__24993),
            .I(n11_adj_845));
    InMux I__3991 (
            .O(N__24990),
            .I(N__24987));
    LocalMux I__3990 (
            .O(N__24987),
            .I(neopxl_color_prev_4));
    InMux I__3989 (
            .O(N__24984),
            .I(N__24980));
    CascadeMux I__3988 (
            .O(N__24983),
            .I(N__24975));
    LocalMux I__3987 (
            .O(N__24980),
            .I(N__24972));
    InMux I__3986 (
            .O(N__24979),
            .I(N__24965));
    InMux I__3985 (
            .O(N__24978),
            .I(N__24965));
    InMux I__3984 (
            .O(N__24975),
            .I(N__24965));
    Span4Mux_h I__3983 (
            .O(N__24972),
            .I(N__24962));
    LocalMux I__3982 (
            .O(N__24965),
            .I(neopxl_color_14));
    Odrv4 I__3981 (
            .O(N__24962),
            .I(neopxl_color_14));
    CascadeMux I__3980 (
            .O(N__24957),
            .I(N__24952));
    CascadeMux I__3979 (
            .O(N__24956),
            .I(N__24949));
    InMux I__3978 (
            .O(N__24955),
            .I(N__24946));
    InMux I__3977 (
            .O(N__24952),
            .I(N__24937));
    InMux I__3976 (
            .O(N__24949),
            .I(N__24934));
    LocalMux I__3975 (
            .O(N__24946),
            .I(N__24930));
    InMux I__3974 (
            .O(N__24945),
            .I(N__24927));
    InMux I__3973 (
            .O(N__24944),
            .I(N__24920));
    InMux I__3972 (
            .O(N__24943),
            .I(N__24920));
    InMux I__3971 (
            .O(N__24942),
            .I(N__24920));
    InMux I__3970 (
            .O(N__24941),
            .I(N__24915));
    InMux I__3969 (
            .O(N__24940),
            .I(N__24915));
    LocalMux I__3968 (
            .O(N__24937),
            .I(N__24912));
    LocalMux I__3967 (
            .O(N__24934),
            .I(N__24909));
    InMux I__3966 (
            .O(N__24933),
            .I(N__24904));
    Span4Mux_h I__3965 (
            .O(N__24930),
            .I(N__24895));
    LocalMux I__3964 (
            .O(N__24927),
            .I(N__24895));
    LocalMux I__3963 (
            .O(N__24920),
            .I(N__24895));
    LocalMux I__3962 (
            .O(N__24915),
            .I(N__24895));
    Span4Mux_h I__3961 (
            .O(N__24912),
            .I(N__24892));
    Span4Mux_h I__3960 (
            .O(N__24909),
            .I(N__24889));
    InMux I__3959 (
            .O(N__24908),
            .I(N__24884));
    InMux I__3958 (
            .O(N__24907),
            .I(N__24884));
    LocalMux I__3957 (
            .O(N__24904),
            .I(\nx.neo_pixel_transmitter_done ));
    Odrv4 I__3956 (
            .O(N__24895),
            .I(\nx.neo_pixel_transmitter_done ));
    Odrv4 I__3955 (
            .O(N__24892),
            .I(\nx.neo_pixel_transmitter_done ));
    Odrv4 I__3954 (
            .O(N__24889),
            .I(\nx.neo_pixel_transmitter_done ));
    LocalMux I__3953 (
            .O(N__24884),
            .I(\nx.neo_pixel_transmitter_done ));
    IoInMux I__3952 (
            .O(N__24873),
            .I(N__24870));
    LocalMux I__3951 (
            .O(N__24870),
            .I(N__24867));
    Odrv12 I__3950 (
            .O(N__24867),
            .I(NEOPXL_c));
    CEMux I__3949 (
            .O(N__24864),
            .I(N__24861));
    LocalMux I__3948 (
            .O(N__24861),
            .I(N__24858));
    Odrv12 I__3947 (
            .O(N__24858),
            .I(\nx.n11988 ));
    SRMux I__3946 (
            .O(N__24855),
            .I(N__24852));
    LocalMux I__3945 (
            .O(N__24852),
            .I(N__24849));
    Odrv4 I__3944 (
            .O(N__24849),
            .I(\nx.n12451 ));
    InMux I__3943 (
            .O(N__24846),
            .I(N__24843));
    LocalMux I__3942 (
            .O(N__24843),
            .I(N__24839));
    InMux I__3941 (
            .O(N__24842),
            .I(N__24836));
    Span4Mux_v I__3940 (
            .O(N__24839),
            .I(N__24833));
    LocalMux I__3939 (
            .O(N__24836),
            .I(\nx.bit_ctr_1 ));
    Odrv4 I__3938 (
            .O(N__24833),
            .I(\nx.bit_ctr_1 ));
    InMux I__3937 (
            .O(N__24828),
            .I(N__24825));
    LocalMux I__3936 (
            .O(N__24825),
            .I(\nx.n13364 ));
    CascadeMux I__3935 (
            .O(N__24822),
            .I(\nx.n11156_cascade_ ));
    InMux I__3934 (
            .O(N__24819),
            .I(N__24816));
    LocalMux I__3933 (
            .O(N__24816),
            .I(\nx.n13363 ));
    CascadeMux I__3932 (
            .O(N__24813),
            .I(\nx.n13619_cascade_ ));
    InMux I__3931 (
            .O(N__24810),
            .I(N__24807));
    LocalMux I__3930 (
            .O(N__24807),
            .I(\nx.n11156 ));
    InMux I__3929 (
            .O(N__24804),
            .I(N__24801));
    LocalMux I__3928 (
            .O(N__24801),
            .I(N__24798));
    Span4Mux_h I__3927 (
            .O(N__24798),
            .I(N__24795));
    Odrv4 I__3926 (
            .O(N__24795),
            .I(n11966));
    IoInMux I__3925 (
            .O(N__24792),
            .I(N__24789));
    LocalMux I__3924 (
            .O(N__24789),
            .I(N__24786));
    Span4Mux_s2_h I__3923 (
            .O(N__24786),
            .I(N__24783));
    Span4Mux_h I__3922 (
            .O(N__24783),
            .I(N__24779));
    InMux I__3921 (
            .O(N__24782),
            .I(N__24776));
    Odrv4 I__3920 (
            .O(N__24779),
            .I(pin_oe_2));
    LocalMux I__3919 (
            .O(N__24776),
            .I(pin_oe_2));
    InMux I__3918 (
            .O(N__24771),
            .I(N__24768));
    LocalMux I__3917 (
            .O(N__24768),
            .I(\nx.n13372 ));
    CascadeMux I__3916 (
            .O(N__24765),
            .I(N__24760));
    InMux I__3915 (
            .O(N__24764),
            .I(N__24757));
    InMux I__3914 (
            .O(N__24763),
            .I(N__24754));
    InMux I__3913 (
            .O(N__24760),
            .I(N__24750));
    LocalMux I__3912 (
            .O(N__24757),
            .I(N__24747));
    LocalMux I__3911 (
            .O(N__24754),
            .I(N__24744));
    InMux I__3910 (
            .O(N__24753),
            .I(N__24740));
    LocalMux I__3909 (
            .O(N__24750),
            .I(N__24737));
    Span12Mux_s5_h I__3908 (
            .O(N__24747),
            .I(N__24734));
    Span4Mux_v I__3907 (
            .O(N__24744),
            .I(N__24731));
    InMux I__3906 (
            .O(N__24743),
            .I(N__24728));
    LocalMux I__3905 (
            .O(N__24740),
            .I(\nx.bit_ctr_18 ));
    Odrv12 I__3904 (
            .O(N__24737),
            .I(\nx.bit_ctr_18 ));
    Odrv12 I__3903 (
            .O(N__24734),
            .I(\nx.bit_ctr_18 ));
    Odrv4 I__3902 (
            .O(N__24731),
            .I(\nx.bit_ctr_18 ));
    LocalMux I__3901 (
            .O(N__24728),
            .I(\nx.bit_ctr_18 ));
    CascadeMux I__3900 (
            .O(N__24717),
            .I(N__24714));
    InMux I__3899 (
            .O(N__24714),
            .I(N__24711));
    LocalMux I__3898 (
            .O(N__24711),
            .I(N__24708));
    Span4Mux_h I__3897 (
            .O(N__24708),
            .I(N__24705));
    Odrv4 I__3896 (
            .O(N__24705),
            .I(\nx.n48_adj_778 ));
    InMux I__3895 (
            .O(N__24702),
            .I(N__24699));
    LocalMux I__3894 (
            .O(N__24699),
            .I(\nx.n18_adj_716 ));
    InMux I__3893 (
            .O(N__24696),
            .I(N__24691));
    InMux I__3892 (
            .O(N__24695),
            .I(N__24688));
    InMux I__3891 (
            .O(N__24694),
            .I(N__24685));
    LocalMux I__3890 (
            .O(N__24691),
            .I(\nx.n1799 ));
    LocalMux I__3889 (
            .O(N__24688),
            .I(\nx.n1799 ));
    LocalMux I__3888 (
            .O(N__24685),
            .I(\nx.n1799 ));
    CascadeMux I__3887 (
            .O(N__24678),
            .I(N__24675));
    InMux I__3886 (
            .O(N__24675),
            .I(N__24670));
    InMux I__3885 (
            .O(N__24674),
            .I(N__24667));
    InMux I__3884 (
            .O(N__24673),
            .I(N__24664));
    LocalMux I__3883 (
            .O(N__24670),
            .I(N__24661));
    LocalMux I__3882 (
            .O(N__24667),
            .I(\nx.n1805 ));
    LocalMux I__3881 (
            .O(N__24664),
            .I(\nx.n1805 ));
    Odrv4 I__3880 (
            .O(N__24661),
            .I(\nx.n1805 ));
    InMux I__3879 (
            .O(N__24654),
            .I(N__24651));
    LocalMux I__3878 (
            .O(N__24651),
            .I(\nx.n24_adj_717 ));
    InMux I__3877 (
            .O(N__24648),
            .I(N__24644));
    InMux I__3876 (
            .O(N__24647),
            .I(N__24641));
    LocalMux I__3875 (
            .O(N__24644),
            .I(N__24635));
    LocalMux I__3874 (
            .O(N__24641),
            .I(N__24635));
    InMux I__3873 (
            .O(N__24640),
            .I(N__24632));
    Odrv4 I__3872 (
            .O(N__24635),
            .I(\nx.n1798 ));
    LocalMux I__3871 (
            .O(N__24632),
            .I(\nx.n1798 ));
    InMux I__3870 (
            .O(N__24627),
            .I(N__24622));
    InMux I__3869 (
            .O(N__24626),
            .I(N__24619));
    InMux I__3868 (
            .O(N__24625),
            .I(N__24616));
    LocalMux I__3867 (
            .O(N__24622),
            .I(N__24613));
    LocalMux I__3866 (
            .O(N__24619),
            .I(\nx.n1808 ));
    LocalMux I__3865 (
            .O(N__24616),
            .I(\nx.n1808 ));
    Odrv4 I__3864 (
            .O(N__24613),
            .I(\nx.n1808 ));
    CascadeMux I__3863 (
            .O(N__24606),
            .I(\nx.n26_adj_719_cascade_ ));
    InMux I__3862 (
            .O(N__24603),
            .I(N__24598));
    InMux I__3861 (
            .O(N__24602),
            .I(N__24595));
    InMux I__3860 (
            .O(N__24601),
            .I(N__24592));
    LocalMux I__3859 (
            .O(N__24598),
            .I(N__24589));
    LocalMux I__3858 (
            .O(N__24595),
            .I(\nx.n1809 ));
    LocalMux I__3857 (
            .O(N__24592),
            .I(\nx.n1809 ));
    Odrv4 I__3856 (
            .O(N__24589),
            .I(\nx.n1809 ));
    InMux I__3855 (
            .O(N__24582),
            .I(N__24577));
    InMux I__3854 (
            .O(N__24581),
            .I(N__24574));
    InMux I__3853 (
            .O(N__24580),
            .I(N__24571));
    LocalMux I__3852 (
            .O(N__24577),
            .I(N__24568));
    LocalMux I__3851 (
            .O(N__24574),
            .I(\nx.n1803 ));
    LocalMux I__3850 (
            .O(N__24571),
            .I(\nx.n1803 ));
    Odrv4 I__3849 (
            .O(N__24568),
            .I(\nx.n1803 ));
    InMux I__3848 (
            .O(N__24561),
            .I(N__24556));
    InMux I__3847 (
            .O(N__24560),
            .I(N__24553));
    InMux I__3846 (
            .O(N__24559),
            .I(N__24550));
    LocalMux I__3845 (
            .O(N__24556),
            .I(\nx.n1800 ));
    LocalMux I__3844 (
            .O(N__24553),
            .I(\nx.n1800 ));
    LocalMux I__3843 (
            .O(N__24550),
            .I(\nx.n1800 ));
    CascadeMux I__3842 (
            .O(N__24543),
            .I(\nx.n9717_cascade_ ));
    InMux I__3841 (
            .O(N__24540),
            .I(N__24535));
    InMux I__3840 (
            .O(N__24539),
            .I(N__24532));
    InMux I__3839 (
            .O(N__24538),
            .I(N__24529));
    LocalMux I__3838 (
            .O(N__24535),
            .I(\nx.n1796 ));
    LocalMux I__3837 (
            .O(N__24532),
            .I(\nx.n1796 ));
    LocalMux I__3836 (
            .O(N__24529),
            .I(\nx.n1796 ));
    InMux I__3835 (
            .O(N__24522),
            .I(N__24519));
    LocalMux I__3834 (
            .O(N__24519),
            .I(\nx.n22_adj_718 ));
    CascadeMux I__3833 (
            .O(N__24516),
            .I(N__24501));
    CascadeMux I__3832 (
            .O(N__24515),
            .I(N__24498));
    CascadeMux I__3831 (
            .O(N__24514),
            .I(N__24495));
    CascadeMux I__3830 (
            .O(N__24513),
            .I(N__24492));
    CascadeMux I__3829 (
            .O(N__24512),
            .I(N__24489));
    CascadeMux I__3828 (
            .O(N__24511),
            .I(N__24486));
    CascadeMux I__3827 (
            .O(N__24510),
            .I(N__24483));
    CascadeMux I__3826 (
            .O(N__24509),
            .I(N__24480));
    CascadeMux I__3825 (
            .O(N__24508),
            .I(N__24477));
    CascadeMux I__3824 (
            .O(N__24507),
            .I(N__24474));
    CascadeMux I__3823 (
            .O(N__24506),
            .I(N__24471));
    CascadeMux I__3822 (
            .O(N__24505),
            .I(N__24468));
    CascadeMux I__3821 (
            .O(N__24504),
            .I(N__24465));
    InMux I__3820 (
            .O(N__24501),
            .I(N__24458));
    InMux I__3819 (
            .O(N__24498),
            .I(N__24458));
    InMux I__3818 (
            .O(N__24495),
            .I(N__24458));
    InMux I__3817 (
            .O(N__24492),
            .I(N__24451));
    InMux I__3816 (
            .O(N__24489),
            .I(N__24451));
    InMux I__3815 (
            .O(N__24486),
            .I(N__24451));
    InMux I__3814 (
            .O(N__24483),
            .I(N__24443));
    InMux I__3813 (
            .O(N__24480),
            .I(N__24443));
    InMux I__3812 (
            .O(N__24477),
            .I(N__24443));
    InMux I__3811 (
            .O(N__24474),
            .I(N__24434));
    InMux I__3810 (
            .O(N__24471),
            .I(N__24434));
    InMux I__3809 (
            .O(N__24468),
            .I(N__24434));
    InMux I__3808 (
            .O(N__24465),
            .I(N__24434));
    LocalMux I__3807 (
            .O(N__24458),
            .I(N__24429));
    LocalMux I__3806 (
            .O(N__24451),
            .I(N__24429));
    InMux I__3805 (
            .O(N__24450),
            .I(N__24426));
    LocalMux I__3804 (
            .O(N__24443),
            .I(\nx.n1829 ));
    LocalMux I__3803 (
            .O(N__24434),
            .I(\nx.n1829 ));
    Odrv4 I__3802 (
            .O(N__24429),
            .I(\nx.n1829 ));
    LocalMux I__3801 (
            .O(N__24426),
            .I(\nx.n1829 ));
    CascadeMux I__3800 (
            .O(N__24417),
            .I(N__24413));
    CascadeMux I__3799 (
            .O(N__24416),
            .I(N__24410));
    InMux I__3798 (
            .O(N__24413),
            .I(N__24407));
    InMux I__3797 (
            .O(N__24410),
            .I(N__24404));
    LocalMux I__3796 (
            .O(N__24407),
            .I(N__24399));
    LocalMux I__3795 (
            .O(N__24404),
            .I(N__24399));
    Odrv4 I__3794 (
            .O(N__24399),
            .I(\nx.n13605 ));
    IoInMux I__3793 (
            .O(N__24396),
            .I(N__24393));
    LocalMux I__3792 (
            .O(N__24393),
            .I(N__24390));
    Span12Mux_s1_h I__3791 (
            .O(N__24390),
            .I(N__24387));
    Span12Mux_h I__3790 (
            .O(N__24387),
            .I(N__24384));
    Span12Mux_v I__3789 (
            .O(N__24384),
            .I(N__24380));
    InMux I__3788 (
            .O(N__24383),
            .I(N__24377));
    Odrv12 I__3787 (
            .O(N__24380),
            .I(pin_oe_7));
    LocalMux I__3786 (
            .O(N__24377),
            .I(pin_oe_7));
    InMux I__3785 (
            .O(N__24372),
            .I(N__24367));
    InMux I__3784 (
            .O(N__24371),
            .I(N__24364));
    InMux I__3783 (
            .O(N__24370),
            .I(N__24361));
    LocalMux I__3782 (
            .O(N__24367),
            .I(N__24358));
    LocalMux I__3781 (
            .O(N__24364),
            .I(\nx.n1804 ));
    LocalMux I__3780 (
            .O(N__24361),
            .I(\nx.n1804 ));
    Odrv4 I__3779 (
            .O(N__24358),
            .I(\nx.n1804 ));
    InMux I__3778 (
            .O(N__24351),
            .I(\nx.n10824 ));
    InMux I__3777 (
            .O(N__24348),
            .I(\nx.n10825 ));
    InMux I__3776 (
            .O(N__24345),
            .I(N__24340));
    InMux I__3775 (
            .O(N__24344),
            .I(N__24337));
    InMux I__3774 (
            .O(N__24343),
            .I(N__24334));
    LocalMux I__3773 (
            .O(N__24340),
            .I(N__24331));
    LocalMux I__3772 (
            .O(N__24337),
            .I(\nx.n1802 ));
    LocalMux I__3771 (
            .O(N__24334),
            .I(\nx.n1802 ));
    Odrv4 I__3770 (
            .O(N__24331),
            .I(\nx.n1802 ));
    InMux I__3769 (
            .O(N__24324),
            .I(bfn_6_28_0_));
    CascadeMux I__3768 (
            .O(N__24321),
            .I(N__24316));
    InMux I__3767 (
            .O(N__24320),
            .I(N__24313));
    InMux I__3766 (
            .O(N__24319),
            .I(N__24310));
    InMux I__3765 (
            .O(N__24316),
            .I(N__24307));
    LocalMux I__3764 (
            .O(N__24313),
            .I(\nx.n1801 ));
    LocalMux I__3763 (
            .O(N__24310),
            .I(\nx.n1801 ));
    LocalMux I__3762 (
            .O(N__24307),
            .I(\nx.n1801 ));
    InMux I__3761 (
            .O(N__24300),
            .I(\nx.n10827 ));
    InMux I__3760 (
            .O(N__24297),
            .I(\nx.n10828 ));
    InMux I__3759 (
            .O(N__24294),
            .I(\nx.n10829 ));
    InMux I__3758 (
            .O(N__24291),
            .I(\nx.n10830 ));
    InMux I__3757 (
            .O(N__24288),
            .I(N__24283));
    InMux I__3756 (
            .O(N__24287),
            .I(N__24280));
    InMux I__3755 (
            .O(N__24286),
            .I(N__24277));
    LocalMux I__3754 (
            .O(N__24283),
            .I(\nx.n1797 ));
    LocalMux I__3753 (
            .O(N__24280),
            .I(\nx.n1797 ));
    LocalMux I__3752 (
            .O(N__24277),
            .I(\nx.n1797 ));
    InMux I__3751 (
            .O(N__24270),
            .I(\nx.n10831 ));
    InMux I__3750 (
            .O(N__24267),
            .I(\nx.n10832 ));
    InMux I__3749 (
            .O(N__24264),
            .I(\nx.n10641 ));
    InMux I__3748 (
            .O(N__24261),
            .I(\nx.n10642 ));
    InMux I__3747 (
            .O(N__24258),
            .I(\nx.n10643 ));
    CEMux I__3746 (
            .O(N__24255),
            .I(N__24251));
    CEMux I__3745 (
            .O(N__24254),
            .I(N__24247));
    LocalMux I__3744 (
            .O(N__24251),
            .I(N__24244));
    CEMux I__3743 (
            .O(N__24250),
            .I(N__24241));
    LocalMux I__3742 (
            .O(N__24247),
            .I(N__24237));
    Span4Mux_h I__3741 (
            .O(N__24244),
            .I(N__24232));
    LocalMux I__3740 (
            .O(N__24241),
            .I(N__24232));
    CEMux I__3739 (
            .O(N__24240),
            .I(N__24229));
    Span4Mux_v I__3738 (
            .O(N__24237),
            .I(N__24226));
    Span4Mux_v I__3737 (
            .O(N__24232),
            .I(N__24223));
    LocalMux I__3736 (
            .O(N__24229),
            .I(N__24220));
    Odrv4 I__3735 (
            .O(N__24226),
            .I(\nx.n7657 ));
    Odrv4 I__3734 (
            .O(N__24223),
            .I(\nx.n7657 ));
    Odrv12 I__3733 (
            .O(N__24220),
            .I(\nx.n7657 ));
    SRMux I__3732 (
            .O(N__24213),
            .I(N__24209));
    SRMux I__3731 (
            .O(N__24212),
            .I(N__24205));
    LocalMux I__3730 (
            .O(N__24209),
            .I(N__24201));
    SRMux I__3729 (
            .O(N__24208),
            .I(N__24198));
    LocalMux I__3728 (
            .O(N__24205),
            .I(N__24195));
    SRMux I__3727 (
            .O(N__24204),
            .I(N__24192));
    Span4Mux_v I__3726 (
            .O(N__24201),
            .I(N__24189));
    LocalMux I__3725 (
            .O(N__24198),
            .I(N__24184));
    Span4Mux_v I__3724 (
            .O(N__24195),
            .I(N__24184));
    LocalMux I__3723 (
            .O(N__24192),
            .I(N__24181));
    Sp12to4 I__3722 (
            .O(N__24189),
            .I(N__24178));
    Span4Mux_v I__3721 (
            .O(N__24184),
            .I(N__24175));
    Odrv12 I__3720 (
            .O(N__24181),
            .I(\nx.n7994 ));
    Odrv12 I__3719 (
            .O(N__24178),
            .I(\nx.n7994 ));
    Odrv4 I__3718 (
            .O(N__24175),
            .I(\nx.n7994 ));
    InMux I__3717 (
            .O(N__24168),
            .I(bfn_6_27_0_));
    InMux I__3716 (
            .O(N__24165),
            .I(\nx.n10819 ));
    InMux I__3715 (
            .O(N__24162),
            .I(\nx.n10820 ));
    InMux I__3714 (
            .O(N__24159),
            .I(N__24154));
    InMux I__3713 (
            .O(N__24158),
            .I(N__24151));
    InMux I__3712 (
            .O(N__24157),
            .I(N__24148));
    LocalMux I__3711 (
            .O(N__24154),
            .I(\nx.n1807 ));
    LocalMux I__3710 (
            .O(N__24151),
            .I(\nx.n1807 ));
    LocalMux I__3709 (
            .O(N__24148),
            .I(\nx.n1807 ));
    InMux I__3708 (
            .O(N__24141),
            .I(\nx.n10821 ));
    CascadeMux I__3707 (
            .O(N__24138),
            .I(N__24135));
    InMux I__3706 (
            .O(N__24135),
            .I(N__24130));
    InMux I__3705 (
            .O(N__24134),
            .I(N__24127));
    InMux I__3704 (
            .O(N__24133),
            .I(N__24124));
    LocalMux I__3703 (
            .O(N__24130),
            .I(N__24121));
    LocalMux I__3702 (
            .O(N__24127),
            .I(\nx.n1806 ));
    LocalMux I__3701 (
            .O(N__24124),
            .I(\nx.n1806 ));
    Odrv4 I__3700 (
            .O(N__24121),
            .I(\nx.n1806 ));
    InMux I__3699 (
            .O(N__24114),
            .I(\nx.n10822 ));
    InMux I__3698 (
            .O(N__24111),
            .I(\nx.n10823 ));
    InMux I__3697 (
            .O(N__24108),
            .I(\nx.n10632 ));
    InMux I__3696 (
            .O(N__24105),
            .I(N__24100));
    InMux I__3695 (
            .O(N__24104),
            .I(N__24097));
    InMux I__3694 (
            .O(N__24103),
            .I(N__24093));
    LocalMux I__3693 (
            .O(N__24100),
            .I(N__24087));
    LocalMux I__3692 (
            .O(N__24097),
            .I(N__24087));
    InMux I__3691 (
            .O(N__24096),
            .I(N__24084));
    LocalMux I__3690 (
            .O(N__24093),
            .I(N__24081));
    InMux I__3689 (
            .O(N__24092),
            .I(N__24078));
    Span4Mux_v I__3688 (
            .O(N__24087),
            .I(N__24075));
    LocalMux I__3687 (
            .O(N__24084),
            .I(N__24072));
    Span4Mux_h I__3686 (
            .O(N__24081),
            .I(N__24069));
    LocalMux I__3685 (
            .O(N__24078),
            .I(\nx.bit_ctr_21 ));
    Odrv4 I__3684 (
            .O(N__24075),
            .I(\nx.bit_ctr_21 ));
    Odrv12 I__3683 (
            .O(N__24072),
            .I(\nx.bit_ctr_21 ));
    Odrv4 I__3682 (
            .O(N__24069),
            .I(\nx.bit_ctr_21 ));
    InMux I__3681 (
            .O(N__24060),
            .I(\nx.n10633 ));
    InMux I__3680 (
            .O(N__24057),
            .I(\nx.n10634 ));
    InMux I__3679 (
            .O(N__24054),
            .I(N__24049));
    InMux I__3678 (
            .O(N__24053),
            .I(N__24045));
    InMux I__3677 (
            .O(N__24052),
            .I(N__24041));
    LocalMux I__3676 (
            .O(N__24049),
            .I(N__24038));
    InMux I__3675 (
            .O(N__24048),
            .I(N__24035));
    LocalMux I__3674 (
            .O(N__24045),
            .I(N__24032));
    InMux I__3673 (
            .O(N__24044),
            .I(N__24029));
    LocalMux I__3672 (
            .O(N__24041),
            .I(N__24024));
    Span4Mux_h I__3671 (
            .O(N__24038),
            .I(N__24024));
    LocalMux I__3670 (
            .O(N__24035),
            .I(N__24021));
    Span4Mux_h I__3669 (
            .O(N__24032),
            .I(N__24018));
    LocalMux I__3668 (
            .O(N__24029),
            .I(N__24013));
    Span4Mux_v I__3667 (
            .O(N__24024),
            .I(N__24013));
    Span4Mux_h I__3666 (
            .O(N__24021),
            .I(N__24010));
    Odrv4 I__3665 (
            .O(N__24018),
            .I(\nx.bit_ctr_23 ));
    Odrv4 I__3664 (
            .O(N__24013),
            .I(\nx.bit_ctr_23 ));
    Odrv4 I__3663 (
            .O(N__24010),
            .I(\nx.bit_ctr_23 ));
    InMux I__3662 (
            .O(N__24003),
            .I(\nx.n10635 ));
    InMux I__3661 (
            .O(N__24000),
            .I(N__23994));
    InMux I__3660 (
            .O(N__23999),
            .I(N__23991));
    InMux I__3659 (
            .O(N__23998),
            .I(N__23988));
    InMux I__3658 (
            .O(N__23997),
            .I(N__23984));
    LocalMux I__3657 (
            .O(N__23994),
            .I(N__23981));
    LocalMux I__3656 (
            .O(N__23991),
            .I(N__23976));
    LocalMux I__3655 (
            .O(N__23988),
            .I(N__23976));
    InMux I__3654 (
            .O(N__23987),
            .I(N__23973));
    LocalMux I__3653 (
            .O(N__23984),
            .I(N__23970));
    Span4Mux_h I__3652 (
            .O(N__23981),
            .I(N__23967));
    Span4Mux_v I__3651 (
            .O(N__23976),
            .I(N__23964));
    LocalMux I__3650 (
            .O(N__23973),
            .I(\nx.bit_ctr_24 ));
    Odrv4 I__3649 (
            .O(N__23970),
            .I(\nx.bit_ctr_24 ));
    Odrv4 I__3648 (
            .O(N__23967),
            .I(\nx.bit_ctr_24 ));
    Odrv4 I__3647 (
            .O(N__23964),
            .I(\nx.bit_ctr_24 ));
    InMux I__3646 (
            .O(N__23955),
            .I(bfn_6_26_0_));
    InMux I__3645 (
            .O(N__23952),
            .I(N__23947));
    InMux I__3644 (
            .O(N__23951),
            .I(N__23944));
    InMux I__3643 (
            .O(N__23950),
            .I(N__23941));
    LocalMux I__3642 (
            .O(N__23947),
            .I(N__23936));
    LocalMux I__3641 (
            .O(N__23944),
            .I(N__23933));
    LocalMux I__3640 (
            .O(N__23941),
            .I(N__23930));
    InMux I__3639 (
            .O(N__23940),
            .I(N__23927));
    InMux I__3638 (
            .O(N__23939),
            .I(N__23924));
    Span4Mux_h I__3637 (
            .O(N__23936),
            .I(N__23921));
    Span4Mux_v I__3636 (
            .O(N__23933),
            .I(N__23918));
    Span4Mux_v I__3635 (
            .O(N__23930),
            .I(N__23915));
    LocalMux I__3634 (
            .O(N__23927),
            .I(N__23912));
    LocalMux I__3633 (
            .O(N__23924),
            .I(\nx.bit_ctr_25 ));
    Odrv4 I__3632 (
            .O(N__23921),
            .I(\nx.bit_ctr_25 ));
    Odrv4 I__3631 (
            .O(N__23918),
            .I(\nx.bit_ctr_25 ));
    Odrv4 I__3630 (
            .O(N__23915),
            .I(\nx.bit_ctr_25 ));
    Odrv12 I__3629 (
            .O(N__23912),
            .I(\nx.bit_ctr_25 ));
    InMux I__3628 (
            .O(N__23901),
            .I(\nx.n10637 ));
    InMux I__3627 (
            .O(N__23898),
            .I(\nx.n10638 ));
    InMux I__3626 (
            .O(N__23895),
            .I(\nx.n10639 ));
    InMux I__3625 (
            .O(N__23892),
            .I(\nx.n10640 ));
    InMux I__3624 (
            .O(N__23889),
            .I(\nx.n10624 ));
    InMux I__3623 (
            .O(N__23886),
            .I(\nx.n10625 ));
    InMux I__3622 (
            .O(N__23883),
            .I(\nx.n10626 ));
    InMux I__3621 (
            .O(N__23880),
            .I(\nx.n10627 ));
    InMux I__3620 (
            .O(N__23877),
            .I(bfn_6_25_0_));
    InMux I__3619 (
            .O(N__23874),
            .I(\nx.n10629 ));
    InMux I__3618 (
            .O(N__23871),
            .I(\nx.n10630 ));
    InMux I__3617 (
            .O(N__23868),
            .I(N__23861));
    InMux I__3616 (
            .O(N__23867),
            .I(N__23858));
    InMux I__3615 (
            .O(N__23866),
            .I(N__23855));
    InMux I__3614 (
            .O(N__23865),
            .I(N__23852));
    InMux I__3613 (
            .O(N__23864),
            .I(N__23849));
    LocalMux I__3612 (
            .O(N__23861),
            .I(N__23844));
    LocalMux I__3611 (
            .O(N__23858),
            .I(N__23844));
    LocalMux I__3610 (
            .O(N__23855),
            .I(N__23841));
    LocalMux I__3609 (
            .O(N__23852),
            .I(\nx.bit_ctr_19 ));
    LocalMux I__3608 (
            .O(N__23849),
            .I(\nx.bit_ctr_19 ));
    Odrv4 I__3607 (
            .O(N__23844),
            .I(\nx.bit_ctr_19 ));
    Odrv4 I__3606 (
            .O(N__23841),
            .I(\nx.bit_ctr_19 ));
    InMux I__3605 (
            .O(N__23832),
            .I(\nx.n10631 ));
    InMux I__3604 (
            .O(N__23829),
            .I(N__23823));
    InMux I__3603 (
            .O(N__23828),
            .I(N__23820));
    InMux I__3602 (
            .O(N__23827),
            .I(N__23817));
    InMux I__3601 (
            .O(N__23826),
            .I(N__23814));
    LocalMux I__3600 (
            .O(N__23823),
            .I(N__23810));
    LocalMux I__3599 (
            .O(N__23820),
            .I(N__23805));
    LocalMux I__3598 (
            .O(N__23817),
            .I(N__23805));
    LocalMux I__3597 (
            .O(N__23814),
            .I(N__23802));
    InMux I__3596 (
            .O(N__23813),
            .I(N__23799));
    Span4Mux_v I__3595 (
            .O(N__23810),
            .I(N__23796));
    Span4Mux_v I__3594 (
            .O(N__23805),
            .I(N__23791));
    Span4Mux_v I__3593 (
            .O(N__23802),
            .I(N__23791));
    LocalMux I__3592 (
            .O(N__23799),
            .I(\nx.bit_ctr_20 ));
    Odrv4 I__3591 (
            .O(N__23796),
            .I(\nx.bit_ctr_20 ));
    Odrv4 I__3590 (
            .O(N__23791),
            .I(\nx.bit_ctr_20 ));
    InMux I__3589 (
            .O(N__23784),
            .I(\nx.n10614 ));
    InMux I__3588 (
            .O(N__23781),
            .I(\nx.n10615 ));
    InMux I__3587 (
            .O(N__23778),
            .I(\nx.n10616 ));
    InMux I__3586 (
            .O(N__23775),
            .I(\nx.n10617 ));
    InMux I__3585 (
            .O(N__23772),
            .I(\nx.n10618 ));
    InMux I__3584 (
            .O(N__23769),
            .I(\nx.n10619 ));
    InMux I__3583 (
            .O(N__23766),
            .I(bfn_6_24_0_));
    InMux I__3582 (
            .O(N__23763),
            .I(\nx.n10621 ));
    InMux I__3581 (
            .O(N__23760),
            .I(\nx.n10622 ));
    InMux I__3580 (
            .O(N__23757),
            .I(\nx.n10623 ));
    CascadeMux I__3579 (
            .O(N__23754),
            .I(\nx.n7899_cascade_ ));
    CascadeMux I__3578 (
            .O(N__23751),
            .I(N__23748));
    InMux I__3577 (
            .O(N__23748),
            .I(N__23745));
    LocalMux I__3576 (
            .O(N__23745),
            .I(\nx.n740 ));
    CascadeMux I__3575 (
            .O(N__23742),
            .I(\nx.n740_cascade_ ));
    CascadeMux I__3574 (
            .O(N__23739),
            .I(\nx.n11866_cascade_ ));
    CascadeMux I__3573 (
            .O(N__23736),
            .I(\nx.n838_cascade_ ));
    InMux I__3572 (
            .O(N__23733),
            .I(N__23730));
    LocalMux I__3571 (
            .O(N__23730),
            .I(N__23727));
    Span4Mux_h I__3570 (
            .O(N__23727),
            .I(N__23724));
    Span4Mux_h I__3569 (
            .O(N__23724),
            .I(N__23721));
    Odrv4 I__3568 (
            .O(N__23721),
            .I(n18_adj_815));
    InMux I__3567 (
            .O(N__23718),
            .I(N__23715));
    LocalMux I__3566 (
            .O(N__23715),
            .I(N__23712));
    Span4Mux_h I__3565 (
            .O(N__23712),
            .I(N__23708));
    InMux I__3564 (
            .O(N__23711),
            .I(N__23705));
    Span4Mux_h I__3563 (
            .O(N__23708),
            .I(N__23702));
    LocalMux I__3562 (
            .O(N__23705),
            .I(delay_counter_31));
    Odrv4 I__3561 (
            .O(N__23702),
            .I(delay_counter_31));
    CascadeMux I__3560 (
            .O(N__23697),
            .I(N__23694));
    InMux I__3559 (
            .O(N__23694),
            .I(N__23691));
    LocalMux I__3558 (
            .O(N__23691),
            .I(N__23688));
    Span4Mux_h I__3557 (
            .O(N__23688),
            .I(N__23685));
    Odrv4 I__3556 (
            .O(N__23685),
            .I(n19_adj_814));
    InMux I__3555 (
            .O(N__23682),
            .I(N__23679));
    LocalMux I__3554 (
            .O(N__23679),
            .I(N__23676));
    Span4Mux_h I__3553 (
            .O(N__23676),
            .I(N__23673));
    Odrv4 I__3552 (
            .O(N__23673),
            .I(n17_adj_816));
    InMux I__3551 (
            .O(N__23670),
            .I(bfn_6_23_0_));
    InMux I__3550 (
            .O(N__23667),
            .I(\nx.n10613 ));
    InMux I__3549 (
            .O(N__23664),
            .I(N__23661));
    LocalMux I__3548 (
            .O(N__23661),
            .I(N__23658));
    Span12Mux_s11_v I__3547 (
            .O(N__23658),
            .I(N__23655));
    Odrv12 I__3546 (
            .O(N__23655),
            .I(\nx.n5 ));
    CascadeMux I__3545 (
            .O(N__23652),
            .I(N__23648));
    CascadeMux I__3544 (
            .O(N__23651),
            .I(N__23645));
    InMux I__3543 (
            .O(N__23648),
            .I(N__23642));
    InMux I__3542 (
            .O(N__23645),
            .I(N__23639));
    LocalMux I__3541 (
            .O(N__23642),
            .I(\nx.n1007 ));
    LocalMux I__3540 (
            .O(N__23639),
            .I(\nx.n1007 ));
    InMux I__3539 (
            .O(N__23634),
            .I(N__23631));
    LocalMux I__3538 (
            .O(N__23631),
            .I(\nx.n1075 ));
    InMux I__3537 (
            .O(N__23628),
            .I(N__23624));
    CascadeMux I__3536 (
            .O(N__23627),
            .I(N__23620));
    LocalMux I__3535 (
            .O(N__23624),
            .I(N__23617));
    InMux I__3534 (
            .O(N__23623),
            .I(N__23614));
    InMux I__3533 (
            .O(N__23620),
            .I(N__23611));
    Odrv4 I__3532 (
            .O(N__23617),
            .I(\nx.n1107 ));
    LocalMux I__3531 (
            .O(N__23614),
            .I(\nx.n1107 ));
    LocalMux I__3530 (
            .O(N__23611),
            .I(\nx.n1107 ));
    CascadeMux I__3529 (
            .O(N__23604),
            .I(N__23600));
    CascadeMux I__3528 (
            .O(N__23603),
            .I(N__23597));
    InMux I__3527 (
            .O(N__23600),
            .I(N__23594));
    InMux I__3526 (
            .O(N__23597),
            .I(N__23591));
    LocalMux I__3525 (
            .O(N__23594),
            .I(\nx.n1005 ));
    LocalMux I__3524 (
            .O(N__23591),
            .I(\nx.n1005 ));
    CascadeMux I__3523 (
            .O(N__23586),
            .I(\nx.n1005_cascade_ ));
    CascadeMux I__3522 (
            .O(N__23583),
            .I(N__23578));
    InMux I__3521 (
            .O(N__23582),
            .I(N__23575));
    InMux I__3520 (
            .O(N__23581),
            .I(N__23572));
    InMux I__3519 (
            .O(N__23578),
            .I(N__23569));
    LocalMux I__3518 (
            .O(N__23575),
            .I(\nx.n1009 ));
    LocalMux I__3517 (
            .O(N__23572),
            .I(\nx.n1009 ));
    LocalMux I__3516 (
            .O(N__23569),
            .I(\nx.n1009 ));
    CascadeMux I__3515 (
            .O(N__23562),
            .I(\nx.n7_adj_690_cascade_ ));
    CascadeMux I__3514 (
            .O(N__23559),
            .I(N__23555));
    CascadeMux I__3513 (
            .O(N__23558),
            .I(N__23549));
    InMux I__3512 (
            .O(N__23555),
            .I(N__23545));
    InMux I__3511 (
            .O(N__23554),
            .I(N__23542));
    InMux I__3510 (
            .O(N__23553),
            .I(N__23533));
    InMux I__3509 (
            .O(N__23552),
            .I(N__23533));
    InMux I__3508 (
            .O(N__23549),
            .I(N__23533));
    InMux I__3507 (
            .O(N__23548),
            .I(N__23533));
    LocalMux I__3506 (
            .O(N__23545),
            .I(\nx.n1037 ));
    LocalMux I__3505 (
            .O(N__23542),
            .I(\nx.n1037 ));
    LocalMux I__3504 (
            .O(N__23533),
            .I(\nx.n1037 ));
    CascadeMux I__3503 (
            .O(N__23526),
            .I(\nx.n1037_cascade_ ));
    InMux I__3502 (
            .O(N__23523),
            .I(N__23520));
    LocalMux I__3501 (
            .O(N__23520),
            .I(\nx.n1073 ));
    InMux I__3500 (
            .O(N__23517),
            .I(N__23513));
    CascadeMux I__3499 (
            .O(N__23516),
            .I(N__23510));
    LocalMux I__3498 (
            .O(N__23513),
            .I(N__23506));
    InMux I__3497 (
            .O(N__23510),
            .I(N__23503));
    InMux I__3496 (
            .O(N__23509),
            .I(N__23500));
    Odrv4 I__3495 (
            .O(N__23506),
            .I(\nx.n1105 ));
    LocalMux I__3494 (
            .O(N__23503),
            .I(\nx.n1105 ));
    LocalMux I__3493 (
            .O(N__23500),
            .I(\nx.n1105 ));
    InMux I__3492 (
            .O(N__23493),
            .I(N__23489));
    InMux I__3491 (
            .O(N__23492),
            .I(N__23486));
    LocalMux I__3490 (
            .O(N__23489),
            .I(N__23483));
    LocalMux I__3489 (
            .O(N__23486),
            .I(N__23466));
    Span4Mux_h I__3488 (
            .O(N__23483),
            .I(N__23463));
    InMux I__3487 (
            .O(N__23482),
            .I(N__23458));
    InMux I__3486 (
            .O(N__23481),
            .I(N__23458));
    InMux I__3485 (
            .O(N__23480),
            .I(N__23453));
    InMux I__3484 (
            .O(N__23479),
            .I(N__23453));
    InMux I__3483 (
            .O(N__23478),
            .I(N__23450));
    InMux I__3482 (
            .O(N__23477),
            .I(N__23445));
    InMux I__3481 (
            .O(N__23476),
            .I(N__23445));
    InMux I__3480 (
            .O(N__23475),
            .I(N__23440));
    InMux I__3479 (
            .O(N__23474),
            .I(N__23440));
    InMux I__3478 (
            .O(N__23473),
            .I(N__23433));
    InMux I__3477 (
            .O(N__23472),
            .I(N__23433));
    InMux I__3476 (
            .O(N__23471),
            .I(N__23433));
    InMux I__3475 (
            .O(N__23470),
            .I(N__23428));
    InMux I__3474 (
            .O(N__23469),
            .I(N__23428));
    Odrv4 I__3473 (
            .O(N__23466),
            .I(state_1_adj_791));
    Odrv4 I__3472 (
            .O(N__23463),
            .I(state_1_adj_791));
    LocalMux I__3471 (
            .O(N__23458),
            .I(state_1_adj_791));
    LocalMux I__3470 (
            .O(N__23453),
            .I(state_1_adj_791));
    LocalMux I__3469 (
            .O(N__23450),
            .I(state_1_adj_791));
    LocalMux I__3468 (
            .O(N__23445),
            .I(state_1_adj_791));
    LocalMux I__3467 (
            .O(N__23440),
            .I(state_1_adj_791));
    LocalMux I__3466 (
            .O(N__23433),
            .I(state_1_adj_791));
    LocalMux I__3465 (
            .O(N__23428),
            .I(state_1_adj_791));
    CascadeMux I__3464 (
            .O(N__23409),
            .I(\nx.n3901_cascade_ ));
    InMux I__3463 (
            .O(N__23406),
            .I(N__23403));
    LocalMux I__3462 (
            .O(N__23403),
            .I(N__23400));
    Odrv4 I__3461 (
            .O(N__23400),
            .I(\nx.n13435 ));
    InMux I__3460 (
            .O(N__23397),
            .I(N__23394));
    LocalMux I__3459 (
            .O(N__23394),
            .I(\nx.n1077 ));
    InMux I__3458 (
            .O(N__23391),
            .I(bfn_6_20_0_));
    CascadeMux I__3457 (
            .O(N__23388),
            .I(N__23385));
    InMux I__3456 (
            .O(N__23385),
            .I(N__23382));
    LocalMux I__3455 (
            .O(N__23382),
            .I(\nx.n1076 ));
    InMux I__3454 (
            .O(N__23379),
            .I(\nx.n10743 ));
    InMux I__3453 (
            .O(N__23376),
            .I(\nx.n10744 ));
    InMux I__3452 (
            .O(N__23373),
            .I(N__23370));
    LocalMux I__3451 (
            .O(N__23370),
            .I(\nx.n1074 ));
    InMux I__3450 (
            .O(N__23367),
            .I(\nx.n10745 ));
    InMux I__3449 (
            .O(N__23364),
            .I(\nx.n10746 ));
    InMux I__3448 (
            .O(N__23361),
            .I(N__23358));
    LocalMux I__3447 (
            .O(N__23358),
            .I(\nx.n1072 ));
    InMux I__3446 (
            .O(N__23355),
            .I(\nx.n10747 ));
    InMux I__3445 (
            .O(N__23352),
            .I(\nx.n10748 ));
    CascadeMux I__3444 (
            .O(N__23349),
            .I(N__23345));
    InMux I__3443 (
            .O(N__23348),
            .I(N__23342));
    InMux I__3442 (
            .O(N__23345),
            .I(N__23339));
    LocalMux I__3441 (
            .O(N__23342),
            .I(N__23336));
    LocalMux I__3440 (
            .O(N__23339),
            .I(\nx.n1103 ));
    Odrv4 I__3439 (
            .O(N__23336),
            .I(\nx.n1103 ));
    InMux I__3438 (
            .O(N__23331),
            .I(N__23328));
    LocalMux I__3437 (
            .O(N__23328),
            .I(N__23324));
    CascadeMux I__3436 (
            .O(N__23327),
            .I(N__23320));
    Span4Mux_h I__3435 (
            .O(N__23324),
            .I(N__23317));
    InMux I__3434 (
            .O(N__23323),
            .I(N__23314));
    InMux I__3433 (
            .O(N__23320),
            .I(N__23311));
    Odrv4 I__3432 (
            .O(N__23317),
            .I(timer_26));
    LocalMux I__3431 (
            .O(N__23314),
            .I(timer_26));
    LocalMux I__3430 (
            .O(N__23311),
            .I(timer_26));
    InMux I__3429 (
            .O(N__23304),
            .I(N__23298));
    InMux I__3428 (
            .O(N__23303),
            .I(N__23298));
    LocalMux I__3427 (
            .O(N__23298),
            .I(neo_pixel_transmitter_t0_26));
    InMux I__3426 (
            .O(N__23295),
            .I(N__23292));
    LocalMux I__3425 (
            .O(N__23292),
            .I(N__23289));
    Span4Mux_v I__3424 (
            .O(N__23289),
            .I(N__23286));
    Odrv4 I__3423 (
            .O(N__23286),
            .I(\nx.n7 ));
    InMux I__3422 (
            .O(N__23283),
            .I(N__23280));
    LocalMux I__3421 (
            .O(N__23280),
            .I(\nx.n10_adj_760 ));
    CascadeMux I__3420 (
            .O(N__23277),
            .I(N__23274));
    InMux I__3419 (
            .O(N__23274),
            .I(N__23271));
    LocalMux I__3418 (
            .O(N__23271),
            .I(N__23268));
    Span4Mux_h I__3417 (
            .O(N__23268),
            .I(N__23265));
    Odrv4 I__3416 (
            .O(N__23265),
            .I(n12_adj_844));
    InMux I__3415 (
            .O(N__23262),
            .I(N__23256));
    InMux I__3414 (
            .O(N__23261),
            .I(N__23251));
    InMux I__3413 (
            .O(N__23260),
            .I(N__23251));
    CascadeMux I__3412 (
            .O(N__23259),
            .I(N__23245));
    LocalMux I__3411 (
            .O(N__23256),
            .I(N__23240));
    LocalMux I__3410 (
            .O(N__23251),
            .I(N__23237));
    InMux I__3409 (
            .O(N__23250),
            .I(N__23234));
    InMux I__3408 (
            .O(N__23249),
            .I(N__23231));
    InMux I__3407 (
            .O(N__23248),
            .I(N__23222));
    InMux I__3406 (
            .O(N__23245),
            .I(N__23222));
    InMux I__3405 (
            .O(N__23244),
            .I(N__23222));
    InMux I__3404 (
            .O(N__23243),
            .I(N__23222));
    Span4Mux_v I__3403 (
            .O(N__23240),
            .I(N__23219));
    Span4Mux_h I__3402 (
            .O(N__23237),
            .I(N__23216));
    LocalMux I__3401 (
            .O(N__23234),
            .I(\nx.start ));
    LocalMux I__3400 (
            .O(N__23231),
            .I(\nx.start ));
    LocalMux I__3399 (
            .O(N__23222),
            .I(\nx.start ));
    Odrv4 I__3398 (
            .O(N__23219),
            .I(\nx.start ));
    Odrv4 I__3397 (
            .O(N__23216),
            .I(\nx.start ));
    InMux I__3396 (
            .O(N__23205),
            .I(N__23200));
    InMux I__3395 (
            .O(N__23204),
            .I(N__23197));
    InMux I__3394 (
            .O(N__23203),
            .I(N__23194));
    LocalMux I__3393 (
            .O(N__23200),
            .I(\nx.n11908 ));
    LocalMux I__3392 (
            .O(N__23197),
            .I(\nx.n11908 ));
    LocalMux I__3391 (
            .O(N__23194),
            .I(\nx.n11908 ));
    CascadeMux I__3390 (
            .O(N__23187),
            .I(N__23184));
    InMux I__3389 (
            .O(N__23184),
            .I(N__23178));
    InMux I__3388 (
            .O(N__23183),
            .I(N__23175));
    InMux I__3387 (
            .O(N__23182),
            .I(N__23170));
    InMux I__3386 (
            .O(N__23181),
            .I(N__23170));
    LocalMux I__3385 (
            .O(N__23178),
            .I(N__23161));
    LocalMux I__3384 (
            .O(N__23175),
            .I(N__23161));
    LocalMux I__3383 (
            .O(N__23170),
            .I(N__23161));
    InMux I__3382 (
            .O(N__23169),
            .I(N__23158));
    InMux I__3381 (
            .O(N__23168),
            .I(N__23155));
    Span4Mux_h I__3380 (
            .O(N__23161),
            .I(N__23152));
    LocalMux I__3379 (
            .O(N__23158),
            .I(N__23149));
    LocalMux I__3378 (
            .O(N__23155),
            .I(\nx.n7564 ));
    Odrv4 I__3377 (
            .O(N__23152),
            .I(\nx.n7564 ));
    Odrv12 I__3376 (
            .O(N__23149),
            .I(\nx.n7564 ));
    InMux I__3375 (
            .O(N__23142),
            .I(N__23138));
    InMux I__3374 (
            .O(N__23141),
            .I(N__23135));
    LocalMux I__3373 (
            .O(N__23138),
            .I(update_color));
    LocalMux I__3372 (
            .O(N__23135),
            .I(update_color));
    CascadeMux I__3371 (
            .O(N__23130),
            .I(\nx.n13436_cascade_ ));
    InMux I__3370 (
            .O(N__23127),
            .I(N__23124));
    LocalMux I__3369 (
            .O(N__23124),
            .I(\nx.n3901 ));
    InMux I__3368 (
            .O(N__23121),
            .I(N__23118));
    LocalMux I__3367 (
            .O(N__23118),
            .I(N__23115));
    Odrv4 I__3366 (
            .O(N__23115),
            .I(\nx.n16_adj_766 ));
    InMux I__3365 (
            .O(N__23112),
            .I(N__23107));
    InMux I__3364 (
            .O(N__23111),
            .I(N__23104));
    InMux I__3363 (
            .O(N__23110),
            .I(N__23101));
    LocalMux I__3362 (
            .O(N__23107),
            .I(N__23094));
    LocalMux I__3361 (
            .O(N__23104),
            .I(N__23094));
    LocalMux I__3360 (
            .O(N__23101),
            .I(N__23094));
    Odrv12 I__3359 (
            .O(N__23094),
            .I(\nx.n1702 ));
    CascadeMux I__3358 (
            .O(N__23091),
            .I(\nx.n22_adj_774_cascade_ ));
    InMux I__3357 (
            .O(N__23088),
            .I(N__23083));
    InMux I__3356 (
            .O(N__23087),
            .I(N__23080));
    InMux I__3355 (
            .O(N__23086),
            .I(N__23077));
    LocalMux I__3354 (
            .O(N__23083),
            .I(N__23074));
    LocalMux I__3353 (
            .O(N__23080),
            .I(N__23069));
    LocalMux I__3352 (
            .O(N__23077),
            .I(N__23069));
    Odrv4 I__3351 (
            .O(N__23074),
            .I(\nx.n1698 ));
    Odrv4 I__3350 (
            .O(N__23069),
            .I(\nx.n1698 ));
    InMux I__3349 (
            .O(N__23064),
            .I(N__23059));
    InMux I__3348 (
            .O(N__23063),
            .I(N__23056));
    InMux I__3347 (
            .O(N__23062),
            .I(N__23053));
    LocalMux I__3346 (
            .O(N__23059),
            .I(N__23046));
    LocalMux I__3345 (
            .O(N__23056),
            .I(N__23046));
    LocalMux I__3344 (
            .O(N__23053),
            .I(N__23046));
    Odrv4 I__3343 (
            .O(N__23046),
            .I(\nx.n1699 ));
    InMux I__3342 (
            .O(N__23043),
            .I(N__23038));
    InMux I__3341 (
            .O(N__23042),
            .I(N__23035));
    InMux I__3340 (
            .O(N__23041),
            .I(N__23032));
    LocalMux I__3339 (
            .O(N__23038),
            .I(N__23029));
    LocalMux I__3338 (
            .O(N__23035),
            .I(N__23026));
    LocalMux I__3337 (
            .O(N__23032),
            .I(N__23023));
    Odrv4 I__3336 (
            .O(N__23029),
            .I(\nx.n1697 ));
    Odrv12 I__3335 (
            .O(N__23026),
            .I(\nx.n1697 ));
    Odrv4 I__3334 (
            .O(N__23023),
            .I(\nx.n1697 ));
    CascadeMux I__3333 (
            .O(N__23016),
            .I(\nx.n24_adj_776_cascade_ ));
    InMux I__3332 (
            .O(N__23013),
            .I(N__23010));
    LocalMux I__3331 (
            .O(N__23010),
            .I(N__23007));
    Odrv4 I__3330 (
            .O(N__23007),
            .I(\nx.n20_adj_775 ));
    CascadeMux I__3329 (
            .O(N__23004),
            .I(N__22990));
    CascadeMux I__3328 (
            .O(N__23003),
            .I(N__22987));
    CascadeMux I__3327 (
            .O(N__23002),
            .I(N__22984));
    CascadeMux I__3326 (
            .O(N__23001),
            .I(N__22981));
    CascadeMux I__3325 (
            .O(N__23000),
            .I(N__22978));
    CascadeMux I__3324 (
            .O(N__22999),
            .I(N__22975));
    CascadeMux I__3323 (
            .O(N__22998),
            .I(N__22972));
    CascadeMux I__3322 (
            .O(N__22997),
            .I(N__22969));
    CascadeMux I__3321 (
            .O(N__22996),
            .I(N__22966));
    CascadeMux I__3320 (
            .O(N__22995),
            .I(N__22963));
    CascadeMux I__3319 (
            .O(N__22994),
            .I(N__22960));
    CascadeMux I__3318 (
            .O(N__22993),
            .I(N__22957));
    InMux I__3317 (
            .O(N__22990),
            .I(N__22950));
    InMux I__3316 (
            .O(N__22987),
            .I(N__22950));
    InMux I__3315 (
            .O(N__22984),
            .I(N__22950));
    InMux I__3314 (
            .O(N__22981),
            .I(N__22943));
    InMux I__3313 (
            .O(N__22978),
            .I(N__22943));
    InMux I__3312 (
            .O(N__22975),
            .I(N__22943));
    InMux I__3311 (
            .O(N__22972),
            .I(N__22936));
    InMux I__3310 (
            .O(N__22969),
            .I(N__22936));
    InMux I__3309 (
            .O(N__22966),
            .I(N__22936));
    InMux I__3308 (
            .O(N__22963),
            .I(N__22929));
    InMux I__3307 (
            .O(N__22960),
            .I(N__22929));
    InMux I__3306 (
            .O(N__22957),
            .I(N__22929));
    LocalMux I__3305 (
            .O(N__22950),
            .I(N__22924));
    LocalMux I__3304 (
            .O(N__22943),
            .I(N__22924));
    LocalMux I__3303 (
            .O(N__22936),
            .I(\nx.n1730 ));
    LocalMux I__3302 (
            .O(N__22929),
            .I(\nx.n1730 ));
    Odrv4 I__3301 (
            .O(N__22924),
            .I(\nx.n1730 ));
    CascadeMux I__3300 (
            .O(N__22917),
            .I(\nx.n1730_cascade_ ));
    CascadeMux I__3299 (
            .O(N__22914),
            .I(N__22910));
    CascadeMux I__3298 (
            .O(N__22913),
            .I(N__22907));
    InMux I__3297 (
            .O(N__22910),
            .I(N__22904));
    InMux I__3296 (
            .O(N__22907),
            .I(N__22901));
    LocalMux I__3295 (
            .O(N__22904),
            .I(N__22896));
    LocalMux I__3294 (
            .O(N__22901),
            .I(N__22896));
    Odrv4 I__3293 (
            .O(N__22896),
            .I(\nx.n13601 ));
    InMux I__3292 (
            .O(N__22893),
            .I(N__22890));
    LocalMux I__3291 (
            .O(N__22890),
            .I(n11972));
    InMux I__3290 (
            .O(N__22887),
            .I(N__22884));
    LocalMux I__3289 (
            .O(N__22884),
            .I(\nx.n13514 ));
    CascadeMux I__3288 (
            .O(N__22881),
            .I(N__22878));
    InMux I__3287 (
            .O(N__22878),
            .I(N__22875));
    LocalMux I__3286 (
            .O(N__22875),
            .I(\nx.n13513 ));
    InMux I__3285 (
            .O(N__22872),
            .I(N__22869));
    LocalMux I__3284 (
            .O(N__22869),
            .I(N__22865));
    InMux I__3283 (
            .O(N__22868),
            .I(N__22862));
    Odrv4 I__3282 (
            .O(N__22865),
            .I(\nx.n7598 ));
    LocalMux I__3281 (
            .O(N__22862),
            .I(\nx.n7598 ));
    InMux I__3280 (
            .O(N__22857),
            .I(N__22849));
    InMux I__3279 (
            .O(N__22856),
            .I(N__22849));
    InMux I__3278 (
            .O(N__22855),
            .I(N__22846));
    InMux I__3277 (
            .O(N__22854),
            .I(N__22843));
    LocalMux I__3276 (
            .O(N__22849),
            .I(\nx.n11113 ));
    LocalMux I__3275 (
            .O(N__22846),
            .I(\nx.n11113 ));
    LocalMux I__3274 (
            .O(N__22843),
            .I(\nx.n11113 ));
    CascadeMux I__3273 (
            .O(N__22836),
            .I(\nx.n7598_cascade_ ));
    InMux I__3272 (
            .O(N__22833),
            .I(bfn_5_28_0_));
    InMux I__3271 (
            .O(N__22830),
            .I(N__22826));
    InMux I__3270 (
            .O(N__22829),
            .I(N__22823));
    LocalMux I__3269 (
            .O(N__22826),
            .I(N__22817));
    LocalMux I__3268 (
            .O(N__22823),
            .I(N__22817));
    InMux I__3267 (
            .O(N__22822),
            .I(N__22814));
    Odrv4 I__3266 (
            .O(N__22817),
            .I(\nx.n1701 ));
    LocalMux I__3265 (
            .O(N__22814),
            .I(\nx.n1701 ));
    InMux I__3264 (
            .O(N__22809),
            .I(\nx.n10814 ));
    InMux I__3263 (
            .O(N__22806),
            .I(\nx.n10815 ));
    InMux I__3262 (
            .O(N__22803),
            .I(\nx.n10816 ));
    InMux I__3261 (
            .O(N__22800),
            .I(\nx.n10817 ));
    InMux I__3260 (
            .O(N__22797),
            .I(\nx.n10818 ));
    InMux I__3259 (
            .O(N__22794),
            .I(N__22791));
    LocalMux I__3258 (
            .O(N__22791),
            .I(N__22788));
    Span4Mux_v I__3257 (
            .O(N__22788),
            .I(N__22783));
    InMux I__3256 (
            .O(N__22787),
            .I(N__22780));
    InMux I__3255 (
            .O(N__22786),
            .I(N__22777));
    Span4Mux_h I__3254 (
            .O(N__22783),
            .I(N__22772));
    LocalMux I__3253 (
            .O(N__22780),
            .I(N__22772));
    LocalMux I__3252 (
            .O(N__22777),
            .I(N__22769));
    Odrv4 I__3251 (
            .O(N__22772),
            .I(\nx.n1703 ));
    Odrv12 I__3250 (
            .O(N__22769),
            .I(\nx.n1703 ));
    InMux I__3249 (
            .O(N__22764),
            .I(N__22759));
    InMux I__3248 (
            .O(N__22763),
            .I(N__22756));
    InMux I__3247 (
            .O(N__22762),
            .I(N__22753));
    LocalMux I__3246 (
            .O(N__22759),
            .I(N__22746));
    LocalMux I__3245 (
            .O(N__22756),
            .I(N__22746));
    LocalMux I__3244 (
            .O(N__22753),
            .I(N__22746));
    Odrv12 I__3243 (
            .O(N__22746),
            .I(\nx.n1706 ));
    CascadeMux I__3242 (
            .O(N__22743),
            .I(N__22738));
    InMux I__3241 (
            .O(N__22742),
            .I(N__22735));
    InMux I__3240 (
            .O(N__22741),
            .I(N__22732));
    InMux I__3239 (
            .O(N__22738),
            .I(N__22729));
    LocalMux I__3238 (
            .O(N__22735),
            .I(N__22724));
    LocalMux I__3237 (
            .O(N__22732),
            .I(N__22724));
    LocalMux I__3236 (
            .O(N__22729),
            .I(N__22721));
    Odrv4 I__3235 (
            .O(N__22724),
            .I(\nx.n1705 ));
    Odrv12 I__3234 (
            .O(N__22721),
            .I(\nx.n1705 ));
    InMux I__3233 (
            .O(N__22716),
            .I(N__22711));
    InMux I__3232 (
            .O(N__22715),
            .I(N__22708));
    InMux I__3231 (
            .O(N__22714),
            .I(N__22705));
    LocalMux I__3230 (
            .O(N__22711),
            .I(N__22698));
    LocalMux I__3229 (
            .O(N__22708),
            .I(N__22698));
    LocalMux I__3228 (
            .O(N__22705),
            .I(N__22698));
    Odrv12 I__3227 (
            .O(N__22698),
            .I(\nx.n1700 ));
    InMux I__3226 (
            .O(N__22695),
            .I(bfn_5_27_0_));
    InMux I__3225 (
            .O(N__22692),
            .I(N__22687));
    InMux I__3224 (
            .O(N__22691),
            .I(N__22684));
    CascadeMux I__3223 (
            .O(N__22690),
            .I(N__22681));
    LocalMux I__3222 (
            .O(N__22687),
            .I(N__22676));
    LocalMux I__3221 (
            .O(N__22684),
            .I(N__22676));
    InMux I__3220 (
            .O(N__22681),
            .I(N__22673));
    Odrv12 I__3219 (
            .O(N__22676),
            .I(\nx.n1709 ));
    LocalMux I__3218 (
            .O(N__22673),
            .I(\nx.n1709 ));
    InMux I__3217 (
            .O(N__22668),
            .I(\nx.n10806 ));
    InMux I__3216 (
            .O(N__22665),
            .I(N__22662));
    LocalMux I__3215 (
            .O(N__22662),
            .I(N__22658));
    InMux I__3214 (
            .O(N__22661),
            .I(N__22655));
    Span4Mux_h I__3213 (
            .O(N__22658),
            .I(N__22649));
    LocalMux I__3212 (
            .O(N__22655),
            .I(N__22649));
    InMux I__3211 (
            .O(N__22654),
            .I(N__22646));
    Odrv4 I__3210 (
            .O(N__22649),
            .I(\nx.n1708 ));
    LocalMux I__3209 (
            .O(N__22646),
            .I(\nx.n1708 ));
    InMux I__3208 (
            .O(N__22641),
            .I(\nx.n10807 ));
    InMux I__3207 (
            .O(N__22638),
            .I(N__22634));
    InMux I__3206 (
            .O(N__22637),
            .I(N__22631));
    LocalMux I__3205 (
            .O(N__22634),
            .I(N__22625));
    LocalMux I__3204 (
            .O(N__22631),
            .I(N__22625));
    InMux I__3203 (
            .O(N__22630),
            .I(N__22622));
    Odrv4 I__3202 (
            .O(N__22625),
            .I(\nx.n1707 ));
    LocalMux I__3201 (
            .O(N__22622),
            .I(\nx.n1707 ));
    InMux I__3200 (
            .O(N__22617),
            .I(\nx.n10808 ));
    InMux I__3199 (
            .O(N__22614),
            .I(\nx.n10809 ));
    InMux I__3198 (
            .O(N__22611),
            .I(\nx.n10810 ));
    InMux I__3197 (
            .O(N__22608),
            .I(N__22603));
    InMux I__3196 (
            .O(N__22607),
            .I(N__22600));
    CascadeMux I__3195 (
            .O(N__22606),
            .I(N__22597));
    LocalMux I__3194 (
            .O(N__22603),
            .I(N__22592));
    LocalMux I__3193 (
            .O(N__22600),
            .I(N__22592));
    InMux I__3192 (
            .O(N__22597),
            .I(N__22589));
    Odrv4 I__3191 (
            .O(N__22592),
            .I(\nx.n1704 ));
    LocalMux I__3190 (
            .O(N__22589),
            .I(\nx.n1704 ));
    InMux I__3189 (
            .O(N__22584),
            .I(\nx.n10811 ));
    InMux I__3188 (
            .O(N__22581),
            .I(\nx.n10812 ));
    InMux I__3187 (
            .O(N__22578),
            .I(N__22573));
    InMux I__3186 (
            .O(N__22577),
            .I(N__22570));
    InMux I__3185 (
            .O(N__22576),
            .I(N__22567));
    LocalMux I__3184 (
            .O(N__22573),
            .I(\nx.n1605 ));
    LocalMux I__3183 (
            .O(N__22570),
            .I(\nx.n1605 ));
    LocalMux I__3182 (
            .O(N__22567),
            .I(\nx.n1605 ));
    InMux I__3181 (
            .O(N__22560),
            .I(\nx.n10798 ));
    InMux I__3180 (
            .O(N__22557),
            .I(N__22552));
    InMux I__3179 (
            .O(N__22556),
            .I(N__22549));
    InMux I__3178 (
            .O(N__22555),
            .I(N__22546));
    LocalMux I__3177 (
            .O(N__22552),
            .I(\nx.n1604 ));
    LocalMux I__3176 (
            .O(N__22549),
            .I(\nx.n1604 ));
    LocalMux I__3175 (
            .O(N__22546),
            .I(\nx.n1604 ));
    InMux I__3174 (
            .O(N__22539),
            .I(\nx.n10799 ));
    CascadeMux I__3173 (
            .O(N__22536),
            .I(N__22531));
    InMux I__3172 (
            .O(N__22535),
            .I(N__22528));
    InMux I__3171 (
            .O(N__22534),
            .I(N__22525));
    InMux I__3170 (
            .O(N__22531),
            .I(N__22522));
    LocalMux I__3169 (
            .O(N__22528),
            .I(\nx.n1603 ));
    LocalMux I__3168 (
            .O(N__22525),
            .I(\nx.n1603 ));
    LocalMux I__3167 (
            .O(N__22522),
            .I(\nx.n1603 ));
    InMux I__3166 (
            .O(N__22515),
            .I(\nx.n10800 ));
    CascadeMux I__3165 (
            .O(N__22512),
            .I(N__22507));
    InMux I__3164 (
            .O(N__22511),
            .I(N__22504));
    InMux I__3163 (
            .O(N__22510),
            .I(N__22501));
    InMux I__3162 (
            .O(N__22507),
            .I(N__22498));
    LocalMux I__3161 (
            .O(N__22504),
            .I(\nx.n1602 ));
    LocalMux I__3160 (
            .O(N__22501),
            .I(\nx.n1602 ));
    LocalMux I__3159 (
            .O(N__22498),
            .I(\nx.n1602 ));
    InMux I__3158 (
            .O(N__22491),
            .I(bfn_5_26_0_));
    InMux I__3157 (
            .O(N__22488),
            .I(N__22484));
    InMux I__3156 (
            .O(N__22487),
            .I(N__22480));
    LocalMux I__3155 (
            .O(N__22484),
            .I(N__22477));
    InMux I__3154 (
            .O(N__22483),
            .I(N__22474));
    LocalMux I__3153 (
            .O(N__22480),
            .I(\nx.n1601 ));
    Odrv4 I__3152 (
            .O(N__22477),
            .I(\nx.n1601 ));
    LocalMux I__3151 (
            .O(N__22474),
            .I(\nx.n1601 ));
    InMux I__3150 (
            .O(N__22467),
            .I(\nx.n10802 ));
    InMux I__3149 (
            .O(N__22464),
            .I(N__22459));
    InMux I__3148 (
            .O(N__22463),
            .I(N__22456));
    CascadeMux I__3147 (
            .O(N__22462),
            .I(N__22453));
    LocalMux I__3146 (
            .O(N__22459),
            .I(N__22448));
    LocalMux I__3145 (
            .O(N__22456),
            .I(N__22448));
    InMux I__3144 (
            .O(N__22453),
            .I(N__22445));
    Odrv4 I__3143 (
            .O(N__22448),
            .I(\nx.n1600 ));
    LocalMux I__3142 (
            .O(N__22445),
            .I(\nx.n1600 ));
    InMux I__3141 (
            .O(N__22440),
            .I(\nx.n10803 ));
    InMux I__3140 (
            .O(N__22437),
            .I(N__22432));
    InMux I__3139 (
            .O(N__22436),
            .I(N__22429));
    InMux I__3138 (
            .O(N__22435),
            .I(N__22426));
    LocalMux I__3137 (
            .O(N__22432),
            .I(\nx.n1599 ));
    LocalMux I__3136 (
            .O(N__22429),
            .I(\nx.n1599 ));
    LocalMux I__3135 (
            .O(N__22426),
            .I(\nx.n1599 ));
    InMux I__3134 (
            .O(N__22419),
            .I(\nx.n10804 ));
    InMux I__3133 (
            .O(N__22416),
            .I(N__22411));
    InMux I__3132 (
            .O(N__22415),
            .I(N__22408));
    InMux I__3131 (
            .O(N__22414),
            .I(N__22405));
    LocalMux I__3130 (
            .O(N__22411),
            .I(N__22402));
    LocalMux I__3129 (
            .O(N__22408),
            .I(\nx.n1598 ));
    LocalMux I__3128 (
            .O(N__22405),
            .I(\nx.n1598 ));
    Odrv4 I__3127 (
            .O(N__22402),
            .I(\nx.n1598 ));
    CascadeMux I__3126 (
            .O(N__22395),
            .I(N__22382));
    CascadeMux I__3125 (
            .O(N__22394),
            .I(N__22379));
    CascadeMux I__3124 (
            .O(N__22393),
            .I(N__22376));
    CascadeMux I__3123 (
            .O(N__22392),
            .I(N__22373));
    CascadeMux I__3122 (
            .O(N__22391),
            .I(N__22370));
    CascadeMux I__3121 (
            .O(N__22390),
            .I(N__22367));
    CascadeMux I__3120 (
            .O(N__22389),
            .I(N__22364));
    CascadeMux I__3119 (
            .O(N__22388),
            .I(N__22361));
    CascadeMux I__3118 (
            .O(N__22387),
            .I(N__22358));
    CascadeMux I__3117 (
            .O(N__22386),
            .I(N__22355));
    CascadeMux I__3116 (
            .O(N__22385),
            .I(N__22352));
    InMux I__3115 (
            .O(N__22382),
            .I(N__22347));
    InMux I__3114 (
            .O(N__22379),
            .I(N__22347));
    InMux I__3113 (
            .O(N__22376),
            .I(N__22340));
    InMux I__3112 (
            .O(N__22373),
            .I(N__22340));
    InMux I__3111 (
            .O(N__22370),
            .I(N__22340));
    InMux I__3110 (
            .O(N__22367),
            .I(N__22333));
    InMux I__3109 (
            .O(N__22364),
            .I(N__22333));
    InMux I__3108 (
            .O(N__22361),
            .I(N__22333));
    InMux I__3107 (
            .O(N__22358),
            .I(N__22326));
    InMux I__3106 (
            .O(N__22355),
            .I(N__22326));
    InMux I__3105 (
            .O(N__22352),
            .I(N__22326));
    LocalMux I__3104 (
            .O(N__22347),
            .I(\nx.n1631 ));
    LocalMux I__3103 (
            .O(N__22340),
            .I(\nx.n1631 ));
    LocalMux I__3102 (
            .O(N__22333),
            .I(\nx.n1631 ));
    LocalMux I__3101 (
            .O(N__22326),
            .I(\nx.n1631 ));
    InMux I__3100 (
            .O(N__22317),
            .I(\nx.n10805 ));
    CEMux I__3099 (
            .O(N__22314),
            .I(N__22311));
    LocalMux I__3098 (
            .O(N__22311),
            .I(N__22307));
    CEMux I__3097 (
            .O(N__22310),
            .I(N__22304));
    Span4Mux_v I__3096 (
            .O(N__22307),
            .I(N__22297));
    LocalMux I__3095 (
            .O(N__22304),
            .I(N__22297));
    CEMux I__3094 (
            .O(N__22303),
            .I(N__22294));
    CEMux I__3093 (
            .O(N__22302),
            .I(N__22291));
    Span4Mux_v I__3092 (
            .O(N__22297),
            .I(N__22286));
    LocalMux I__3091 (
            .O(N__22294),
            .I(N__22286));
    LocalMux I__3090 (
            .O(N__22291),
            .I(N__22283));
    Span4Mux_h I__3089 (
            .O(N__22286),
            .I(N__22280));
    Span4Mux_s2_h I__3088 (
            .O(N__22283),
            .I(N__22277));
    Odrv4 I__3087 (
            .O(N__22280),
            .I(n7664));
    Odrv4 I__3086 (
            .O(N__22277),
            .I(n7664));
    CascadeMux I__3085 (
            .O(N__22272),
            .I(\nx.n30_adj_777_cascade_ ));
    InMux I__3084 (
            .O(N__22269),
            .I(N__22266));
    LocalMux I__3083 (
            .O(N__22266),
            .I(\nx.n43_adj_783 ));
    InMux I__3082 (
            .O(N__22263),
            .I(bfn_5_25_0_));
    CascadeMux I__3081 (
            .O(N__22260),
            .I(N__22255));
    InMux I__3080 (
            .O(N__22259),
            .I(N__22252));
    InMux I__3079 (
            .O(N__22258),
            .I(N__22249));
    InMux I__3078 (
            .O(N__22255),
            .I(N__22246));
    LocalMux I__3077 (
            .O(N__22252),
            .I(\nx.n1609 ));
    LocalMux I__3076 (
            .O(N__22249),
            .I(\nx.n1609 ));
    LocalMux I__3075 (
            .O(N__22246),
            .I(\nx.n1609 ));
    CascadeMux I__3074 (
            .O(N__22239),
            .I(N__22235));
    CascadeMux I__3073 (
            .O(N__22238),
            .I(N__22232));
    InMux I__3072 (
            .O(N__22235),
            .I(N__22229));
    InMux I__3071 (
            .O(N__22232),
            .I(N__22226));
    LocalMux I__3070 (
            .O(N__22229),
            .I(\nx.n13602 ));
    LocalMux I__3069 (
            .O(N__22226),
            .I(\nx.n13602 ));
    InMux I__3068 (
            .O(N__22221),
            .I(\nx.n10794 ));
    InMux I__3067 (
            .O(N__22218),
            .I(N__22213));
    InMux I__3066 (
            .O(N__22217),
            .I(N__22210));
    InMux I__3065 (
            .O(N__22216),
            .I(N__22207));
    LocalMux I__3064 (
            .O(N__22213),
            .I(\nx.n1608 ));
    LocalMux I__3063 (
            .O(N__22210),
            .I(\nx.n1608 ));
    LocalMux I__3062 (
            .O(N__22207),
            .I(\nx.n1608 ));
    InMux I__3061 (
            .O(N__22200),
            .I(\nx.n10795 ));
    InMux I__3060 (
            .O(N__22197),
            .I(N__22192));
    InMux I__3059 (
            .O(N__22196),
            .I(N__22189));
    InMux I__3058 (
            .O(N__22195),
            .I(N__22186));
    LocalMux I__3057 (
            .O(N__22192),
            .I(\nx.n1607 ));
    LocalMux I__3056 (
            .O(N__22189),
            .I(\nx.n1607 ));
    LocalMux I__3055 (
            .O(N__22186),
            .I(\nx.n1607 ));
    InMux I__3054 (
            .O(N__22179),
            .I(\nx.n10796 ));
    InMux I__3053 (
            .O(N__22176),
            .I(N__22171));
    InMux I__3052 (
            .O(N__22175),
            .I(N__22168));
    InMux I__3051 (
            .O(N__22174),
            .I(N__22165));
    LocalMux I__3050 (
            .O(N__22171),
            .I(\nx.n1606 ));
    LocalMux I__3049 (
            .O(N__22168),
            .I(\nx.n1606 ));
    LocalMux I__3048 (
            .O(N__22165),
            .I(\nx.n1606 ));
    InMux I__3047 (
            .O(N__22158),
            .I(\nx.n10797 ));
    CascadeMux I__3046 (
            .O(N__22155),
            .I(N__22152));
    InMux I__3045 (
            .O(N__22152),
            .I(N__22149));
    LocalMux I__3044 (
            .O(N__22149),
            .I(\nx.n1273 ));
    InMux I__3043 (
            .O(N__22146),
            .I(\nx.n10759 ));
    CascadeMux I__3042 (
            .O(N__22143),
            .I(N__22139));
    InMux I__3041 (
            .O(N__22142),
            .I(N__22136));
    InMux I__3040 (
            .O(N__22139),
            .I(N__22133));
    LocalMux I__3039 (
            .O(N__22136),
            .I(\nx.n1205 ));
    LocalMux I__3038 (
            .O(N__22133),
            .I(\nx.n1205 ));
    InMux I__3037 (
            .O(N__22128),
            .I(N__22125));
    LocalMux I__3036 (
            .O(N__22125),
            .I(\nx.n1272 ));
    InMux I__3035 (
            .O(N__22122),
            .I(\nx.n10760 ));
    CascadeMux I__3034 (
            .O(N__22119),
            .I(N__22115));
    CascadeMux I__3033 (
            .O(N__22118),
            .I(N__22112));
    InMux I__3032 (
            .O(N__22115),
            .I(N__22108));
    InMux I__3031 (
            .O(N__22112),
            .I(N__22105));
    InMux I__3030 (
            .O(N__22111),
            .I(N__22102));
    LocalMux I__3029 (
            .O(N__22108),
            .I(\nx.n1204 ));
    LocalMux I__3028 (
            .O(N__22105),
            .I(\nx.n1204 ));
    LocalMux I__3027 (
            .O(N__22102),
            .I(\nx.n1204 ));
    InMux I__3026 (
            .O(N__22095),
            .I(N__22092));
    LocalMux I__3025 (
            .O(N__22092),
            .I(N__22089));
    Odrv4 I__3024 (
            .O(N__22089),
            .I(\nx.n1271 ));
    InMux I__3023 (
            .O(N__22086),
            .I(\nx.n10761 ));
    InMux I__3022 (
            .O(N__22083),
            .I(\nx.n10762 ));
    CascadeMux I__3021 (
            .O(N__22080),
            .I(N__22077));
    InMux I__3020 (
            .O(N__22077),
            .I(N__22074));
    LocalMux I__3019 (
            .O(N__22074),
            .I(N__22070));
    InMux I__3018 (
            .O(N__22073),
            .I(N__22067));
    Odrv4 I__3017 (
            .O(N__22070),
            .I(\nx.n1202 ));
    LocalMux I__3016 (
            .O(N__22067),
            .I(\nx.n1202 ));
    InMux I__3015 (
            .O(N__22062),
            .I(bfn_5_23_0_));
    CascadeMux I__3014 (
            .O(N__22059),
            .I(N__22055));
    CascadeMux I__3013 (
            .O(N__22058),
            .I(N__22052));
    InMux I__3012 (
            .O(N__22055),
            .I(N__22047));
    InMux I__3011 (
            .O(N__22052),
            .I(N__22047));
    LocalMux I__3010 (
            .O(N__22047),
            .I(\nx.n1301 ));
    InMux I__3009 (
            .O(N__22044),
            .I(N__22041));
    LocalMux I__3008 (
            .O(N__22041),
            .I(N__22037));
    InMux I__3007 (
            .O(N__22040),
            .I(N__22034));
    Span4Mux_h I__3006 (
            .O(N__22037),
            .I(N__22031));
    LocalMux I__3005 (
            .O(N__22034),
            .I(delay_counter_19));
    Odrv4 I__3004 (
            .O(N__22031),
            .I(delay_counter_19));
    InMux I__3003 (
            .O(N__22026),
            .I(N__22023));
    LocalMux I__3002 (
            .O(N__22023),
            .I(N__22019));
    InMux I__3001 (
            .O(N__22022),
            .I(N__22016));
    Span4Mux_h I__3000 (
            .O(N__22019),
            .I(N__22013));
    LocalMux I__2999 (
            .O(N__22016),
            .I(delay_counter_20));
    Odrv4 I__2998 (
            .O(N__22013),
            .I(delay_counter_20));
    InMux I__2997 (
            .O(N__22008),
            .I(N__22005));
    LocalMux I__2996 (
            .O(N__22005),
            .I(N__22002));
    Odrv12 I__2995 (
            .O(N__22002),
            .I(n4));
    CascadeMux I__2994 (
            .O(N__21999),
            .I(N__21995));
    InMux I__2993 (
            .O(N__21998),
            .I(N__21992));
    InMux I__2992 (
            .O(N__21995),
            .I(N__21989));
    LocalMux I__2991 (
            .O(N__21992),
            .I(\nx.n1203 ));
    LocalMux I__2990 (
            .O(N__21989),
            .I(\nx.n1203 ));
    CascadeMux I__2989 (
            .O(N__21984),
            .I(N__21977));
    CascadeMux I__2988 (
            .O(N__21983),
            .I(N__21974));
    CascadeMux I__2987 (
            .O(N__21982),
            .I(N__21969));
    CascadeMux I__2986 (
            .O(N__21981),
            .I(N__21966));
    InMux I__2985 (
            .O(N__21980),
            .I(N__21962));
    InMux I__2984 (
            .O(N__21977),
            .I(N__21955));
    InMux I__2983 (
            .O(N__21974),
            .I(N__21955));
    InMux I__2982 (
            .O(N__21973),
            .I(N__21955));
    InMux I__2981 (
            .O(N__21972),
            .I(N__21950));
    InMux I__2980 (
            .O(N__21969),
            .I(N__21950));
    InMux I__2979 (
            .O(N__21966),
            .I(N__21945));
    InMux I__2978 (
            .O(N__21965),
            .I(N__21945));
    LocalMux I__2977 (
            .O(N__21962),
            .I(\nx.n1235 ));
    LocalMux I__2976 (
            .O(N__21955),
            .I(\nx.n1235 ));
    LocalMux I__2975 (
            .O(N__21950),
            .I(\nx.n1235 ));
    LocalMux I__2974 (
            .O(N__21945),
            .I(\nx.n1235 ));
    InMux I__2973 (
            .O(N__21936),
            .I(N__21933));
    LocalMux I__2972 (
            .O(N__21933),
            .I(\nx.n1270 ));
    CascadeMux I__2971 (
            .O(N__21930),
            .I(N__21926));
    InMux I__2970 (
            .O(N__21929),
            .I(N__21918));
    InMux I__2969 (
            .O(N__21926),
            .I(N__21918));
    InMux I__2968 (
            .O(N__21925),
            .I(N__21918));
    LocalMux I__2967 (
            .O(N__21918),
            .I(\nx.n1302 ));
    CascadeMux I__2966 (
            .O(N__21915),
            .I(\nx.n49_adj_784_cascade_ ));
    InMux I__2965 (
            .O(N__21912),
            .I(N__21909));
    LocalMux I__2964 (
            .O(N__21909),
            .I(N__21906));
    Span4Mux_h I__2963 (
            .O(N__21906),
            .I(N__21903));
    Odrv4 I__2962 (
            .O(N__21903),
            .I(\nx.n54 ));
    CascadeMux I__2961 (
            .O(N__21900),
            .I(N__21896));
    InMux I__2960 (
            .O(N__21899),
            .I(N__21892));
    InMux I__2959 (
            .O(N__21896),
            .I(N__21889));
    InMux I__2958 (
            .O(N__21895),
            .I(N__21886));
    LocalMux I__2957 (
            .O(N__21892),
            .I(\nx.n1106 ));
    LocalMux I__2956 (
            .O(N__21889),
            .I(\nx.n1106 ));
    LocalMux I__2955 (
            .O(N__21886),
            .I(\nx.n1106 ));
    InMux I__2954 (
            .O(N__21879),
            .I(N__21876));
    LocalMux I__2953 (
            .O(N__21876),
            .I(\nx.n1173 ));
    InMux I__2952 (
            .O(N__21873),
            .I(\nx.n10752 ));
    InMux I__2951 (
            .O(N__21870),
            .I(N__21867));
    LocalMux I__2950 (
            .O(N__21867),
            .I(\nx.n1172 ));
    InMux I__2949 (
            .O(N__21864),
            .I(\nx.n10753 ));
    InMux I__2948 (
            .O(N__21861),
            .I(N__21857));
    CascadeMux I__2947 (
            .O(N__21860),
            .I(N__21854));
    LocalMux I__2946 (
            .O(N__21857),
            .I(N__21850));
    InMux I__2945 (
            .O(N__21854),
            .I(N__21847));
    InMux I__2944 (
            .O(N__21853),
            .I(N__21844));
    Odrv4 I__2943 (
            .O(N__21850),
            .I(\nx.n1104 ));
    LocalMux I__2942 (
            .O(N__21847),
            .I(\nx.n1104 ));
    LocalMux I__2941 (
            .O(N__21844),
            .I(\nx.n1104 ));
    InMux I__2940 (
            .O(N__21837),
            .I(N__21834));
    LocalMux I__2939 (
            .O(N__21834),
            .I(\nx.n1171 ));
    InMux I__2938 (
            .O(N__21831),
            .I(\nx.n10754 ));
    CascadeMux I__2937 (
            .O(N__21828),
            .I(N__21822));
    CascadeMux I__2936 (
            .O(N__21827),
            .I(N__21817));
    CascadeMux I__2935 (
            .O(N__21826),
            .I(N__21813));
    CascadeMux I__2934 (
            .O(N__21825),
            .I(N__21810));
    InMux I__2933 (
            .O(N__21822),
            .I(N__21804));
    InMux I__2932 (
            .O(N__21821),
            .I(N__21804));
    InMux I__2931 (
            .O(N__21820),
            .I(N__21801));
    InMux I__2930 (
            .O(N__21817),
            .I(N__21790));
    InMux I__2929 (
            .O(N__21816),
            .I(N__21790));
    InMux I__2928 (
            .O(N__21813),
            .I(N__21790));
    InMux I__2927 (
            .O(N__21810),
            .I(N__21790));
    InMux I__2926 (
            .O(N__21809),
            .I(N__21790));
    LocalMux I__2925 (
            .O(N__21804),
            .I(N__21787));
    LocalMux I__2924 (
            .O(N__21801),
            .I(\nx.n1136 ));
    LocalMux I__2923 (
            .O(N__21790),
            .I(\nx.n1136 ));
    Odrv4 I__2922 (
            .O(N__21787),
            .I(\nx.n1136 ));
    InMux I__2921 (
            .O(N__21780),
            .I(\nx.n10755 ));
    InMux I__2920 (
            .O(N__21777),
            .I(N__21774));
    LocalMux I__2919 (
            .O(N__21774),
            .I(N__21771));
    Span4Mux_h I__2918 (
            .O(N__21771),
            .I(N__21768));
    Odrv4 I__2917 (
            .O(N__21768),
            .I(\nx.n1277 ));
    InMux I__2916 (
            .O(N__21765),
            .I(bfn_5_22_0_));
    CascadeMux I__2915 (
            .O(N__21762),
            .I(N__21757));
    InMux I__2914 (
            .O(N__21761),
            .I(N__21754));
    InMux I__2913 (
            .O(N__21760),
            .I(N__21751));
    InMux I__2912 (
            .O(N__21757),
            .I(N__21748));
    LocalMux I__2911 (
            .O(N__21754),
            .I(\nx.n1209 ));
    LocalMux I__2910 (
            .O(N__21751),
            .I(\nx.n1209 ));
    LocalMux I__2909 (
            .O(N__21748),
            .I(\nx.n1209 ));
    InMux I__2908 (
            .O(N__21741),
            .I(N__21738));
    LocalMux I__2907 (
            .O(N__21738),
            .I(N__21735));
    Span4Mux_h I__2906 (
            .O(N__21735),
            .I(N__21732));
    Odrv4 I__2905 (
            .O(N__21732),
            .I(\nx.n1276 ));
    InMux I__2904 (
            .O(N__21729),
            .I(\nx.n10756 ));
    CascadeMux I__2903 (
            .O(N__21726),
            .I(N__21721));
    InMux I__2902 (
            .O(N__21725),
            .I(N__21716));
    InMux I__2901 (
            .O(N__21724),
            .I(N__21716));
    InMux I__2900 (
            .O(N__21721),
            .I(N__21713));
    LocalMux I__2899 (
            .O(N__21716),
            .I(\nx.n1208 ));
    LocalMux I__2898 (
            .O(N__21713),
            .I(\nx.n1208 ));
    InMux I__2897 (
            .O(N__21708),
            .I(N__21705));
    LocalMux I__2896 (
            .O(N__21705),
            .I(\nx.n1275 ));
    InMux I__2895 (
            .O(N__21702),
            .I(\nx.n10757 ));
    CascadeMux I__2894 (
            .O(N__21699),
            .I(N__21694));
    InMux I__2893 (
            .O(N__21698),
            .I(N__21689));
    InMux I__2892 (
            .O(N__21697),
            .I(N__21689));
    InMux I__2891 (
            .O(N__21694),
            .I(N__21686));
    LocalMux I__2890 (
            .O(N__21689),
            .I(\nx.n1207 ));
    LocalMux I__2889 (
            .O(N__21686),
            .I(\nx.n1207 ));
    InMux I__2888 (
            .O(N__21681),
            .I(N__21678));
    LocalMux I__2887 (
            .O(N__21678),
            .I(\nx.n1274 ));
    InMux I__2886 (
            .O(N__21675),
            .I(\nx.n10758 ));
    CascadeMux I__2885 (
            .O(N__21672),
            .I(N__21667));
    InMux I__2884 (
            .O(N__21671),
            .I(N__21662));
    InMux I__2883 (
            .O(N__21670),
            .I(N__21662));
    InMux I__2882 (
            .O(N__21667),
            .I(N__21659));
    LocalMux I__2881 (
            .O(N__21662),
            .I(\nx.n1206 ));
    LocalMux I__2880 (
            .O(N__21659),
            .I(\nx.n1206 ));
    CascadeMux I__2879 (
            .O(N__21654),
            .I(\nx.n1109_cascade_ ));
    CascadeMux I__2878 (
            .O(N__21651),
            .I(\nx.n9737_cascade_ ));
    CascadeMux I__2877 (
            .O(N__21648),
            .I(\nx.n12_adj_673_cascade_ ));
    InMux I__2876 (
            .O(N__21645),
            .I(N__21642));
    LocalMux I__2875 (
            .O(N__21642),
            .I(N__21639));
    Odrv4 I__2874 (
            .O(N__21639),
            .I(\nx.n1177 ));
    InMux I__2873 (
            .O(N__21636),
            .I(bfn_5_21_0_));
    CascadeMux I__2872 (
            .O(N__21633),
            .I(N__21629));
    InMux I__2871 (
            .O(N__21632),
            .I(N__21626));
    InMux I__2870 (
            .O(N__21629),
            .I(N__21623));
    LocalMux I__2869 (
            .O(N__21626),
            .I(\nx.n1109 ));
    LocalMux I__2868 (
            .O(N__21623),
            .I(\nx.n1109 ));
    CascadeMux I__2867 (
            .O(N__21618),
            .I(N__21615));
    InMux I__2866 (
            .O(N__21615),
            .I(N__21612));
    LocalMux I__2865 (
            .O(N__21612),
            .I(\nx.n1176 ));
    InMux I__2864 (
            .O(N__21609),
            .I(\nx.n10749 ));
    CascadeMux I__2863 (
            .O(N__21606),
            .I(N__21602));
    InMux I__2862 (
            .O(N__21605),
            .I(N__21598));
    InMux I__2861 (
            .O(N__21602),
            .I(N__21595));
    InMux I__2860 (
            .O(N__21601),
            .I(N__21592));
    LocalMux I__2859 (
            .O(N__21598),
            .I(\nx.n1108 ));
    LocalMux I__2858 (
            .O(N__21595),
            .I(\nx.n1108 ));
    LocalMux I__2857 (
            .O(N__21592),
            .I(\nx.n1108 ));
    InMux I__2856 (
            .O(N__21585),
            .I(N__21582));
    LocalMux I__2855 (
            .O(N__21582),
            .I(\nx.n1175 ));
    InMux I__2854 (
            .O(N__21579),
            .I(\nx.n10750 ));
    CascadeMux I__2853 (
            .O(N__21576),
            .I(N__21573));
    InMux I__2852 (
            .O(N__21573),
            .I(N__21570));
    LocalMux I__2851 (
            .O(N__21570),
            .I(\nx.n1174 ));
    InMux I__2850 (
            .O(N__21567),
            .I(\nx.n10751 ));
    InMux I__2849 (
            .O(N__21564),
            .I(N__21561));
    LocalMux I__2848 (
            .O(N__21561),
            .I(N__21557));
    CascadeMux I__2847 (
            .O(N__21560),
            .I(N__21553));
    Span4Mux_h I__2846 (
            .O(N__21557),
            .I(N__21550));
    InMux I__2845 (
            .O(N__21556),
            .I(N__21547));
    InMux I__2844 (
            .O(N__21553),
            .I(N__21544));
    Odrv4 I__2843 (
            .O(N__21550),
            .I(timer_11));
    LocalMux I__2842 (
            .O(N__21547),
            .I(timer_11));
    LocalMux I__2841 (
            .O(N__21544),
            .I(timer_11));
    InMux I__2840 (
            .O(N__21537),
            .I(N__21534));
    LocalMux I__2839 (
            .O(N__21534),
            .I(N__21531));
    Sp12to4 I__2838 (
            .O(N__21531),
            .I(N__21528));
    Span12Mux_v I__2837 (
            .O(N__21528),
            .I(N__21525));
    Odrv12 I__2836 (
            .O(N__21525),
            .I(pin_in_0));
    InMux I__2835 (
            .O(N__21522),
            .I(N__21519));
    LocalMux I__2834 (
            .O(N__21519),
            .I(N__21516));
    Span12Mux_h I__2833 (
            .O(N__21516),
            .I(N__21513));
    Span12Mux_v I__2832 (
            .O(N__21513),
            .I(N__21510));
    Odrv12 I__2831 (
            .O(N__21510),
            .I(pin_in_1));
    InMux I__2830 (
            .O(N__21507),
            .I(N__21504));
    LocalMux I__2829 (
            .O(N__21504),
            .I(N__21501));
    Odrv4 I__2828 (
            .O(N__21501),
            .I(n13378));
    InMux I__2827 (
            .O(N__21498),
            .I(N__21495));
    LocalMux I__2826 (
            .O(N__21495),
            .I(N__21492));
    Span4Mux_h I__2825 (
            .O(N__21492),
            .I(N__21489));
    Span4Mux_v I__2824 (
            .O(N__21489),
            .I(N__21486));
    Sp12to4 I__2823 (
            .O(N__21486),
            .I(N__21483));
    Span12Mux_v I__2822 (
            .O(N__21483),
            .I(N__21480));
    Odrv12 I__2821 (
            .O(N__21480),
            .I(pin_in_4));
    InMux I__2820 (
            .O(N__21477),
            .I(N__21474));
    LocalMux I__2819 (
            .O(N__21474),
            .I(N__21471));
    Span4Mux_v I__2818 (
            .O(N__21471),
            .I(N__21468));
    Span4Mux_v I__2817 (
            .O(N__21468),
            .I(N__21465));
    Span4Mux_v I__2816 (
            .O(N__21465),
            .I(N__21462));
    Span4Mux_h I__2815 (
            .O(N__21462),
            .I(N__21459));
    Odrv4 I__2814 (
            .O(N__21459),
            .I(pin_in_5));
    InMux I__2813 (
            .O(N__21456),
            .I(N__21453));
    LocalMux I__2812 (
            .O(N__21453),
            .I(n13382));
    CascadeMux I__2811 (
            .O(N__21450),
            .I(n13381_cascade_));
    InMux I__2810 (
            .O(N__21447),
            .I(N__21444));
    LocalMux I__2809 (
            .O(N__21444),
            .I(N__21441));
    Odrv4 I__2808 (
            .O(N__21441),
            .I(n13613));
    InMux I__2807 (
            .O(N__21438),
            .I(N__21434));
    InMux I__2806 (
            .O(N__21437),
            .I(N__21431));
    LocalMux I__2805 (
            .O(N__21434),
            .I(neo_pixel_transmitter_t0_11));
    LocalMux I__2804 (
            .O(N__21431),
            .I(neo_pixel_transmitter_t0_11));
    InMux I__2803 (
            .O(N__21426),
            .I(N__21423));
    LocalMux I__2802 (
            .O(N__21423),
            .I(N__21420));
    Span4Mux_h I__2801 (
            .O(N__21420),
            .I(N__21417));
    Odrv4 I__2800 (
            .O(N__21417),
            .I(\nx.n22_adj_749 ));
    InMux I__2799 (
            .O(N__21414),
            .I(N__21410));
    InMux I__2798 (
            .O(N__21413),
            .I(N__21407));
    LocalMux I__2797 (
            .O(N__21410),
            .I(neo_pixel_transmitter_t0_19));
    LocalMux I__2796 (
            .O(N__21407),
            .I(neo_pixel_transmitter_t0_19));
    InMux I__2795 (
            .O(N__21402),
            .I(N__21399));
    LocalMux I__2794 (
            .O(N__21399),
            .I(N__21396));
    Span4Mux_h I__2793 (
            .O(N__21396),
            .I(N__21393));
    Odrv4 I__2792 (
            .O(N__21393),
            .I(\nx.n14 ));
    InMux I__2791 (
            .O(N__21390),
            .I(N__21387));
    LocalMux I__2790 (
            .O(N__21387),
            .I(\nx.n13438 ));
    InMux I__2789 (
            .O(N__21384),
            .I(N__21379));
    InMux I__2788 (
            .O(N__21383),
            .I(N__21376));
    InMux I__2787 (
            .O(N__21382),
            .I(N__21372));
    LocalMux I__2786 (
            .O(N__21379),
            .I(N__21367));
    LocalMux I__2785 (
            .O(N__21376),
            .I(N__21367));
    InMux I__2784 (
            .O(N__21375),
            .I(N__21364));
    LocalMux I__2783 (
            .O(N__21372),
            .I(N__21361));
    Span4Mux_v I__2782 (
            .O(N__21367),
            .I(N__21356));
    LocalMux I__2781 (
            .O(N__21364),
            .I(N__21356));
    Odrv4 I__2780 (
            .O(N__21361),
            .I(\nx.one_wire_N_599_3 ));
    Odrv4 I__2779 (
            .O(N__21356),
            .I(\nx.one_wire_N_599_3 ));
    CascadeMux I__2778 (
            .O(N__21351),
            .I(\nx.n11908_cascade_ ));
    InMux I__2777 (
            .O(N__21348),
            .I(N__21342));
    InMux I__2776 (
            .O(N__21347),
            .I(N__21342));
    LocalMux I__2775 (
            .O(N__21342),
            .I(\nx.n11926 ));
    CascadeMux I__2774 (
            .O(N__21339),
            .I(\nx.n11926_cascade_ ));
    CascadeMux I__2773 (
            .O(N__21336),
            .I(n7671_cascade_));
    InMux I__2772 (
            .O(N__21333),
            .I(N__21328));
    InMux I__2771 (
            .O(N__21332),
            .I(N__21322));
    InMux I__2770 (
            .O(N__21331),
            .I(N__21322));
    LocalMux I__2769 (
            .O(N__21328),
            .I(N__21319));
    InMux I__2768 (
            .O(N__21327),
            .I(N__21316));
    LocalMux I__2767 (
            .O(N__21322),
            .I(N__21313));
    Span4Mux_v I__2766 (
            .O(N__21319),
            .I(N__21310));
    LocalMux I__2765 (
            .O(N__21316),
            .I(N__21307));
    Span4Mux_h I__2764 (
            .O(N__21313),
            .I(N__21304));
    Odrv4 I__2763 (
            .O(N__21310),
            .I(\nx.one_wire_N_599_2 ));
    Odrv4 I__2762 (
            .O(N__21307),
            .I(\nx.one_wire_N_599_2 ));
    Odrv4 I__2761 (
            .O(N__21304),
            .I(\nx.one_wire_N_599_2 ));
    InMux I__2760 (
            .O(N__21297),
            .I(N__21293));
    InMux I__2759 (
            .O(N__21296),
            .I(N__21290));
    LocalMux I__2758 (
            .O(N__21293),
            .I(N__21287));
    LocalMux I__2757 (
            .O(N__21290),
            .I(N__21284));
    Span4Mux_v I__2756 (
            .O(N__21287),
            .I(N__21281));
    Odrv4 I__2755 (
            .O(N__21284),
            .I(\nx.n4_adj_771 ));
    Odrv4 I__2754 (
            .O(N__21281),
            .I(\nx.n4_adj_771 ));
    CascadeMux I__2753 (
            .O(N__21276),
            .I(N__21273));
    InMux I__2752 (
            .O(N__21273),
            .I(N__21270));
    LocalMux I__2751 (
            .O(N__21270),
            .I(N__21265));
    InMux I__2750 (
            .O(N__21269),
            .I(N__21262));
    InMux I__2749 (
            .O(N__21268),
            .I(N__21259));
    Span4Mux_v I__2748 (
            .O(N__21265),
            .I(N__21255));
    LocalMux I__2747 (
            .O(N__21262),
            .I(N__21250));
    LocalMux I__2746 (
            .O(N__21259),
            .I(N__21250));
    InMux I__2745 (
            .O(N__21258),
            .I(N__21247));
    Odrv4 I__2744 (
            .O(N__21255),
            .I(\nx.n9747 ));
    Odrv4 I__2743 (
            .O(N__21250),
            .I(\nx.n9747 ));
    LocalMux I__2742 (
            .O(N__21247),
            .I(\nx.n9747 ));
    InMux I__2741 (
            .O(N__21240),
            .I(N__21237));
    LocalMux I__2740 (
            .O(N__21237),
            .I(\nx.n12381 ));
    InMux I__2739 (
            .O(N__21234),
            .I(N__21231));
    LocalMux I__2738 (
            .O(N__21231),
            .I(N__21228));
    Span4Mux_v I__2737 (
            .O(N__21228),
            .I(N__21225));
    Sp12to4 I__2736 (
            .O(N__21225),
            .I(N__21222));
    Span12Mux_h I__2735 (
            .O(N__21222),
            .I(N__21219));
    Odrv12 I__2734 (
            .O(N__21219),
            .I(pin_in_10));
    CascadeMux I__2733 (
            .O(N__21216),
            .I(N__21213));
    InMux I__2732 (
            .O(N__21213),
            .I(N__21210));
    LocalMux I__2731 (
            .O(N__21210),
            .I(N__21207));
    Span4Mux_v I__2730 (
            .O(N__21207),
            .I(N__21204));
    Span4Mux_h I__2729 (
            .O(N__21204),
            .I(N__21201));
    Span4Mux_v I__2728 (
            .O(N__21201),
            .I(N__21198));
    Span4Mux_v I__2727 (
            .O(N__21198),
            .I(N__21195));
    Odrv4 I__2726 (
            .O(N__21195),
            .I(pin_in_11));
    IoInMux I__2725 (
            .O(N__21192),
            .I(N__21189));
    LocalMux I__2724 (
            .O(N__21189),
            .I(N__21186));
    IoSpan4Mux I__2723 (
            .O(N__21186),
            .I(N__21183));
    Span4Mux_s0_h I__2722 (
            .O(N__21183),
            .I(N__21180));
    Sp12to4 I__2721 (
            .O(N__21180),
            .I(N__21177));
    Span12Mux_v I__2720 (
            .O(N__21177),
            .I(N__21173));
    InMux I__2719 (
            .O(N__21176),
            .I(N__21170));
    Odrv12 I__2718 (
            .O(N__21173),
            .I(pin_oe_6));
    LocalMux I__2717 (
            .O(N__21170),
            .I(pin_oe_6));
    InMux I__2716 (
            .O(N__21165),
            .I(N__21162));
    LocalMux I__2715 (
            .O(N__21162),
            .I(N__21159));
    Span4Mux_h I__2714 (
            .O(N__21159),
            .I(N__21156));
    Sp12to4 I__2713 (
            .O(N__21156),
            .I(N__21153));
    Span12Mux_v I__2712 (
            .O(N__21153),
            .I(N__21150));
    Odrv12 I__2711 (
            .O(N__21150),
            .I(pin_in_9));
    CascadeMux I__2710 (
            .O(N__21147),
            .I(N__21144));
    InMux I__2709 (
            .O(N__21144),
            .I(N__21141));
    LocalMux I__2708 (
            .O(N__21141),
            .I(N__21138));
    Span4Mux_h I__2707 (
            .O(N__21138),
            .I(N__21135));
    Sp12to4 I__2706 (
            .O(N__21135),
            .I(N__21132));
    Span12Mux_v I__2705 (
            .O(N__21132),
            .I(N__21129));
    Odrv12 I__2704 (
            .O(N__21129),
            .I(pin_in_8));
    InMux I__2703 (
            .O(N__21126),
            .I(N__21123));
    LocalMux I__2702 (
            .O(N__21123),
            .I(n13649));
    InMux I__2701 (
            .O(N__21120),
            .I(N__21116));
    CascadeMux I__2700 (
            .O(N__21119),
            .I(N__21113));
    LocalMux I__2699 (
            .O(N__21116),
            .I(N__21110));
    InMux I__2698 (
            .O(N__21113),
            .I(N__21106));
    Span12Mux_v I__2697 (
            .O(N__21110),
            .I(N__21103));
    InMux I__2696 (
            .O(N__21109),
            .I(N__21100));
    LocalMux I__2695 (
            .O(N__21106),
            .I(N__21097));
    Odrv12 I__2694 (
            .O(N__21103),
            .I(timer_30));
    LocalMux I__2693 (
            .O(N__21100),
            .I(timer_30));
    Odrv4 I__2692 (
            .O(N__21097),
            .I(timer_30));
    InMux I__2691 (
            .O(N__21090),
            .I(N__21086));
    InMux I__2690 (
            .O(N__21089),
            .I(N__21083));
    LocalMux I__2689 (
            .O(N__21086),
            .I(neo_pixel_transmitter_t0_30));
    LocalMux I__2688 (
            .O(N__21083),
            .I(neo_pixel_transmitter_t0_30));
    InMux I__2687 (
            .O(N__21078),
            .I(N__21075));
    LocalMux I__2686 (
            .O(N__21075),
            .I(\nx.n11946 ));
    InMux I__2685 (
            .O(N__21072),
            .I(N__21069));
    LocalMux I__2684 (
            .O(N__21069),
            .I(\nx.n13445 ));
    CascadeMux I__2683 (
            .O(N__21066),
            .I(\nx.n11948_cascade_ ));
    InMux I__2682 (
            .O(N__21063),
            .I(N__21060));
    LocalMux I__2681 (
            .O(N__21060),
            .I(N__21057));
    Span4Mux_v I__2680 (
            .O(N__21057),
            .I(N__21054));
    Span4Mux_h I__2679 (
            .O(N__21054),
            .I(N__21051));
    Odrv4 I__2678 (
            .O(N__21051),
            .I(pin_in_2));
    InMux I__2677 (
            .O(N__21048),
            .I(N__21045));
    LocalMux I__2676 (
            .O(N__21045),
            .I(N__21042));
    Span4Mux_v I__2675 (
            .O(N__21042),
            .I(N__21039));
    Span4Mux_h I__2674 (
            .O(N__21039),
            .I(N__21036));
    Odrv4 I__2673 (
            .O(N__21036),
            .I(pin_in_3));
    CascadeMux I__2672 (
            .O(N__21033),
            .I(n13379_cascade_));
    InMux I__2671 (
            .O(N__21030),
            .I(N__21025));
    InMux I__2670 (
            .O(N__21029),
            .I(N__21022));
    InMux I__2669 (
            .O(N__21028),
            .I(N__21019));
    LocalMux I__2668 (
            .O(N__21025),
            .I(\nx.n1504 ));
    LocalMux I__2667 (
            .O(N__21022),
            .I(\nx.n1504 ));
    LocalMux I__2666 (
            .O(N__21019),
            .I(\nx.n1504 ));
    InMux I__2665 (
            .O(N__21012),
            .I(\nx.n10788 ));
    InMux I__2664 (
            .O(N__21009),
            .I(N__21004));
    InMux I__2663 (
            .O(N__21008),
            .I(N__21001));
    InMux I__2662 (
            .O(N__21007),
            .I(N__20998));
    LocalMux I__2661 (
            .O(N__21004),
            .I(\nx.n1503 ));
    LocalMux I__2660 (
            .O(N__21001),
            .I(\nx.n1503 ));
    LocalMux I__2659 (
            .O(N__20998),
            .I(\nx.n1503 ));
    InMux I__2658 (
            .O(N__20991),
            .I(\nx.n10789 ));
    InMux I__2657 (
            .O(N__20988),
            .I(N__20984));
    InMux I__2656 (
            .O(N__20987),
            .I(N__20981));
    LocalMux I__2655 (
            .O(N__20984),
            .I(N__20976));
    LocalMux I__2654 (
            .O(N__20981),
            .I(N__20976));
    Odrv4 I__2653 (
            .O(N__20976),
            .I(\nx.n1502 ));
    InMux I__2652 (
            .O(N__20973),
            .I(bfn_4_27_0_));
    InMux I__2651 (
            .O(N__20970),
            .I(N__20966));
    InMux I__2650 (
            .O(N__20969),
            .I(N__20963));
    LocalMux I__2649 (
            .O(N__20966),
            .I(N__20958));
    LocalMux I__2648 (
            .O(N__20963),
            .I(N__20958));
    Span4Mux_h I__2647 (
            .O(N__20958),
            .I(N__20954));
    InMux I__2646 (
            .O(N__20957),
            .I(N__20951));
    Odrv4 I__2645 (
            .O(N__20954),
            .I(\nx.n1501 ));
    LocalMux I__2644 (
            .O(N__20951),
            .I(\nx.n1501 ));
    InMux I__2643 (
            .O(N__20946),
            .I(\nx.n10791 ));
    InMux I__2642 (
            .O(N__20943),
            .I(N__20938));
    InMux I__2641 (
            .O(N__20942),
            .I(N__20935));
    InMux I__2640 (
            .O(N__20941),
            .I(N__20932));
    LocalMux I__2639 (
            .O(N__20938),
            .I(\nx.n1500 ));
    LocalMux I__2638 (
            .O(N__20935),
            .I(\nx.n1500 ));
    LocalMux I__2637 (
            .O(N__20932),
            .I(\nx.n1500 ));
    InMux I__2636 (
            .O(N__20925),
            .I(\nx.n10792 ));
    InMux I__2635 (
            .O(N__20922),
            .I(N__20918));
    InMux I__2634 (
            .O(N__20921),
            .I(N__20915));
    LocalMux I__2633 (
            .O(N__20918),
            .I(N__20910));
    LocalMux I__2632 (
            .O(N__20915),
            .I(N__20910));
    Span4Mux_h I__2631 (
            .O(N__20910),
            .I(N__20906));
    InMux I__2630 (
            .O(N__20909),
            .I(N__20903));
    Odrv4 I__2629 (
            .O(N__20906),
            .I(\nx.n1499 ));
    LocalMux I__2628 (
            .O(N__20903),
            .I(\nx.n1499 ));
    CascadeMux I__2627 (
            .O(N__20898),
            .I(N__20886));
    CascadeMux I__2626 (
            .O(N__20897),
            .I(N__20883));
    CascadeMux I__2625 (
            .O(N__20896),
            .I(N__20880));
    CascadeMux I__2624 (
            .O(N__20895),
            .I(N__20877));
    CascadeMux I__2623 (
            .O(N__20894),
            .I(N__20874));
    CascadeMux I__2622 (
            .O(N__20893),
            .I(N__20871));
    CascadeMux I__2621 (
            .O(N__20892),
            .I(N__20868));
    CascadeMux I__2620 (
            .O(N__20891),
            .I(N__20865));
    CascadeMux I__2619 (
            .O(N__20890),
            .I(N__20862));
    CascadeMux I__2618 (
            .O(N__20889),
            .I(N__20859));
    InMux I__2617 (
            .O(N__20886),
            .I(N__20854));
    InMux I__2616 (
            .O(N__20883),
            .I(N__20854));
    InMux I__2615 (
            .O(N__20880),
            .I(N__20849));
    InMux I__2614 (
            .O(N__20877),
            .I(N__20849));
    InMux I__2613 (
            .O(N__20874),
            .I(N__20842));
    InMux I__2612 (
            .O(N__20871),
            .I(N__20842));
    InMux I__2611 (
            .O(N__20868),
            .I(N__20842));
    InMux I__2610 (
            .O(N__20865),
            .I(N__20835));
    InMux I__2609 (
            .O(N__20862),
            .I(N__20835));
    InMux I__2608 (
            .O(N__20859),
            .I(N__20835));
    LocalMux I__2607 (
            .O(N__20854),
            .I(\nx.n1532 ));
    LocalMux I__2606 (
            .O(N__20849),
            .I(\nx.n1532 ));
    LocalMux I__2605 (
            .O(N__20842),
            .I(\nx.n1532 ));
    LocalMux I__2604 (
            .O(N__20835),
            .I(\nx.n1532 ));
    InMux I__2603 (
            .O(N__20826),
            .I(\nx.n10793 ));
    InMux I__2602 (
            .O(N__20823),
            .I(N__20820));
    LocalMux I__2601 (
            .O(N__20820),
            .I(\nx.n45_adj_781 ));
    InMux I__2600 (
            .O(N__20817),
            .I(N__20814));
    LocalMux I__2599 (
            .O(N__20814),
            .I(N__20811));
    Odrv4 I__2598 (
            .O(N__20811),
            .I(\nx.n19 ));
    InMux I__2597 (
            .O(N__20808),
            .I(N__20805));
    LocalMux I__2596 (
            .O(N__20805),
            .I(N__20802));
    Odrv4 I__2595 (
            .O(N__20802),
            .I(\nx.n47_adj_780 ));
    InMux I__2594 (
            .O(N__20799),
            .I(N__20796));
    LocalMux I__2593 (
            .O(N__20796),
            .I(\nx.n18 ));
    InMux I__2592 (
            .O(N__20793),
            .I(N__20789));
    InMux I__2591 (
            .O(N__20792),
            .I(N__20786));
    LocalMux I__2590 (
            .O(N__20789),
            .I(N__20783));
    LocalMux I__2589 (
            .O(N__20786),
            .I(delay_counter_28));
    Odrv4 I__2588 (
            .O(N__20783),
            .I(delay_counter_28));
    InMux I__2587 (
            .O(N__20778),
            .I(N__20774));
    InMux I__2586 (
            .O(N__20777),
            .I(N__20771));
    LocalMux I__2585 (
            .O(N__20774),
            .I(N__20768));
    LocalMux I__2584 (
            .O(N__20771),
            .I(delay_counter_24));
    Odrv4 I__2583 (
            .O(N__20768),
            .I(delay_counter_24));
    CascadeMux I__2582 (
            .O(N__20763),
            .I(N__20760));
    InMux I__2581 (
            .O(N__20760),
            .I(N__20757));
    LocalMux I__2580 (
            .O(N__20757),
            .I(N__20753));
    InMux I__2579 (
            .O(N__20756),
            .I(N__20750));
    Span4Mux_h I__2578 (
            .O(N__20753),
            .I(N__20747));
    LocalMux I__2577 (
            .O(N__20750),
            .I(delay_counter_22));
    Odrv4 I__2576 (
            .O(N__20747),
            .I(delay_counter_22));
    InMux I__2575 (
            .O(N__20742),
            .I(N__20738));
    InMux I__2574 (
            .O(N__20741),
            .I(N__20735));
    LocalMux I__2573 (
            .O(N__20738),
            .I(N__20732));
    LocalMux I__2572 (
            .O(N__20735),
            .I(delay_counter_26));
    Odrv4 I__2571 (
            .O(N__20732),
            .I(delay_counter_26));
    InMux I__2570 (
            .O(N__20727),
            .I(bfn_4_26_0_));
    InMux I__2569 (
            .O(N__20724),
            .I(N__20720));
    InMux I__2568 (
            .O(N__20723),
            .I(N__20717));
    LocalMux I__2567 (
            .O(N__20720),
            .I(\nx.n1509 ));
    LocalMux I__2566 (
            .O(N__20717),
            .I(\nx.n1509 ));
    CascadeMux I__2565 (
            .O(N__20712),
            .I(N__20708));
    CascadeMux I__2564 (
            .O(N__20711),
            .I(N__20705));
    InMux I__2563 (
            .O(N__20708),
            .I(N__20702));
    InMux I__2562 (
            .O(N__20705),
            .I(N__20699));
    LocalMux I__2561 (
            .O(N__20702),
            .I(\nx.n13604 ));
    LocalMux I__2560 (
            .O(N__20699),
            .I(\nx.n13604 ));
    InMux I__2559 (
            .O(N__20694),
            .I(\nx.n10783 ));
    InMux I__2558 (
            .O(N__20691),
            .I(N__20686));
    InMux I__2557 (
            .O(N__20690),
            .I(N__20683));
    InMux I__2556 (
            .O(N__20689),
            .I(N__20680));
    LocalMux I__2555 (
            .O(N__20686),
            .I(\nx.n1508 ));
    LocalMux I__2554 (
            .O(N__20683),
            .I(\nx.n1508 ));
    LocalMux I__2553 (
            .O(N__20680),
            .I(\nx.n1508 ));
    InMux I__2552 (
            .O(N__20673),
            .I(\nx.n10784 ));
    InMux I__2551 (
            .O(N__20670),
            .I(N__20666));
    InMux I__2550 (
            .O(N__20669),
            .I(N__20663));
    LocalMux I__2549 (
            .O(N__20666),
            .I(\nx.n1507 ));
    LocalMux I__2548 (
            .O(N__20663),
            .I(\nx.n1507 ));
    InMux I__2547 (
            .O(N__20658),
            .I(\nx.n10785 ));
    InMux I__2546 (
            .O(N__20655),
            .I(N__20650));
    InMux I__2545 (
            .O(N__20654),
            .I(N__20647));
    InMux I__2544 (
            .O(N__20653),
            .I(N__20644));
    LocalMux I__2543 (
            .O(N__20650),
            .I(\nx.n1506 ));
    LocalMux I__2542 (
            .O(N__20647),
            .I(\nx.n1506 ));
    LocalMux I__2541 (
            .O(N__20644),
            .I(\nx.n1506 ));
    InMux I__2540 (
            .O(N__20637),
            .I(\nx.n10786 ));
    InMux I__2539 (
            .O(N__20634),
            .I(N__20629));
    InMux I__2538 (
            .O(N__20633),
            .I(N__20626));
    InMux I__2537 (
            .O(N__20632),
            .I(N__20623));
    LocalMux I__2536 (
            .O(N__20629),
            .I(\nx.n1505 ));
    LocalMux I__2535 (
            .O(N__20626),
            .I(\nx.n1505 ));
    LocalMux I__2534 (
            .O(N__20623),
            .I(\nx.n1505 ));
    InMux I__2533 (
            .O(N__20616),
            .I(\nx.n10787 ));
    InMux I__2532 (
            .O(N__20613),
            .I(N__20609));
    InMux I__2531 (
            .O(N__20612),
            .I(N__20606));
    LocalMux I__2530 (
            .O(N__20609),
            .I(N__20603));
    LocalMux I__2529 (
            .O(N__20606),
            .I(delay_counter_18));
    Odrv4 I__2528 (
            .O(N__20603),
            .I(delay_counter_18));
    InMux I__2527 (
            .O(N__20598),
            .I(N__20594));
    InMux I__2526 (
            .O(N__20597),
            .I(N__20591));
    LocalMux I__2525 (
            .O(N__20594),
            .I(N__20588));
    LocalMux I__2524 (
            .O(N__20591),
            .I(delay_counter_16));
    Odrv4 I__2523 (
            .O(N__20588),
            .I(delay_counter_16));
    InMux I__2522 (
            .O(N__20583),
            .I(N__20580));
    LocalMux I__2521 (
            .O(N__20580),
            .I(N__20577));
    Odrv4 I__2520 (
            .O(N__20577),
            .I(n6_adj_843));
    CascadeMux I__2519 (
            .O(N__20574),
            .I(N__20569));
    InMux I__2518 (
            .O(N__20573),
            .I(N__20566));
    InMux I__2517 (
            .O(N__20572),
            .I(N__20563));
    InMux I__2516 (
            .O(N__20569),
            .I(N__20560));
    LocalMux I__2515 (
            .O(N__20566),
            .I(N__20555));
    LocalMux I__2514 (
            .O(N__20563),
            .I(N__20555));
    LocalMux I__2513 (
            .O(N__20560),
            .I(\nx.n1304 ));
    Odrv4 I__2512 (
            .O(N__20555),
            .I(\nx.n1304 ));
    CascadeMux I__2511 (
            .O(N__20550),
            .I(N__20546));
    CascadeMux I__2510 (
            .O(N__20549),
            .I(N__20542));
    InMux I__2509 (
            .O(N__20546),
            .I(N__20539));
    InMux I__2508 (
            .O(N__20545),
            .I(N__20536));
    InMux I__2507 (
            .O(N__20542),
            .I(N__20533));
    LocalMux I__2506 (
            .O(N__20539),
            .I(N__20528));
    LocalMux I__2505 (
            .O(N__20536),
            .I(N__20528));
    LocalMux I__2504 (
            .O(N__20533),
            .I(\nx.n1305 ));
    Odrv4 I__2503 (
            .O(N__20528),
            .I(\nx.n1305 ));
    CascadeMux I__2502 (
            .O(N__20523),
            .I(\nx.n10_adj_668_cascade_ ));
    CascadeMux I__2501 (
            .O(N__20520),
            .I(N__20515));
    InMux I__2500 (
            .O(N__20519),
            .I(N__20512));
    InMux I__2499 (
            .O(N__20518),
            .I(N__20509));
    InMux I__2498 (
            .O(N__20515),
            .I(N__20506));
    LocalMux I__2497 (
            .O(N__20512),
            .I(N__20501));
    LocalMux I__2496 (
            .O(N__20509),
            .I(N__20501));
    LocalMux I__2495 (
            .O(N__20506),
            .I(\nx.n1307 ));
    Odrv4 I__2494 (
            .O(N__20501),
            .I(\nx.n1307 ));
    InMux I__2493 (
            .O(N__20496),
            .I(N__20493));
    LocalMux I__2492 (
            .O(N__20493),
            .I(\nx.n16 ));
    CascadeMux I__2491 (
            .O(N__20490),
            .I(N__20487));
    InMux I__2490 (
            .O(N__20487),
            .I(N__20484));
    LocalMux I__2489 (
            .O(N__20484),
            .I(\nx.n1369 ));
    CascadeMux I__2488 (
            .O(N__20481),
            .I(N__20477));
    CascadeMux I__2487 (
            .O(N__20480),
            .I(N__20471));
    InMux I__2486 (
            .O(N__20477),
            .I(N__20462));
    InMux I__2485 (
            .O(N__20476),
            .I(N__20462));
    InMux I__2484 (
            .O(N__20475),
            .I(N__20453));
    InMux I__2483 (
            .O(N__20474),
            .I(N__20453));
    InMux I__2482 (
            .O(N__20471),
            .I(N__20453));
    InMux I__2481 (
            .O(N__20470),
            .I(N__20453));
    InMux I__2480 (
            .O(N__20469),
            .I(N__20448));
    InMux I__2479 (
            .O(N__20468),
            .I(N__20448));
    InMux I__2478 (
            .O(N__20467),
            .I(N__20445));
    LocalMux I__2477 (
            .O(N__20462),
            .I(\nx.n1334 ));
    LocalMux I__2476 (
            .O(N__20453),
            .I(\nx.n1334 ));
    LocalMux I__2475 (
            .O(N__20448),
            .I(\nx.n1334 ));
    LocalMux I__2474 (
            .O(N__20445),
            .I(\nx.n1334 ));
    CascadeMux I__2473 (
            .O(N__20436),
            .I(N__20433));
    InMux I__2472 (
            .O(N__20433),
            .I(N__20429));
    InMux I__2471 (
            .O(N__20432),
            .I(N__20426));
    LocalMux I__2470 (
            .O(N__20429),
            .I(N__20423));
    LocalMux I__2469 (
            .O(N__20426),
            .I(N__20419));
    Span4Mux_s3_h I__2468 (
            .O(N__20423),
            .I(N__20416));
    InMux I__2467 (
            .O(N__20422),
            .I(N__20413));
    Odrv4 I__2466 (
            .O(N__20419),
            .I(\nx.n1401 ));
    Odrv4 I__2465 (
            .O(N__20416),
            .I(\nx.n1401 ));
    LocalMux I__2464 (
            .O(N__20413),
            .I(\nx.n1401 ));
    SRMux I__2463 (
            .O(N__20406),
            .I(N__20403));
    LocalMux I__2462 (
            .O(N__20403),
            .I(N__20400));
    Sp12to4 I__2461 (
            .O(N__20400),
            .I(N__20397));
    Odrv12 I__2460 (
            .O(N__20397),
            .I(n22_adj_795));
    CascadeMux I__2459 (
            .O(N__20394),
            .I(\nx.n1631_cascade_ ));
    CascadeMux I__2458 (
            .O(N__20391),
            .I(\nx.n15_adj_676_cascade_ ));
    InMux I__2457 (
            .O(N__20388),
            .I(N__20385));
    LocalMux I__2456 (
            .O(N__20385),
            .I(\nx.n22 ));
    CascadeMux I__2455 (
            .O(N__20382),
            .I(N__20378));
    InMux I__2454 (
            .O(N__20381),
            .I(N__20375));
    InMux I__2453 (
            .O(N__20378),
            .I(N__20372));
    LocalMux I__2452 (
            .O(N__20375),
            .I(\nx.n1308 ));
    LocalMux I__2451 (
            .O(N__20372),
            .I(\nx.n1308 ));
    InMux I__2450 (
            .O(N__20367),
            .I(N__20364));
    LocalMux I__2449 (
            .O(N__20364),
            .I(N__20361));
    Span4Mux_s3_h I__2448 (
            .O(N__20361),
            .I(N__20358));
    Odrv4 I__2447 (
            .O(N__20358),
            .I(\nx.n1375 ));
    InMux I__2446 (
            .O(N__20355),
            .I(\nx.n10765 ));
    InMux I__2445 (
            .O(N__20352),
            .I(N__20349));
    LocalMux I__2444 (
            .O(N__20349),
            .I(\nx.n1374 ));
    InMux I__2443 (
            .O(N__20346),
            .I(\nx.n10766 ));
    CascadeMux I__2442 (
            .O(N__20343),
            .I(N__20338));
    InMux I__2441 (
            .O(N__20342),
            .I(N__20333));
    InMux I__2440 (
            .O(N__20341),
            .I(N__20333));
    InMux I__2439 (
            .O(N__20338),
            .I(N__20330));
    LocalMux I__2438 (
            .O(N__20333),
            .I(\nx.n1306 ));
    LocalMux I__2437 (
            .O(N__20330),
            .I(\nx.n1306 ));
    CascadeMux I__2436 (
            .O(N__20325),
            .I(N__20322));
    InMux I__2435 (
            .O(N__20322),
            .I(N__20319));
    LocalMux I__2434 (
            .O(N__20319),
            .I(\nx.n1373 ));
    InMux I__2433 (
            .O(N__20316),
            .I(\nx.n10767 ));
    InMux I__2432 (
            .O(N__20313),
            .I(N__20310));
    LocalMux I__2431 (
            .O(N__20310),
            .I(\nx.n1372 ));
    InMux I__2430 (
            .O(N__20307),
            .I(\nx.n10768 ));
    CascadeMux I__2429 (
            .O(N__20304),
            .I(N__20301));
    InMux I__2428 (
            .O(N__20301),
            .I(N__20298));
    LocalMux I__2427 (
            .O(N__20298),
            .I(\nx.n1371 ));
    InMux I__2426 (
            .O(N__20295),
            .I(\nx.n10769 ));
    CascadeMux I__2425 (
            .O(N__20292),
            .I(N__20287));
    InMux I__2424 (
            .O(N__20291),
            .I(N__20282));
    InMux I__2423 (
            .O(N__20290),
            .I(N__20282));
    InMux I__2422 (
            .O(N__20287),
            .I(N__20279));
    LocalMux I__2421 (
            .O(N__20282),
            .I(\nx.n1303 ));
    LocalMux I__2420 (
            .O(N__20279),
            .I(\nx.n1303 ));
    InMux I__2419 (
            .O(N__20274),
            .I(N__20271));
    LocalMux I__2418 (
            .O(N__20271),
            .I(\nx.n1370 ));
    InMux I__2417 (
            .O(N__20268),
            .I(\nx.n10770 ));
    InMux I__2416 (
            .O(N__20265),
            .I(bfn_4_24_0_));
    InMux I__2415 (
            .O(N__20262),
            .I(\nx.n10772 ));
    InMux I__2414 (
            .O(N__20259),
            .I(N__20256));
    LocalMux I__2413 (
            .O(N__20256),
            .I(N__20253));
    Span4Mux_s3_h I__2412 (
            .O(N__20253),
            .I(N__20249));
    InMux I__2411 (
            .O(N__20252),
            .I(N__20246));
    Odrv4 I__2410 (
            .O(N__20249),
            .I(\nx.n1400 ));
    LocalMux I__2409 (
            .O(N__20246),
            .I(\nx.n1400 ));
    CascadeMux I__2408 (
            .O(N__20241),
            .I(\nx.n1235_cascade_ ));
    CascadeMux I__2407 (
            .O(N__20238),
            .I(\nx.n1203_cascade_ ));
    CascadeMux I__2406 (
            .O(N__20235),
            .I(N__20232));
    InMux I__2405 (
            .O(N__20232),
            .I(N__20229));
    LocalMux I__2404 (
            .O(N__20229),
            .I(\nx.n13_adj_675 ));
    InMux I__2403 (
            .O(N__20226),
            .I(N__20223));
    LocalMux I__2402 (
            .O(N__20223),
            .I(N__20220));
    Span4Mux_s3_h I__2401 (
            .O(N__20220),
            .I(N__20217));
    Odrv4 I__2400 (
            .O(N__20217),
            .I(\nx.n1377 ));
    InMux I__2399 (
            .O(N__20214),
            .I(bfn_4_23_0_));
    CascadeMux I__2398 (
            .O(N__20211),
            .I(N__20207));
    InMux I__2397 (
            .O(N__20210),
            .I(N__20204));
    InMux I__2396 (
            .O(N__20207),
            .I(N__20201));
    LocalMux I__2395 (
            .O(N__20204),
            .I(\nx.n1309 ));
    LocalMux I__2394 (
            .O(N__20201),
            .I(\nx.n1309 ));
    CascadeMux I__2393 (
            .O(N__20196),
            .I(N__20193));
    InMux I__2392 (
            .O(N__20193),
            .I(N__20190));
    LocalMux I__2391 (
            .O(N__20190),
            .I(\nx.n1376 ));
    InMux I__2390 (
            .O(N__20187),
            .I(\nx.n10764 ));
    CascadeMux I__2389 (
            .O(N__20184),
            .I(N__20181));
    InMux I__2388 (
            .O(N__20181),
            .I(N__20178));
    LocalMux I__2387 (
            .O(N__20178),
            .I(N__20173));
    InMux I__2386 (
            .O(N__20177),
            .I(N__20170));
    InMux I__2385 (
            .O(N__20176),
            .I(N__20167));
    Span4Mux_v I__2384 (
            .O(N__20173),
            .I(N__20164));
    LocalMux I__2383 (
            .O(N__20170),
            .I(timer_29));
    LocalMux I__2382 (
            .O(N__20167),
            .I(timer_29));
    Odrv4 I__2381 (
            .O(N__20164),
            .I(timer_29));
    InMux I__2380 (
            .O(N__20157),
            .I(N__20154));
    LocalMux I__2379 (
            .O(N__20154),
            .I(N__20150));
    InMux I__2378 (
            .O(N__20153),
            .I(N__20147));
    Span4Mux_h I__2377 (
            .O(N__20150),
            .I(N__20144));
    LocalMux I__2376 (
            .O(N__20147),
            .I(neo_pixel_transmitter_t0_29));
    Odrv4 I__2375 (
            .O(N__20144),
            .I(neo_pixel_transmitter_t0_29));
    InMux I__2374 (
            .O(N__20139),
            .I(N__20135));
    InMux I__2373 (
            .O(N__20138),
            .I(N__20132));
    LocalMux I__2372 (
            .O(N__20135),
            .I(neo_pixel_transmitter_t0_25));
    LocalMux I__2371 (
            .O(N__20132),
            .I(neo_pixel_transmitter_t0_25));
    CascadeMux I__2370 (
            .O(N__20127),
            .I(N__20124));
    InMux I__2369 (
            .O(N__20124),
            .I(N__20121));
    LocalMux I__2368 (
            .O(N__20121),
            .I(N__20118));
    Span4Mux_s3_h I__2367 (
            .O(N__20118),
            .I(N__20115));
    Odrv4 I__2366 (
            .O(N__20115),
            .I(\nx.n8 ));
    CascadeMux I__2365 (
            .O(N__20112),
            .I(\nx.n1205_cascade_ ));
    InMux I__2364 (
            .O(N__20109),
            .I(N__20106));
    LocalMux I__2363 (
            .O(N__20106),
            .I(\nx.n11_adj_674 ));
    CascadeMux I__2362 (
            .O(N__20103),
            .I(\nx.n6_adj_786_cascade_ ));
    InMux I__2361 (
            .O(N__20100),
            .I(N__20096));
    InMux I__2360 (
            .O(N__20099),
            .I(N__20093));
    LocalMux I__2359 (
            .O(N__20096),
            .I(N__20090));
    LocalMux I__2358 (
            .O(N__20093),
            .I(N__20087));
    Span4Mux_h I__2357 (
            .O(N__20090),
            .I(N__20084));
    Odrv4 I__2356 (
            .O(N__20087),
            .I(\nx.one_wire_N_599_5 ));
    Odrv4 I__2355 (
            .O(N__20084),
            .I(\nx.one_wire_N_599_5 ));
    CEMux I__2354 (
            .O(N__20079),
            .I(N__20076));
    LocalMux I__2353 (
            .O(N__20076),
            .I(N__20073));
    Span4Mux_v I__2352 (
            .O(N__20073),
            .I(N__20070));
    Odrv4 I__2351 (
            .O(N__20070),
            .I(\nx.n13659 ));
    InMux I__2350 (
            .O(N__20067),
            .I(N__20064));
    LocalMux I__2349 (
            .O(N__20064),
            .I(N__20060));
    InMux I__2348 (
            .O(N__20063),
            .I(N__20057));
    Span4Mux_v I__2347 (
            .O(N__20060),
            .I(N__20052));
    LocalMux I__2346 (
            .O(N__20057),
            .I(N__20052));
    Odrv4 I__2345 (
            .O(N__20052),
            .I(\nx.one_wire_N_599_7 ));
    InMux I__2344 (
            .O(N__20049),
            .I(N__20040));
    InMux I__2343 (
            .O(N__20048),
            .I(N__20040));
    InMux I__2342 (
            .O(N__20047),
            .I(N__20040));
    LocalMux I__2341 (
            .O(N__20040),
            .I(N__20037));
    Span4Mux_v I__2340 (
            .O(N__20037),
            .I(N__20034));
    Odrv4 I__2339 (
            .O(N__20034),
            .I(\nx.one_wire_N_599_8 ));
    CascadeMux I__2338 (
            .O(N__20031),
            .I(N__20027));
    InMux I__2337 (
            .O(N__20030),
            .I(N__20022));
    InMux I__2336 (
            .O(N__20027),
            .I(N__20022));
    LocalMux I__2335 (
            .O(N__20022),
            .I(N__20019));
    Odrv4 I__2334 (
            .O(N__20019),
            .I(\nx.one_wire_N_599_6 ));
    InMux I__2333 (
            .O(N__20016),
            .I(N__20013));
    LocalMux I__2332 (
            .O(N__20013),
            .I(\nx.n13211 ));
    CascadeMux I__2331 (
            .O(N__20010),
            .I(N__20006));
    InMux I__2330 (
            .O(N__20009),
            .I(N__19998));
    InMux I__2329 (
            .O(N__20006),
            .I(N__19998));
    InMux I__2328 (
            .O(N__20005),
            .I(N__19998));
    LocalMux I__2327 (
            .O(N__19998),
            .I(N__19995));
    Span4Mux_h I__2326 (
            .O(N__19995),
            .I(N__19992));
    Odrv4 I__2325 (
            .O(N__19992),
            .I(\nx.one_wire_N_599_10 ));
    InMux I__2324 (
            .O(N__19989),
            .I(N__19984));
    InMux I__2323 (
            .O(N__19988),
            .I(N__19979));
    InMux I__2322 (
            .O(N__19987),
            .I(N__19979));
    LocalMux I__2321 (
            .O(N__19984),
            .I(N__19976));
    LocalMux I__2320 (
            .O(N__19979),
            .I(N__19973));
    Span4Mux_v I__2319 (
            .O(N__19976),
            .I(N__19968));
    Span4Mux_v I__2318 (
            .O(N__19973),
            .I(N__19968));
    Odrv4 I__2317 (
            .O(N__19968),
            .I(\nx.one_wire_N_599_9 ));
    CascadeMux I__2316 (
            .O(N__19965),
            .I(\nx.n13217_cascade_ ));
    InMux I__2315 (
            .O(N__19962),
            .I(N__19953));
    InMux I__2314 (
            .O(N__19961),
            .I(N__19953));
    InMux I__2313 (
            .O(N__19960),
            .I(N__19953));
    LocalMux I__2312 (
            .O(N__19953),
            .I(N__19950));
    Span4Mux_h I__2311 (
            .O(N__19950),
            .I(N__19947));
    Odrv4 I__2310 (
            .O(N__19947),
            .I(\nx.n7608 ));
    InMux I__2309 (
            .O(N__19944),
            .I(N__19941));
    LocalMux I__2308 (
            .O(N__19941),
            .I(N__19938));
    Span4Mux_s3_h I__2307 (
            .O(N__19938),
            .I(N__19935));
    Odrv4 I__2306 (
            .O(N__19935),
            .I(\nx.n20_adj_726 ));
    CascadeMux I__2305 (
            .O(N__19932),
            .I(N__19929));
    InMux I__2304 (
            .O(N__19929),
            .I(N__19924));
    InMux I__2303 (
            .O(N__19928),
            .I(N__19921));
    InMux I__2302 (
            .O(N__19927),
            .I(N__19918));
    LocalMux I__2301 (
            .O(N__19924),
            .I(N__19915));
    LocalMux I__2300 (
            .O(N__19921),
            .I(timer_13));
    LocalMux I__2299 (
            .O(N__19918),
            .I(timer_13));
    Odrv4 I__2298 (
            .O(N__19915),
            .I(timer_13));
    InMux I__2297 (
            .O(N__19908),
            .I(N__19902));
    InMux I__2296 (
            .O(N__19907),
            .I(N__19902));
    LocalMux I__2295 (
            .O(N__19902),
            .I(neo_pixel_transmitter_t0_13));
    InMux I__2294 (
            .O(N__19899),
            .I(N__19894));
    InMux I__2293 (
            .O(N__19898),
            .I(N__19891));
    InMux I__2292 (
            .O(N__19897),
            .I(N__19888));
    LocalMux I__2291 (
            .O(N__19894),
            .I(timer_25));
    LocalMux I__2290 (
            .O(N__19891),
            .I(timer_25));
    LocalMux I__2289 (
            .O(N__19888),
            .I(timer_25));
    CascadeMux I__2288 (
            .O(N__19881),
            .I(N__19876));
    InMux I__2287 (
            .O(N__19880),
            .I(N__19873));
    InMux I__2286 (
            .O(N__19879),
            .I(N__19870));
    InMux I__2285 (
            .O(N__19876),
            .I(N__19867));
    LocalMux I__2284 (
            .O(N__19873),
            .I(timer_19));
    LocalMux I__2283 (
            .O(N__19870),
            .I(timer_19));
    LocalMux I__2282 (
            .O(N__19867),
            .I(timer_19));
    InMux I__2281 (
            .O(N__19860),
            .I(N__19857));
    LocalMux I__2280 (
            .O(N__19857),
            .I(N__19854));
    Span4Mux_h I__2279 (
            .O(N__19854),
            .I(N__19851));
    Span4Mux_v I__2278 (
            .O(N__19851),
            .I(N__19848));
    Span4Mux_v I__2277 (
            .O(N__19848),
            .I(N__19845));
    Odrv4 I__2276 (
            .O(N__19845),
            .I(pin_in_7));
    InMux I__2275 (
            .O(N__19842),
            .I(N__19839));
    LocalMux I__2274 (
            .O(N__19839),
            .I(N__19836));
    Span12Mux_v I__2273 (
            .O(N__19836),
            .I(N__19833));
    Odrv12 I__2272 (
            .O(N__19833),
            .I(pin_in_6));
    InMux I__2271 (
            .O(N__19830),
            .I(N__19827));
    LocalMux I__2270 (
            .O(N__19827),
            .I(\nx.n103 ));
    CascadeMux I__2269 (
            .O(N__19824),
            .I(N__19821));
    InMux I__2268 (
            .O(N__19821),
            .I(N__19818));
    LocalMux I__2267 (
            .O(N__19818),
            .I(\nx.n11892 ));
    InMux I__2266 (
            .O(N__19815),
            .I(N__19812));
    LocalMux I__2265 (
            .O(N__19812),
            .I(N__19809));
    Span4Mux_s3_h I__2264 (
            .O(N__19809),
            .I(N__19806));
    Odrv4 I__2263 (
            .O(N__19806),
            .I(\nx.n30_adj_712 ));
    InMux I__2262 (
            .O(N__19803),
            .I(N__19800));
    LocalMux I__2261 (
            .O(N__19800),
            .I(N__19797));
    Span4Mux_s3_h I__2260 (
            .O(N__19797),
            .I(N__19794));
    Odrv4 I__2259 (
            .O(N__19794),
            .I(\nx.n32 ));
    CascadeMux I__2258 (
            .O(N__19791),
            .I(N__19788));
    InMux I__2257 (
            .O(N__19788),
            .I(N__19785));
    LocalMux I__2256 (
            .O(N__19785),
            .I(N__19782));
    Span4Mux_v I__2255 (
            .O(N__19782),
            .I(N__19779));
    Sp12to4 I__2254 (
            .O(N__19779),
            .I(N__19776));
    Odrv12 I__2253 (
            .O(N__19776),
            .I(\nx.n28_adj_715 ));
    InMux I__2252 (
            .O(N__19773),
            .I(N__19768));
    InMux I__2251 (
            .O(N__19772),
            .I(N__19765));
    InMux I__2250 (
            .O(N__19771),
            .I(N__19762));
    LocalMux I__2249 (
            .O(N__19768),
            .I(timer_5));
    LocalMux I__2248 (
            .O(N__19765),
            .I(timer_5));
    LocalMux I__2247 (
            .O(N__19762),
            .I(timer_5));
    CascadeMux I__2246 (
            .O(N__19755),
            .I(N__19752));
    InMux I__2245 (
            .O(N__19752),
            .I(N__19746));
    InMux I__2244 (
            .O(N__19751),
            .I(N__19746));
    LocalMux I__2243 (
            .O(N__19746),
            .I(neo_pixel_transmitter_t0_5));
    CascadeMux I__2242 (
            .O(N__19743),
            .I(N__19738));
    InMux I__2241 (
            .O(N__19742),
            .I(N__19735));
    InMux I__2240 (
            .O(N__19741),
            .I(N__19732));
    InMux I__2239 (
            .O(N__19738),
            .I(N__19729));
    LocalMux I__2238 (
            .O(N__19735),
            .I(timer_1));
    LocalMux I__2237 (
            .O(N__19732),
            .I(timer_1));
    LocalMux I__2236 (
            .O(N__19729),
            .I(timer_1));
    CascadeMux I__2235 (
            .O(N__19722),
            .I(N__19719));
    InMux I__2234 (
            .O(N__19719),
            .I(N__19713));
    InMux I__2233 (
            .O(N__19718),
            .I(N__19713));
    LocalMux I__2232 (
            .O(N__19713),
            .I(neo_pixel_transmitter_t0_1));
    CascadeMux I__2231 (
            .O(N__19710),
            .I(N__19705));
    InMux I__2230 (
            .O(N__19709),
            .I(N__19702));
    InMux I__2229 (
            .O(N__19708),
            .I(N__19699));
    InMux I__2228 (
            .O(N__19705),
            .I(N__19696));
    LocalMux I__2227 (
            .O(N__19702),
            .I(timer_3));
    LocalMux I__2226 (
            .O(N__19699),
            .I(timer_3));
    LocalMux I__2225 (
            .O(N__19696),
            .I(timer_3));
    InMux I__2224 (
            .O(N__19689),
            .I(N__19685));
    InMux I__2223 (
            .O(N__19688),
            .I(N__19682));
    LocalMux I__2222 (
            .O(N__19685),
            .I(neo_pixel_transmitter_t0_3));
    LocalMux I__2221 (
            .O(N__19682),
            .I(neo_pixel_transmitter_t0_3));
    InMux I__2220 (
            .O(N__19677),
            .I(N__19674));
    LocalMux I__2219 (
            .O(N__19674),
            .I(\nx.n16_adj_785 ));
    CascadeMux I__2218 (
            .O(N__19671),
            .I(N__19667));
    InMux I__2217 (
            .O(N__19670),
            .I(N__19664));
    InMux I__2216 (
            .O(N__19667),
            .I(N__19661));
    LocalMux I__2215 (
            .O(N__19664),
            .I(N__19658));
    LocalMux I__2214 (
            .O(N__19661),
            .I(N__19655));
    Span4Mux_h I__2213 (
            .O(N__19658),
            .I(N__19652));
    Odrv4 I__2212 (
            .O(N__19655),
            .I(\nx.one_wire_N_599_4 ));
    Odrv4 I__2211 (
            .O(N__19652),
            .I(\nx.one_wire_N_599_4 ));
    InMux I__2210 (
            .O(N__19647),
            .I(N__19644));
    LocalMux I__2209 (
            .O(N__19644),
            .I(\nx.n46_adj_779 ));
    InMux I__2208 (
            .O(N__19641),
            .I(N__19638));
    LocalMux I__2207 (
            .O(N__19638),
            .I(N__19635));
    Span4Mux_v I__2206 (
            .O(N__19635),
            .I(N__19632));
    Span4Mux_v I__2205 (
            .O(N__19632),
            .I(N__19629));
    Odrv4 I__2204 (
            .O(N__19629),
            .I(\nx.n3 ));
    CascadeMux I__2203 (
            .O(N__19626),
            .I(\nx.n7_adj_764_cascade_ ));
    CascadeMux I__2202 (
            .O(N__19623),
            .I(\nx.n11864_cascade_ ));
    CEMux I__2201 (
            .O(N__19620),
            .I(N__19617));
    LocalMux I__2200 (
            .O(N__19617),
            .I(\nx.n7_adj_667 ));
    InMux I__2199 (
            .O(N__19614),
            .I(N__19611));
    LocalMux I__2198 (
            .O(N__19611),
            .I(\nx.n1476 ));
    CascadeMux I__2197 (
            .O(N__19608),
            .I(N__19604));
    InMux I__2196 (
            .O(N__19607),
            .I(N__19600));
    InMux I__2195 (
            .O(N__19604),
            .I(N__19597));
    InMux I__2194 (
            .O(N__19603),
            .I(N__19594));
    LocalMux I__2193 (
            .O(N__19600),
            .I(\nx.n1409 ));
    LocalMux I__2192 (
            .O(N__19597),
            .I(\nx.n1409 ));
    LocalMux I__2191 (
            .O(N__19594),
            .I(\nx.n1409 ));
    CascadeMux I__2190 (
            .O(N__19587),
            .I(N__19584));
    InMux I__2189 (
            .O(N__19584),
            .I(N__19581));
    LocalMux I__2188 (
            .O(N__19581),
            .I(\nx.n1468 ));
    InMux I__2187 (
            .O(N__19578),
            .I(N__19575));
    LocalMux I__2186 (
            .O(N__19575),
            .I(\nx.n1475 ));
    InMux I__2185 (
            .O(N__19572),
            .I(N__19568));
    CascadeMux I__2184 (
            .O(N__19571),
            .I(N__19565));
    LocalMux I__2183 (
            .O(N__19568),
            .I(N__19561));
    InMux I__2182 (
            .O(N__19565),
            .I(N__19558));
    InMux I__2181 (
            .O(N__19564),
            .I(N__19555));
    Odrv4 I__2180 (
            .O(N__19561),
            .I(\nx.n1408 ));
    LocalMux I__2179 (
            .O(N__19558),
            .I(\nx.n1408 ));
    LocalMux I__2178 (
            .O(N__19555),
            .I(\nx.n1408 ));
    CascadeMux I__2177 (
            .O(N__19548),
            .I(\nx.n1507_cascade_ ));
    CascadeMux I__2176 (
            .O(N__19545),
            .I(\nx.n18_adj_731_cascade_ ));
    CascadeMux I__2175 (
            .O(N__19542),
            .I(\nx.n20_adj_733_cascade_ ));
    InMux I__2174 (
            .O(N__19539),
            .I(N__19536));
    LocalMux I__2173 (
            .O(N__19536),
            .I(\nx.n16_adj_732 ));
    CascadeMux I__2172 (
            .O(N__19533),
            .I(\nx.n1532_cascade_ ));
    InMux I__2171 (
            .O(N__19530),
            .I(N__19527));
    LocalMux I__2170 (
            .O(N__19527),
            .I(N__19524));
    Odrv4 I__2169 (
            .O(N__19524),
            .I(\nx.n1477 ));
    CascadeMux I__2168 (
            .O(N__19521),
            .I(N__19515));
    CascadeMux I__2167 (
            .O(N__19520),
            .I(N__19510));
    CascadeMux I__2166 (
            .O(N__19519),
            .I(N__19506));
    CascadeMux I__2165 (
            .O(N__19518),
            .I(N__19502));
    InMux I__2164 (
            .O(N__19515),
            .I(N__19495));
    InMux I__2163 (
            .O(N__19514),
            .I(N__19495));
    InMux I__2162 (
            .O(N__19513),
            .I(N__19484));
    InMux I__2161 (
            .O(N__19510),
            .I(N__19484));
    InMux I__2160 (
            .O(N__19509),
            .I(N__19484));
    InMux I__2159 (
            .O(N__19506),
            .I(N__19484));
    InMux I__2158 (
            .O(N__19505),
            .I(N__19484));
    InMux I__2157 (
            .O(N__19502),
            .I(N__19477));
    InMux I__2156 (
            .O(N__19501),
            .I(N__19477));
    InMux I__2155 (
            .O(N__19500),
            .I(N__19477));
    LocalMux I__2154 (
            .O(N__19495),
            .I(\nx.n1433 ));
    LocalMux I__2153 (
            .O(N__19484),
            .I(\nx.n1433 ));
    LocalMux I__2152 (
            .O(N__19477),
            .I(\nx.n1433 ));
    CascadeMux I__2151 (
            .O(N__19470),
            .I(\nx.n1509_cascade_ ));
    InMux I__2150 (
            .O(N__19467),
            .I(N__19464));
    LocalMux I__2149 (
            .O(N__19464),
            .I(\nx.n9729 ));
    CascadeMux I__2148 (
            .O(N__19461),
            .I(\nx.n16_adj_727_cascade_ ));
    CascadeMux I__2147 (
            .O(N__19458),
            .I(N__19455));
    InMux I__2146 (
            .O(N__19455),
            .I(N__19452));
    LocalMux I__2145 (
            .O(N__19452),
            .I(\nx.n1471 ));
    InMux I__2144 (
            .O(N__19449),
            .I(N__19446));
    LocalMux I__2143 (
            .O(N__19446),
            .I(\nx.n1473 ));
    CascadeMux I__2142 (
            .O(N__19443),
            .I(N__19439));
    InMux I__2141 (
            .O(N__19442),
            .I(N__19435));
    InMux I__2140 (
            .O(N__19439),
            .I(N__19432));
    InMux I__2139 (
            .O(N__19438),
            .I(N__19429));
    LocalMux I__2138 (
            .O(N__19435),
            .I(\nx.n1406 ));
    LocalMux I__2137 (
            .O(N__19432),
            .I(\nx.n1406 ));
    LocalMux I__2136 (
            .O(N__19429),
            .I(\nx.n1406 ));
    CascadeMux I__2135 (
            .O(N__19422),
            .I(N__19419));
    InMux I__2134 (
            .O(N__19419),
            .I(N__19414));
    InMux I__2133 (
            .O(N__19418),
            .I(N__19409));
    InMux I__2132 (
            .O(N__19417),
            .I(N__19409));
    LocalMux I__2131 (
            .O(N__19414),
            .I(\nx.n1404 ));
    LocalMux I__2130 (
            .O(N__19409),
            .I(\nx.n1404 ));
    CascadeMux I__2129 (
            .O(N__19404),
            .I(N__19401));
    InMux I__2128 (
            .O(N__19401),
            .I(N__19398));
    LocalMux I__2127 (
            .O(N__19398),
            .I(\nx.n13_adj_729 ));
    InMux I__2126 (
            .O(N__19395),
            .I(N__19392));
    LocalMux I__2125 (
            .O(N__19392),
            .I(\nx.n18_adj_728 ));
    InMux I__2124 (
            .O(N__19389),
            .I(N__19384));
    InMux I__2123 (
            .O(N__19388),
            .I(N__19381));
    CascadeMux I__2122 (
            .O(N__19387),
            .I(N__19378));
    LocalMux I__2121 (
            .O(N__19384),
            .I(N__19373));
    LocalMux I__2120 (
            .O(N__19381),
            .I(N__19373));
    InMux I__2119 (
            .O(N__19378),
            .I(N__19370));
    Odrv4 I__2118 (
            .O(N__19373),
            .I(\nx.n1405 ));
    LocalMux I__2117 (
            .O(N__19370),
            .I(\nx.n1405 ));
    CascadeMux I__2116 (
            .O(N__19365),
            .I(\nx.n1433_cascade_ ));
    InMux I__2115 (
            .O(N__19362),
            .I(N__19359));
    LocalMux I__2114 (
            .O(N__19359),
            .I(\nx.n1472 ));
    InMux I__2113 (
            .O(N__19356),
            .I(N__19353));
    LocalMux I__2112 (
            .O(N__19353),
            .I(\nx.n1470 ));
    CascadeMux I__2111 (
            .O(N__19350),
            .I(N__19346));
    CascadeMux I__2110 (
            .O(N__19349),
            .I(N__19343));
    InMux I__2109 (
            .O(N__19346),
            .I(N__19340));
    InMux I__2108 (
            .O(N__19343),
            .I(N__19337));
    LocalMux I__2107 (
            .O(N__19340),
            .I(\nx.n1403 ));
    LocalMux I__2106 (
            .O(N__19337),
            .I(\nx.n1403 ));
    CascadeMux I__2105 (
            .O(N__19332),
            .I(\nx.n1502_cascade_ ));
    InMux I__2104 (
            .O(N__19329),
            .I(N__19326));
    LocalMux I__2103 (
            .O(N__19326),
            .I(\nx.n1474 ));
    CascadeMux I__2102 (
            .O(N__19323),
            .I(N__19319));
    CascadeMux I__2101 (
            .O(N__19322),
            .I(N__19315));
    InMux I__2100 (
            .O(N__19319),
            .I(N__19310));
    InMux I__2099 (
            .O(N__19318),
            .I(N__19310));
    InMux I__2098 (
            .O(N__19315),
            .I(N__19307));
    LocalMux I__2097 (
            .O(N__19310),
            .I(\nx.n1407 ));
    LocalMux I__2096 (
            .O(N__19307),
            .I(\nx.n1407 ));
    InMux I__2095 (
            .O(N__19302),
            .I(N__19299));
    LocalMux I__2094 (
            .O(N__19299),
            .I(N__19295));
    InMux I__2093 (
            .O(N__19298),
            .I(N__19292));
    Span4Mux_h I__2092 (
            .O(N__19295),
            .I(N__19289));
    LocalMux I__2091 (
            .O(N__19292),
            .I(delay_counter_21));
    Odrv4 I__2090 (
            .O(N__19289),
            .I(delay_counter_21));
    CascadeMux I__2089 (
            .O(N__19284),
            .I(N__19281));
    InMux I__2088 (
            .O(N__19281),
            .I(N__19278));
    LocalMux I__2087 (
            .O(N__19278),
            .I(N__19274));
    InMux I__2086 (
            .O(N__19277),
            .I(N__19271));
    Span4Mux_h I__2085 (
            .O(N__19274),
            .I(N__19268));
    LocalMux I__2084 (
            .O(N__19271),
            .I(delay_counter_29));
    Odrv4 I__2083 (
            .O(N__19268),
            .I(delay_counter_29));
    InMux I__2082 (
            .O(N__19263),
            .I(N__19260));
    LocalMux I__2081 (
            .O(N__19260),
            .I(n12379));
    InMux I__2080 (
            .O(N__19257),
            .I(N__19254));
    LocalMux I__2079 (
            .O(N__19254),
            .I(\nx.n12_adj_669 ));
    CascadeMux I__2078 (
            .O(N__19251),
            .I(\nx.n1308_cascade_ ));
    CascadeMux I__2077 (
            .O(N__19248),
            .I(\nx.n1334_cascade_ ));
    CascadeMux I__2076 (
            .O(N__19245),
            .I(\nx.n1403_cascade_ ));
    CascadeMux I__2075 (
            .O(N__19242),
            .I(N__19239));
    InMux I__2074 (
            .O(N__19239),
            .I(N__19233));
    InMux I__2073 (
            .O(N__19238),
            .I(N__19233));
    LocalMux I__2072 (
            .O(N__19233),
            .I(N__19229));
    InMux I__2071 (
            .O(N__19232),
            .I(N__19226));
    Odrv4 I__2070 (
            .O(N__19229),
            .I(\nx.n1402 ));
    LocalMux I__2069 (
            .O(N__19226),
            .I(\nx.n1402 ));
    InMux I__2068 (
            .O(N__19221),
            .I(N__19218));
    LocalMux I__2067 (
            .O(N__19218),
            .I(N__19214));
    InMux I__2066 (
            .O(N__19217),
            .I(N__19211));
    Span4Mux_h I__2065 (
            .O(N__19214),
            .I(N__19208));
    LocalMux I__2064 (
            .O(N__19211),
            .I(delay_counter_17));
    Odrv4 I__2063 (
            .O(N__19208),
            .I(delay_counter_17));
    CascadeMux I__2062 (
            .O(N__19203),
            .I(N__19200));
    InMux I__2061 (
            .O(N__19200),
            .I(N__19197));
    LocalMux I__2060 (
            .O(N__19197),
            .I(N__19193));
    InMux I__2059 (
            .O(N__19196),
            .I(N__19190));
    Span4Mux_h I__2058 (
            .O(N__19193),
            .I(N__19187));
    LocalMux I__2057 (
            .O(N__19190),
            .I(delay_counter_15));
    Odrv4 I__2056 (
            .O(N__19187),
            .I(delay_counter_15));
    InMux I__2055 (
            .O(N__19182),
            .I(N__19179));
    LocalMux I__2054 (
            .O(N__19179),
            .I(N__19176));
    Span4Mux_h I__2053 (
            .O(N__19176),
            .I(N__19173));
    Odrv4 I__2052 (
            .O(N__19173),
            .I(n12382));
    CascadeMux I__2051 (
            .O(N__19170),
            .I(n11828_cascade_));
    IoInMux I__2050 (
            .O(N__19167),
            .I(N__19164));
    LocalMux I__2049 (
            .O(N__19164),
            .I(N__19161));
    Span4Mux_s0_h I__2048 (
            .O(N__19161),
            .I(N__19158));
    Span4Mux_v I__2047 (
            .O(N__19158),
            .I(N__19155));
    Span4Mux_v I__2046 (
            .O(N__19155),
            .I(N__19151));
    InMux I__2045 (
            .O(N__19154),
            .I(N__19148));
    Odrv4 I__2044 (
            .O(N__19151),
            .I(pin_oe_5));
    LocalMux I__2043 (
            .O(N__19148),
            .I(pin_oe_5));
    InMux I__2042 (
            .O(N__19143),
            .I(N__19140));
    LocalMux I__2041 (
            .O(N__19140),
            .I(N__19135));
    InMux I__2040 (
            .O(N__19139),
            .I(N__19132));
    InMux I__2039 (
            .O(N__19138),
            .I(N__19129));
    Odrv4 I__2038 (
            .O(N__19135),
            .I(timer_16));
    LocalMux I__2037 (
            .O(N__19132),
            .I(timer_16));
    LocalMux I__2036 (
            .O(N__19129),
            .I(timer_16));
    InMux I__2035 (
            .O(N__19122),
            .I(N__19118));
    InMux I__2034 (
            .O(N__19121),
            .I(N__19115));
    LocalMux I__2033 (
            .O(N__19118),
            .I(neo_pixel_transmitter_t0_16));
    LocalMux I__2032 (
            .O(N__19115),
            .I(neo_pixel_transmitter_t0_16));
    CascadeMux I__2031 (
            .O(N__19110),
            .I(N__19107));
    InMux I__2030 (
            .O(N__19107),
            .I(N__19104));
    LocalMux I__2029 (
            .O(N__19104),
            .I(N__19101));
    Odrv4 I__2028 (
            .O(N__19101),
            .I(\nx.n17 ));
    CascadeMux I__2027 (
            .O(N__19098),
            .I(\nx.n1309_cascade_ ));
    InMux I__2026 (
            .O(N__19095),
            .I(\nx.n10731 ));
    InMux I__2025 (
            .O(N__19092),
            .I(\nx.n10732 ));
    CascadeMux I__2024 (
            .O(N__19089),
            .I(N__19085));
    InMux I__2023 (
            .O(N__19088),
            .I(N__19081));
    InMux I__2022 (
            .O(N__19085),
            .I(N__19078));
    InMux I__2021 (
            .O(N__19084),
            .I(N__19075));
    LocalMux I__2020 (
            .O(N__19081),
            .I(N__19070));
    LocalMux I__2019 (
            .O(N__19078),
            .I(N__19070));
    LocalMux I__2018 (
            .O(N__19075),
            .I(N__19065));
    Span4Mux_v I__2017 (
            .O(N__19070),
            .I(N__19065));
    Odrv4 I__2016 (
            .O(N__19065),
            .I(timer_27));
    InMux I__2015 (
            .O(N__19062),
            .I(\nx.n10733 ));
    InMux I__2014 (
            .O(N__19059),
            .I(\nx.n10734 ));
    InMux I__2013 (
            .O(N__19056),
            .I(\nx.n10735 ));
    InMux I__2012 (
            .O(N__19053),
            .I(\nx.n10736 ));
    InMux I__2011 (
            .O(N__19050),
            .I(\nx.n10737 ));
    InMux I__2010 (
            .O(N__19047),
            .I(N__19042));
    InMux I__2009 (
            .O(N__19046),
            .I(N__19039));
    InMux I__2008 (
            .O(N__19045),
            .I(N__19036));
    LocalMux I__2007 (
            .O(N__19042),
            .I(N__19033));
    LocalMux I__2006 (
            .O(N__19039),
            .I(N__19030));
    LocalMux I__2005 (
            .O(N__19036),
            .I(timer_31));
    Odrv12 I__2004 (
            .O(N__19033),
            .I(timer_31));
    Odrv4 I__2003 (
            .O(N__19030),
            .I(timer_31));
    CascadeMux I__2002 (
            .O(N__19023),
            .I(n11826_cascade_));
    IoInMux I__2001 (
            .O(N__19020),
            .I(N__19017));
    LocalMux I__2000 (
            .O(N__19017),
            .I(N__19014));
    Span4Mux_s2_v I__1999 (
            .O(N__19014),
            .I(N__19011));
    Span4Mux_v I__1998 (
            .O(N__19011),
            .I(N__19008));
    Span4Mux_v I__1997 (
            .O(N__19008),
            .I(N__19004));
    InMux I__1996 (
            .O(N__19007),
            .I(N__19001));
    Odrv4 I__1995 (
            .O(N__19004),
            .I(pin_oe_1));
    LocalMux I__1994 (
            .O(N__19001),
            .I(pin_oe_1));
    InMux I__1993 (
            .O(N__18996),
            .I(bfn_3_20_0_));
    InMux I__1992 (
            .O(N__18993),
            .I(N__18989));
    CascadeMux I__1991 (
            .O(N__18992),
            .I(N__18985));
    LocalMux I__1990 (
            .O(N__18989),
            .I(N__18982));
    InMux I__1989 (
            .O(N__18988),
            .I(N__18979));
    InMux I__1988 (
            .O(N__18985),
            .I(N__18976));
    Odrv4 I__1987 (
            .O(N__18982),
            .I(timer_17));
    LocalMux I__1986 (
            .O(N__18979),
            .I(timer_17));
    LocalMux I__1985 (
            .O(N__18976),
            .I(timer_17));
    InMux I__1984 (
            .O(N__18969),
            .I(\nx.n10723 ));
    InMux I__1983 (
            .O(N__18966),
            .I(N__18962));
    CascadeMux I__1982 (
            .O(N__18965),
            .I(N__18959));
    LocalMux I__1981 (
            .O(N__18962),
            .I(N__18955));
    InMux I__1980 (
            .O(N__18959),
            .I(N__18952));
    InMux I__1979 (
            .O(N__18958),
            .I(N__18949));
    Span4Mux_s2_h I__1978 (
            .O(N__18955),
            .I(N__18944));
    LocalMux I__1977 (
            .O(N__18952),
            .I(N__18944));
    LocalMux I__1976 (
            .O(N__18949),
            .I(timer_18));
    Odrv4 I__1975 (
            .O(N__18944),
            .I(timer_18));
    InMux I__1974 (
            .O(N__18939),
            .I(\nx.n10724 ));
    InMux I__1973 (
            .O(N__18936),
            .I(\nx.n10725 ));
    InMux I__1972 (
            .O(N__18933),
            .I(N__18930));
    LocalMux I__1971 (
            .O(N__18930),
            .I(N__18927));
    Span4Mux_s2_h I__1970 (
            .O(N__18927),
            .I(N__18922));
    InMux I__1969 (
            .O(N__18926),
            .I(N__18919));
    InMux I__1968 (
            .O(N__18925),
            .I(N__18916));
    Odrv4 I__1967 (
            .O(N__18922),
            .I(timer_20));
    LocalMux I__1966 (
            .O(N__18919),
            .I(timer_20));
    LocalMux I__1965 (
            .O(N__18916),
            .I(timer_20));
    InMux I__1964 (
            .O(N__18909),
            .I(\nx.n10726 ));
    InMux I__1963 (
            .O(N__18906),
            .I(N__18903));
    LocalMux I__1962 (
            .O(N__18903),
            .I(N__18899));
    InMux I__1961 (
            .O(N__18902),
            .I(N__18895));
    Span4Mux_v I__1960 (
            .O(N__18899),
            .I(N__18892));
    InMux I__1959 (
            .O(N__18898),
            .I(N__18889));
    LocalMux I__1958 (
            .O(N__18895),
            .I(N__18886));
    Odrv4 I__1957 (
            .O(N__18892),
            .I(timer_21));
    LocalMux I__1956 (
            .O(N__18889),
            .I(timer_21));
    Odrv4 I__1955 (
            .O(N__18886),
            .I(timer_21));
    InMux I__1954 (
            .O(N__18879),
            .I(\nx.n10727 ));
    InMux I__1953 (
            .O(N__18876),
            .I(N__18872));
    CascadeMux I__1952 (
            .O(N__18875),
            .I(N__18869));
    LocalMux I__1951 (
            .O(N__18872),
            .I(N__18865));
    InMux I__1950 (
            .O(N__18869),
            .I(N__18862));
    InMux I__1949 (
            .O(N__18868),
            .I(N__18859));
    Span4Mux_v I__1948 (
            .O(N__18865),
            .I(N__18854));
    LocalMux I__1947 (
            .O(N__18862),
            .I(N__18854));
    LocalMux I__1946 (
            .O(N__18859),
            .I(timer_22));
    Odrv4 I__1945 (
            .O(N__18854),
            .I(timer_22));
    InMux I__1944 (
            .O(N__18849),
            .I(\nx.n10728 ));
    InMux I__1943 (
            .O(N__18846),
            .I(N__18843));
    LocalMux I__1942 (
            .O(N__18843),
            .I(N__18838));
    InMux I__1941 (
            .O(N__18842),
            .I(N__18835));
    InMux I__1940 (
            .O(N__18841),
            .I(N__18832));
    Span4Mux_v I__1939 (
            .O(N__18838),
            .I(N__18827));
    LocalMux I__1938 (
            .O(N__18835),
            .I(N__18827));
    LocalMux I__1937 (
            .O(N__18832),
            .I(timer_23));
    Odrv4 I__1936 (
            .O(N__18827),
            .I(timer_23));
    InMux I__1935 (
            .O(N__18822),
            .I(\nx.n10729 ));
    InMux I__1934 (
            .O(N__18819),
            .I(N__18815));
    CascadeMux I__1933 (
            .O(N__18818),
            .I(N__18811));
    LocalMux I__1932 (
            .O(N__18815),
            .I(N__18808));
    InMux I__1931 (
            .O(N__18814),
            .I(N__18805));
    InMux I__1930 (
            .O(N__18811),
            .I(N__18802));
    Odrv4 I__1929 (
            .O(N__18808),
            .I(timer_24));
    LocalMux I__1928 (
            .O(N__18805),
            .I(timer_24));
    LocalMux I__1927 (
            .O(N__18802),
            .I(timer_24));
    InMux I__1926 (
            .O(N__18795),
            .I(bfn_3_21_0_));
    InMux I__1925 (
            .O(N__18792),
            .I(N__18789));
    LocalMux I__1924 (
            .O(N__18789),
            .I(N__18784));
    InMux I__1923 (
            .O(N__18788),
            .I(N__18781));
    InMux I__1922 (
            .O(N__18787),
            .I(N__18778));
    Odrv4 I__1921 (
            .O(N__18784),
            .I(timer_8));
    LocalMux I__1920 (
            .O(N__18781),
            .I(timer_8));
    LocalMux I__1919 (
            .O(N__18778),
            .I(timer_8));
    InMux I__1918 (
            .O(N__18771),
            .I(bfn_3_19_0_));
    InMux I__1917 (
            .O(N__18768),
            .I(N__18765));
    LocalMux I__1916 (
            .O(N__18765),
            .I(N__18760));
    InMux I__1915 (
            .O(N__18764),
            .I(N__18757));
    InMux I__1914 (
            .O(N__18763),
            .I(N__18754));
    Odrv4 I__1913 (
            .O(N__18760),
            .I(timer_9));
    LocalMux I__1912 (
            .O(N__18757),
            .I(timer_9));
    LocalMux I__1911 (
            .O(N__18754),
            .I(timer_9));
    InMux I__1910 (
            .O(N__18747),
            .I(\nx.n10715 ));
    InMux I__1909 (
            .O(N__18744),
            .I(N__18740));
    CascadeMux I__1908 (
            .O(N__18743),
            .I(N__18736));
    LocalMux I__1907 (
            .O(N__18740),
            .I(N__18733));
    InMux I__1906 (
            .O(N__18739),
            .I(N__18730));
    InMux I__1905 (
            .O(N__18736),
            .I(N__18727));
    Odrv4 I__1904 (
            .O(N__18733),
            .I(timer_10));
    LocalMux I__1903 (
            .O(N__18730),
            .I(timer_10));
    LocalMux I__1902 (
            .O(N__18727),
            .I(timer_10));
    InMux I__1901 (
            .O(N__18720),
            .I(\nx.n10716 ));
    InMux I__1900 (
            .O(N__18717),
            .I(\nx.n10717 ));
    InMux I__1899 (
            .O(N__18714),
            .I(N__18711));
    LocalMux I__1898 (
            .O(N__18711),
            .I(N__18707));
    CascadeMux I__1897 (
            .O(N__18710),
            .I(N__18703));
    Span4Mux_s2_h I__1896 (
            .O(N__18707),
            .I(N__18700));
    InMux I__1895 (
            .O(N__18706),
            .I(N__18697));
    InMux I__1894 (
            .O(N__18703),
            .I(N__18694));
    Odrv4 I__1893 (
            .O(N__18700),
            .I(timer_12));
    LocalMux I__1892 (
            .O(N__18697),
            .I(timer_12));
    LocalMux I__1891 (
            .O(N__18694),
            .I(timer_12));
    InMux I__1890 (
            .O(N__18687),
            .I(\nx.n10718 ));
    InMux I__1889 (
            .O(N__18684),
            .I(\nx.n10719 ));
    InMux I__1888 (
            .O(N__18681),
            .I(N__18677));
    CascadeMux I__1887 (
            .O(N__18680),
            .I(N__18673));
    LocalMux I__1886 (
            .O(N__18677),
            .I(N__18670));
    InMux I__1885 (
            .O(N__18676),
            .I(N__18667));
    InMux I__1884 (
            .O(N__18673),
            .I(N__18664));
    Odrv12 I__1883 (
            .O(N__18670),
            .I(timer_14));
    LocalMux I__1882 (
            .O(N__18667),
            .I(timer_14));
    LocalMux I__1881 (
            .O(N__18664),
            .I(timer_14));
    InMux I__1880 (
            .O(N__18657),
            .I(\nx.n10720 ));
    InMux I__1879 (
            .O(N__18654),
            .I(N__18651));
    LocalMux I__1878 (
            .O(N__18651),
            .I(N__18646));
    InMux I__1877 (
            .O(N__18650),
            .I(N__18643));
    InMux I__1876 (
            .O(N__18649),
            .I(N__18640));
    Span4Mux_v I__1875 (
            .O(N__18646),
            .I(N__18635));
    LocalMux I__1874 (
            .O(N__18643),
            .I(N__18635));
    LocalMux I__1873 (
            .O(N__18640),
            .I(timer_15));
    Odrv4 I__1872 (
            .O(N__18635),
            .I(timer_15));
    InMux I__1871 (
            .O(N__18630),
            .I(\nx.n10721 ));
    CascadeMux I__1870 (
            .O(N__18627),
            .I(\nx.n11834_cascade_ ));
    InMux I__1869 (
            .O(N__18624),
            .I(N__18621));
    LocalMux I__1868 (
            .O(N__18621),
            .I(N__18617));
    CascadeMux I__1867 (
            .O(N__18620),
            .I(N__18613));
    Span4Mux_v I__1866 (
            .O(N__18617),
            .I(N__18610));
    InMux I__1865 (
            .O(N__18616),
            .I(N__18607));
    InMux I__1864 (
            .O(N__18613),
            .I(N__18604));
    Odrv4 I__1863 (
            .O(N__18610),
            .I(timer_0));
    LocalMux I__1862 (
            .O(N__18607),
            .I(timer_0));
    LocalMux I__1861 (
            .O(N__18604),
            .I(timer_0));
    InMux I__1860 (
            .O(N__18597),
            .I(bfn_3_18_0_));
    InMux I__1859 (
            .O(N__18594),
            .I(\nx.n10707 ));
    CascadeMux I__1858 (
            .O(N__18591),
            .I(N__18586));
    InMux I__1857 (
            .O(N__18590),
            .I(N__18583));
    InMux I__1856 (
            .O(N__18589),
            .I(N__18580));
    InMux I__1855 (
            .O(N__18586),
            .I(N__18577));
    LocalMux I__1854 (
            .O(N__18583),
            .I(timer_2));
    LocalMux I__1853 (
            .O(N__18580),
            .I(timer_2));
    LocalMux I__1852 (
            .O(N__18577),
            .I(timer_2));
    InMux I__1851 (
            .O(N__18570),
            .I(\nx.n10708 ));
    InMux I__1850 (
            .O(N__18567),
            .I(\nx.n10709 ));
    InMux I__1849 (
            .O(N__18564),
            .I(N__18560));
    CascadeMux I__1848 (
            .O(N__18563),
            .I(N__18556));
    LocalMux I__1847 (
            .O(N__18560),
            .I(N__18553));
    InMux I__1846 (
            .O(N__18559),
            .I(N__18550));
    InMux I__1845 (
            .O(N__18556),
            .I(N__18547));
    Odrv4 I__1844 (
            .O(N__18553),
            .I(timer_4));
    LocalMux I__1843 (
            .O(N__18550),
            .I(timer_4));
    LocalMux I__1842 (
            .O(N__18547),
            .I(timer_4));
    InMux I__1841 (
            .O(N__18540),
            .I(\nx.n10710 ));
    InMux I__1840 (
            .O(N__18537),
            .I(\nx.n10711 ));
    CascadeMux I__1839 (
            .O(N__18534),
            .I(N__18529));
    InMux I__1838 (
            .O(N__18533),
            .I(N__18526));
    InMux I__1837 (
            .O(N__18532),
            .I(N__18523));
    InMux I__1836 (
            .O(N__18529),
            .I(N__18520));
    LocalMux I__1835 (
            .O(N__18526),
            .I(timer_6));
    LocalMux I__1834 (
            .O(N__18523),
            .I(timer_6));
    LocalMux I__1833 (
            .O(N__18520),
            .I(timer_6));
    InMux I__1832 (
            .O(N__18513),
            .I(\nx.n10712 ));
    InMux I__1831 (
            .O(N__18510),
            .I(N__18506));
    CascadeMux I__1830 (
            .O(N__18509),
            .I(N__18502));
    LocalMux I__1829 (
            .O(N__18506),
            .I(N__18499));
    InMux I__1828 (
            .O(N__18505),
            .I(N__18496));
    InMux I__1827 (
            .O(N__18502),
            .I(N__18493));
    Odrv4 I__1826 (
            .O(N__18499),
            .I(timer_7));
    LocalMux I__1825 (
            .O(N__18496),
            .I(timer_7));
    LocalMux I__1824 (
            .O(N__18493),
            .I(timer_7));
    InMux I__1823 (
            .O(N__18486),
            .I(\nx.n10713 ));
    InMux I__1822 (
            .O(N__18483),
            .I(bfn_2_26_0_));
    InMux I__1821 (
            .O(N__18480),
            .I(\nx.n10781 ));
    InMux I__1820 (
            .O(N__18477),
            .I(\nx.n10782 ));
    InMux I__1819 (
            .O(N__18474),
            .I(N__18471));
    LocalMux I__1818 (
            .O(N__18471),
            .I(\nx.n1469 ));
    InMux I__1817 (
            .O(N__18468),
            .I(N__18462));
    InMux I__1816 (
            .O(N__18467),
            .I(N__18462));
    LocalMux I__1815 (
            .O(N__18462),
            .I(neo_pixel_transmitter_t0_14));
    InMux I__1814 (
            .O(N__18459),
            .I(N__18456));
    LocalMux I__1813 (
            .O(N__18456),
            .I(N__18453));
    Span4Mux_v I__1812 (
            .O(N__18453),
            .I(N__18450));
    Odrv4 I__1811 (
            .O(N__18450),
            .I(\nx.n19_adj_725 ));
    InMux I__1810 (
            .O(N__18447),
            .I(bfn_2_25_0_));
    InMux I__1809 (
            .O(N__18444),
            .I(\nx.n10773 ));
    InMux I__1808 (
            .O(N__18441),
            .I(\nx.n10774 ));
    InMux I__1807 (
            .O(N__18438),
            .I(\nx.n10775 ));
    InMux I__1806 (
            .O(N__18435),
            .I(\nx.n10776 ));
    InMux I__1805 (
            .O(N__18432),
            .I(\nx.n10777 ));
    InMux I__1804 (
            .O(N__18429),
            .I(\nx.n10778 ));
    InMux I__1803 (
            .O(N__18426),
            .I(\nx.n10779 ));
    InMux I__1802 (
            .O(N__18423),
            .I(N__18420));
    LocalMux I__1801 (
            .O(N__18420),
            .I(\nx.n13201 ));
    InMux I__1800 (
            .O(N__18417),
            .I(bfn_2_23_0_));
    InMux I__1799 (
            .O(N__18414),
            .I(N__18411));
    LocalMux I__1798 (
            .O(N__18411),
            .I(\nx.n13203 ));
    InMux I__1797 (
            .O(N__18408),
            .I(\nx.n10696 ));
    InMux I__1796 (
            .O(N__18405),
            .I(N__18402));
    LocalMux I__1795 (
            .O(N__18402),
            .I(\nx.n13205 ));
    InMux I__1794 (
            .O(N__18399),
            .I(N__18396));
    LocalMux I__1793 (
            .O(N__18396),
            .I(N__18393));
    Span4Mux_v I__1792 (
            .O(N__18393),
            .I(N__18390));
    Odrv4 I__1791 (
            .O(N__18390),
            .I(\nx.n4_adj_710 ));
    InMux I__1790 (
            .O(N__18387),
            .I(\nx.n10697 ));
    InMux I__1789 (
            .O(N__18384),
            .I(N__18381));
    LocalMux I__1788 (
            .O(N__18381),
            .I(\nx.n13207 ));
    InMux I__1787 (
            .O(N__18378),
            .I(\nx.n10698 ));
    InMux I__1786 (
            .O(N__18375),
            .I(N__18372));
    LocalMux I__1785 (
            .O(N__18372),
            .I(N__18369));
    Odrv4 I__1784 (
            .O(N__18369),
            .I(\nx.n2 ));
    CascadeMux I__1783 (
            .O(N__18366),
            .I(N__18363));
    InMux I__1782 (
            .O(N__18363),
            .I(N__18360));
    LocalMux I__1781 (
            .O(N__18360),
            .I(\nx.n13209 ));
    InMux I__1780 (
            .O(N__18357),
            .I(\nx.n10699 ));
    InMux I__1779 (
            .O(N__18354),
            .I(N__18351));
    LocalMux I__1778 (
            .O(N__18351),
            .I(\nx.n6 ));
    InMux I__1777 (
            .O(N__18348),
            .I(N__18342));
    InMux I__1776 (
            .O(N__18347),
            .I(N__18342));
    LocalMux I__1775 (
            .O(N__18342),
            .I(neo_pixel_transmitter_t0_27));
    InMux I__1774 (
            .O(N__18339),
            .I(N__18336));
    LocalMux I__1773 (
            .O(N__18336),
            .I(\nx.n13189 ));
    CascadeMux I__1772 (
            .O(N__18333),
            .I(N__18330));
    InMux I__1771 (
            .O(N__18330),
            .I(N__18327));
    LocalMux I__1770 (
            .O(N__18327),
            .I(N__18324));
    Span4Mux_v I__1769 (
            .O(N__18324),
            .I(N__18321));
    Odrv4 I__1768 (
            .O(N__18321),
            .I(\nx.n12 ));
    InMux I__1767 (
            .O(N__18318),
            .I(bfn_2_22_0_));
    InMux I__1766 (
            .O(N__18315),
            .I(N__18312));
    LocalMux I__1765 (
            .O(N__18312),
            .I(\nx.n13191 ));
    InMux I__1764 (
            .O(N__18309),
            .I(N__18306));
    LocalMux I__1763 (
            .O(N__18306),
            .I(N__18303));
    Odrv12 I__1762 (
            .O(N__18303),
            .I(\nx.n11 ));
    InMux I__1761 (
            .O(N__18300),
            .I(\nx.n10690 ));
    InMux I__1760 (
            .O(N__18297),
            .I(N__18294));
    LocalMux I__1759 (
            .O(N__18294),
            .I(\nx.n13193 ));
    CascadeMux I__1758 (
            .O(N__18291),
            .I(N__18288));
    InMux I__1757 (
            .O(N__18288),
            .I(N__18285));
    LocalMux I__1756 (
            .O(N__18285),
            .I(N__18282));
    Odrv12 I__1755 (
            .O(N__18282),
            .I(\nx.n10 ));
    InMux I__1754 (
            .O(N__18279),
            .I(\nx.n10691 ));
    InMux I__1753 (
            .O(N__18276),
            .I(N__18273));
    LocalMux I__1752 (
            .O(N__18273),
            .I(N__18270));
    Odrv4 I__1751 (
            .O(N__18270),
            .I(\nx.n13195 ));
    InMux I__1750 (
            .O(N__18267),
            .I(N__18264));
    LocalMux I__1749 (
            .O(N__18264),
            .I(\nx.n9 ));
    InMux I__1748 (
            .O(N__18261),
            .I(\nx.n10692 ));
    InMux I__1747 (
            .O(N__18258),
            .I(N__18255));
    LocalMux I__1746 (
            .O(N__18255),
            .I(N__18252));
    Odrv4 I__1745 (
            .O(N__18252),
            .I(\nx.n13197 ));
    InMux I__1744 (
            .O(N__18249),
            .I(\nx.n10693 ));
    InMux I__1743 (
            .O(N__18246),
            .I(N__18243));
    LocalMux I__1742 (
            .O(N__18243),
            .I(N__18240));
    Odrv4 I__1741 (
            .O(N__18240),
            .I(\nx.n13199 ));
    InMux I__1740 (
            .O(N__18237),
            .I(\nx.n10694 ));
    InMux I__1739 (
            .O(N__18234),
            .I(N__18231));
    LocalMux I__1738 (
            .O(N__18231),
            .I(\nx.n13177 ));
    CascadeMux I__1737 (
            .O(N__18228),
            .I(N__18225));
    InMux I__1736 (
            .O(N__18225),
            .I(N__18222));
    LocalMux I__1735 (
            .O(N__18222),
            .I(N__18219));
    Odrv12 I__1734 (
            .O(N__18219),
            .I(\nx.n18_adj_723 ));
    InMux I__1733 (
            .O(N__18216),
            .I(bfn_2_21_0_));
    InMux I__1732 (
            .O(N__18213),
            .I(N__18210));
    LocalMux I__1731 (
            .O(N__18210),
            .I(\nx.n13179 ));
    InMux I__1730 (
            .O(N__18207),
            .I(\nx.n10684 ));
    InMux I__1729 (
            .O(N__18204),
            .I(N__18201));
    LocalMux I__1728 (
            .O(N__18201),
            .I(\nx.n13181 ));
    InMux I__1727 (
            .O(N__18198),
            .I(N__18195));
    LocalMux I__1726 (
            .O(N__18195),
            .I(N__18192));
    Odrv4 I__1725 (
            .O(N__18192),
            .I(\nx.n16_adj_672 ));
    InMux I__1724 (
            .O(N__18189),
            .I(\nx.n10685 ));
    InMux I__1723 (
            .O(N__18186),
            .I(N__18183));
    LocalMux I__1722 (
            .O(N__18183),
            .I(N__18180));
    Odrv4 I__1721 (
            .O(N__18180),
            .I(\nx.n13183 ));
    InMux I__1720 (
            .O(N__18177),
            .I(N__18174));
    LocalMux I__1719 (
            .O(N__18174),
            .I(\nx.n15 ));
    InMux I__1718 (
            .O(N__18171),
            .I(\nx.n10686 ));
    InMux I__1717 (
            .O(N__18168),
            .I(N__18165));
    LocalMux I__1716 (
            .O(N__18165),
            .I(\nx.n13185 ));
    InMux I__1715 (
            .O(N__18162),
            .I(\nx.n10687 ));
    InMux I__1714 (
            .O(N__18159),
            .I(N__18156));
    LocalMux I__1713 (
            .O(N__18156),
            .I(N__18153));
    Odrv4 I__1712 (
            .O(N__18153),
            .I(\nx.n13187 ));
    CascadeMux I__1711 (
            .O(N__18150),
            .I(N__18147));
    InMux I__1710 (
            .O(N__18147),
            .I(N__18144));
    LocalMux I__1709 (
            .O(N__18144),
            .I(\nx.n13 ));
    InMux I__1708 (
            .O(N__18141),
            .I(\nx.n10688 ));
    InMux I__1707 (
            .O(N__18138),
            .I(N__18135));
    LocalMux I__1706 (
            .O(N__18135),
            .I(\nx.n26_adj_722 ));
    InMux I__1705 (
            .O(N__18132),
            .I(\nx.n10675 ));
    CascadeMux I__1704 (
            .O(N__18129),
            .I(N__18126));
    InMux I__1703 (
            .O(N__18126),
            .I(N__18123));
    LocalMux I__1702 (
            .O(N__18123),
            .I(N__18120));
    Odrv12 I__1701 (
            .O(N__18120),
            .I(\nx.n25_adj_724 ));
    InMux I__1700 (
            .O(N__18117),
            .I(bfn_2_20_0_));
    CascadeMux I__1699 (
            .O(N__18114),
            .I(N__18111));
    InMux I__1698 (
            .O(N__18111),
            .I(N__18108));
    LocalMux I__1697 (
            .O(N__18108),
            .I(\nx.n24_adj_734 ));
    InMux I__1696 (
            .O(N__18105),
            .I(\nx.n10677 ));
    InMux I__1695 (
            .O(N__18102),
            .I(N__18099));
    LocalMux I__1694 (
            .O(N__18099),
            .I(N__18096));
    Odrv4 I__1693 (
            .O(N__18096),
            .I(\nx.n23 ));
    InMux I__1692 (
            .O(N__18093),
            .I(\nx.n10678 ));
    InMux I__1691 (
            .O(N__18090),
            .I(\nx.n10679 ));
    InMux I__1690 (
            .O(N__18087),
            .I(N__18084));
    LocalMux I__1689 (
            .O(N__18084),
            .I(\nx.one_wire_N_599_11 ));
    InMux I__1688 (
            .O(N__18081),
            .I(N__18078));
    LocalMux I__1687 (
            .O(N__18078),
            .I(N__18075));
    Span4Mux_h I__1686 (
            .O(N__18075),
            .I(N__18072));
    Odrv4 I__1685 (
            .O(N__18072),
            .I(\nx.n21_adj_737 ));
    InMux I__1684 (
            .O(N__18069),
            .I(\nx.n10680 ));
    InMux I__1683 (
            .O(N__18066),
            .I(N__18063));
    LocalMux I__1682 (
            .O(N__18063),
            .I(\nx.n13173 ));
    InMux I__1681 (
            .O(N__18060),
            .I(\nx.n10681 ));
    InMux I__1680 (
            .O(N__18057),
            .I(N__18054));
    LocalMux I__1679 (
            .O(N__18054),
            .I(\nx.n13175 ));
    InMux I__1678 (
            .O(N__18051),
            .I(\nx.n10682 ));
    InMux I__1677 (
            .O(N__18048),
            .I(N__18042));
    InMux I__1676 (
            .O(N__18047),
            .I(N__18042));
    LocalMux I__1675 (
            .O(N__18042),
            .I(neo_pixel_transmitter_t0_22));
    InMux I__1674 (
            .O(N__18039),
            .I(N__18033));
    InMux I__1673 (
            .O(N__18038),
            .I(N__18033));
    LocalMux I__1672 (
            .O(N__18033),
            .I(neo_pixel_transmitter_t0_10));
    InMux I__1671 (
            .O(N__18030),
            .I(N__18027));
    LocalMux I__1670 (
            .O(N__18027),
            .I(N__18024));
    Odrv4 I__1669 (
            .O(N__18024),
            .I(\nx.n33 ));
    InMux I__1668 (
            .O(N__18021),
            .I(\nx.n10669 ));
    InMux I__1667 (
            .O(N__18018),
            .I(N__18015));
    LocalMux I__1666 (
            .O(N__18015),
            .I(N__18012));
    Odrv4 I__1665 (
            .O(N__18012),
            .I(\nx.n31_adj_711 ));
    InMux I__1664 (
            .O(N__18009),
            .I(\nx.n10670 ));
    InMux I__1663 (
            .O(N__18006),
            .I(\nx.n10671 ));
    InMux I__1662 (
            .O(N__18003),
            .I(N__18000));
    LocalMux I__1661 (
            .O(N__18000),
            .I(\nx.n29_adj_714 ));
    InMux I__1660 (
            .O(N__17997),
            .I(\nx.n10672 ));
    InMux I__1659 (
            .O(N__17994),
            .I(\nx.n10673 ));
    InMux I__1658 (
            .O(N__17991),
            .I(N__17988));
    LocalMux I__1657 (
            .O(N__17988),
            .I(\nx.n27_adj_720 ));
    InMux I__1656 (
            .O(N__17985),
            .I(\nx.n10674 ));
    InMux I__1655 (
            .O(N__17982),
            .I(N__17976));
    InMux I__1654 (
            .O(N__17981),
            .I(N__17976));
    LocalMux I__1653 (
            .O(N__17976),
            .I(neo_pixel_transmitter_t0_23));
    InMux I__1652 (
            .O(N__17973),
            .I(N__17967));
    InMux I__1651 (
            .O(N__17972),
            .I(N__17967));
    LocalMux I__1650 (
            .O(N__17967),
            .I(neo_pixel_transmitter_t0_15));
    InMux I__1649 (
            .O(N__17964),
            .I(N__17958));
    InMux I__1648 (
            .O(N__17963),
            .I(N__17958));
    LocalMux I__1647 (
            .O(N__17958),
            .I(neo_pixel_transmitter_t0_8));
    InMux I__1646 (
            .O(N__17955),
            .I(N__17949));
    InMux I__1645 (
            .O(N__17954),
            .I(N__17949));
    LocalMux I__1644 (
            .O(N__17949),
            .I(neo_pixel_transmitter_t0_2));
    InMux I__1643 (
            .O(N__17946),
            .I(N__17942));
    InMux I__1642 (
            .O(N__17945),
            .I(N__17939));
    LocalMux I__1641 (
            .O(N__17942),
            .I(neo_pixel_transmitter_t0_6));
    LocalMux I__1640 (
            .O(N__17939),
            .I(neo_pixel_transmitter_t0_6));
    InMux I__1639 (
            .O(N__17934),
            .I(N__17928));
    InMux I__1638 (
            .O(N__17933),
            .I(N__17928));
    LocalMux I__1637 (
            .O(N__17928),
            .I(neo_pixel_transmitter_t0_17));
    InMux I__1636 (
            .O(N__17925),
            .I(N__17921));
    InMux I__1635 (
            .O(N__17924),
            .I(N__17918));
    LocalMux I__1634 (
            .O(N__17921),
            .I(N__17915));
    LocalMux I__1633 (
            .O(N__17918),
            .I(delay_counter_27));
    Odrv12 I__1632 (
            .O(N__17915),
            .I(delay_counter_27));
    InMux I__1631 (
            .O(N__17910),
            .I(n10608));
    InMux I__1630 (
            .O(N__17907),
            .I(n10609));
    InMux I__1629 (
            .O(N__17904),
            .I(n10610));
    InMux I__1628 (
            .O(N__17901),
            .I(N__17897));
    InMux I__1627 (
            .O(N__17900),
            .I(N__17894));
    LocalMux I__1626 (
            .O(N__17897),
            .I(N__17891));
    LocalMux I__1625 (
            .O(N__17894),
            .I(delay_counter_30));
    Odrv12 I__1624 (
            .O(N__17891),
            .I(delay_counter_30));
    InMux I__1623 (
            .O(N__17886),
            .I(n10611));
    InMux I__1622 (
            .O(N__17883),
            .I(n10612));
    InMux I__1621 (
            .O(N__17880),
            .I(n10599));
    InMux I__1620 (
            .O(N__17877),
            .I(n10600));
    InMux I__1619 (
            .O(N__17874),
            .I(n10601));
    InMux I__1618 (
            .O(N__17871),
            .I(n10602));
    InMux I__1617 (
            .O(N__17868),
            .I(n10603));
    CascadeMux I__1616 (
            .O(N__17865),
            .I(N__17862));
    InMux I__1615 (
            .O(N__17862),
            .I(N__17858));
    InMux I__1614 (
            .O(N__17861),
            .I(N__17855));
    LocalMux I__1613 (
            .O(N__17858),
            .I(N__17852));
    LocalMux I__1612 (
            .O(N__17855),
            .I(delay_counter_23));
    Odrv12 I__1611 (
            .O(N__17852),
            .I(delay_counter_23));
    InMux I__1610 (
            .O(N__17847),
            .I(n10604));
    InMux I__1609 (
            .O(N__17844),
            .I(bfn_1_25_0_));
    InMux I__1608 (
            .O(N__17841),
            .I(N__17837));
    InMux I__1607 (
            .O(N__17840),
            .I(N__17834));
    LocalMux I__1606 (
            .O(N__17837),
            .I(N__17831));
    LocalMux I__1605 (
            .O(N__17834),
            .I(delay_counter_25));
    Odrv12 I__1604 (
            .O(N__17831),
            .I(delay_counter_25));
    InMux I__1603 (
            .O(N__17826),
            .I(n10606));
    InMux I__1602 (
            .O(N__17823),
            .I(n10607));
    CascadeMux I__1601 (
            .O(N__17820),
            .I(N__17817));
    InMux I__1600 (
            .O(N__17817),
            .I(N__17813));
    InMux I__1599 (
            .O(N__17816),
            .I(N__17810));
    LocalMux I__1598 (
            .O(N__17813),
            .I(N__17807));
    LocalMux I__1597 (
            .O(N__17810),
            .I(delay_counter_9));
    Odrv4 I__1596 (
            .O(N__17807),
            .I(delay_counter_9));
    InMux I__1595 (
            .O(N__17802),
            .I(n10590));
    InMux I__1594 (
            .O(N__17799),
            .I(N__17795));
    InMux I__1593 (
            .O(N__17798),
            .I(N__17792));
    LocalMux I__1592 (
            .O(N__17795),
            .I(N__17789));
    LocalMux I__1591 (
            .O(N__17792),
            .I(delay_counter_10));
    Odrv4 I__1590 (
            .O(N__17789),
            .I(delay_counter_10));
    InMux I__1589 (
            .O(N__17784),
            .I(n10591));
    InMux I__1588 (
            .O(N__17781),
            .I(N__17777));
    InMux I__1587 (
            .O(N__17780),
            .I(N__17774));
    LocalMux I__1586 (
            .O(N__17777),
            .I(N__17771));
    LocalMux I__1585 (
            .O(N__17774),
            .I(delay_counter_11));
    Odrv4 I__1584 (
            .O(N__17771),
            .I(delay_counter_11));
    InMux I__1583 (
            .O(N__17766),
            .I(n10592));
    InMux I__1582 (
            .O(N__17763),
            .I(N__17759));
    InMux I__1581 (
            .O(N__17762),
            .I(N__17756));
    LocalMux I__1580 (
            .O(N__17759),
            .I(N__17753));
    LocalMux I__1579 (
            .O(N__17756),
            .I(delay_counter_12));
    Odrv4 I__1578 (
            .O(N__17753),
            .I(delay_counter_12));
    InMux I__1577 (
            .O(N__17748),
            .I(n10593));
    InMux I__1576 (
            .O(N__17745),
            .I(N__17741));
    InMux I__1575 (
            .O(N__17744),
            .I(N__17738));
    LocalMux I__1574 (
            .O(N__17741),
            .I(N__17735));
    LocalMux I__1573 (
            .O(N__17738),
            .I(delay_counter_13));
    Odrv4 I__1572 (
            .O(N__17735),
            .I(delay_counter_13));
    InMux I__1571 (
            .O(N__17730),
            .I(n10594));
    InMux I__1570 (
            .O(N__17727),
            .I(N__17723));
    InMux I__1569 (
            .O(N__17726),
            .I(N__17720));
    LocalMux I__1568 (
            .O(N__17723),
            .I(N__17717));
    LocalMux I__1567 (
            .O(N__17720),
            .I(delay_counter_14));
    Odrv12 I__1566 (
            .O(N__17717),
            .I(delay_counter_14));
    InMux I__1565 (
            .O(N__17712),
            .I(n10595));
    InMux I__1564 (
            .O(N__17709),
            .I(n10596));
    InMux I__1563 (
            .O(N__17706),
            .I(bfn_1_24_0_));
    InMux I__1562 (
            .O(N__17703),
            .I(n10598));
    InMux I__1561 (
            .O(N__17700),
            .I(N__17696));
    InMux I__1560 (
            .O(N__17699),
            .I(N__17693));
    LocalMux I__1559 (
            .O(N__17696),
            .I(delay_counter_1));
    LocalMux I__1558 (
            .O(N__17693),
            .I(delay_counter_1));
    InMux I__1557 (
            .O(N__17688),
            .I(n10582));
    CascadeMux I__1556 (
            .O(N__17685),
            .I(N__17681));
    InMux I__1555 (
            .O(N__17684),
            .I(N__17678));
    InMux I__1554 (
            .O(N__17681),
            .I(N__17675));
    LocalMux I__1553 (
            .O(N__17678),
            .I(delay_counter_2));
    LocalMux I__1552 (
            .O(N__17675),
            .I(delay_counter_2));
    InMux I__1551 (
            .O(N__17670),
            .I(n10583));
    InMux I__1550 (
            .O(N__17667),
            .I(N__17663));
    InMux I__1549 (
            .O(N__17666),
            .I(N__17660));
    LocalMux I__1548 (
            .O(N__17663),
            .I(delay_counter_3));
    LocalMux I__1547 (
            .O(N__17660),
            .I(delay_counter_3));
    InMux I__1546 (
            .O(N__17655),
            .I(n10584));
    InMux I__1545 (
            .O(N__17652),
            .I(N__17648));
    InMux I__1544 (
            .O(N__17651),
            .I(N__17645));
    LocalMux I__1543 (
            .O(N__17648),
            .I(delay_counter_4));
    LocalMux I__1542 (
            .O(N__17645),
            .I(delay_counter_4));
    InMux I__1541 (
            .O(N__17640),
            .I(n10585));
    InMux I__1540 (
            .O(N__17637),
            .I(N__17633));
    InMux I__1539 (
            .O(N__17636),
            .I(N__17630));
    LocalMux I__1538 (
            .O(N__17633),
            .I(delay_counter_5));
    LocalMux I__1537 (
            .O(N__17630),
            .I(delay_counter_5));
    InMux I__1536 (
            .O(N__17625),
            .I(n10586));
    InMux I__1535 (
            .O(N__17622),
            .I(N__17618));
    InMux I__1534 (
            .O(N__17621),
            .I(N__17615));
    LocalMux I__1533 (
            .O(N__17618),
            .I(delay_counter_6));
    LocalMux I__1532 (
            .O(N__17615),
            .I(delay_counter_6));
    InMux I__1531 (
            .O(N__17610),
            .I(n10587));
    CascadeMux I__1530 (
            .O(N__17607),
            .I(N__17604));
    InMux I__1529 (
            .O(N__17604),
            .I(N__17600));
    InMux I__1528 (
            .O(N__17603),
            .I(N__17597));
    LocalMux I__1527 (
            .O(N__17600),
            .I(N__17594));
    LocalMux I__1526 (
            .O(N__17597),
            .I(delay_counter_7));
    Odrv4 I__1525 (
            .O(N__17594),
            .I(delay_counter_7));
    InMux I__1524 (
            .O(N__17589),
            .I(n10588));
    InMux I__1523 (
            .O(N__17586),
            .I(N__17582));
    InMux I__1522 (
            .O(N__17585),
            .I(N__17579));
    LocalMux I__1521 (
            .O(N__17582),
            .I(N__17576));
    LocalMux I__1520 (
            .O(N__17579),
            .I(delay_counter_8));
    Odrv4 I__1519 (
            .O(N__17576),
            .I(delay_counter_8));
    InMux I__1518 (
            .O(N__17571),
            .I(bfn_1_23_0_));
    InMux I__1517 (
            .O(N__17568),
            .I(N__17564));
    InMux I__1516 (
            .O(N__17567),
            .I(N__17561));
    LocalMux I__1515 (
            .O(N__17564),
            .I(neo_pixel_transmitter_t0_18));
    LocalMux I__1514 (
            .O(N__17561),
            .I(neo_pixel_transmitter_t0_18));
    InMux I__1513 (
            .O(N__17556),
            .I(N__17552));
    InMux I__1512 (
            .O(N__17555),
            .I(N__17549));
    LocalMux I__1511 (
            .O(N__17552),
            .I(neo_pixel_transmitter_t0_20));
    LocalMux I__1510 (
            .O(N__17549),
            .I(neo_pixel_transmitter_t0_20));
    InMux I__1509 (
            .O(N__17544),
            .I(N__17538));
    InMux I__1508 (
            .O(N__17543),
            .I(N__17538));
    LocalMux I__1507 (
            .O(N__17538),
            .I(neo_pixel_transmitter_t0_24));
    InMux I__1506 (
            .O(N__17535),
            .I(N__17529));
    InMux I__1505 (
            .O(N__17534),
            .I(N__17529));
    LocalMux I__1504 (
            .O(N__17529),
            .I(neo_pixel_transmitter_t0_31));
    InMux I__1503 (
            .O(N__17526),
            .I(N__17523));
    LocalMux I__1502 (
            .O(N__17523),
            .I(n15_adj_841));
    InMux I__1501 (
            .O(N__17520),
            .I(N__17517));
    LocalMux I__1500 (
            .O(N__17517),
            .I(n14_adj_842));
    InMux I__1499 (
            .O(N__17514),
            .I(N__17510));
    InMux I__1498 (
            .O(N__17513),
            .I(N__17507));
    LocalMux I__1497 (
            .O(N__17510),
            .I(N__17504));
    LocalMux I__1496 (
            .O(N__17507),
            .I(delay_counter_0));
    Odrv4 I__1495 (
            .O(N__17504),
            .I(delay_counter_0));
    InMux I__1494 (
            .O(N__17499),
            .I(bfn_1_22_0_));
    InMux I__1493 (
            .O(N__17496),
            .I(N__17490));
    InMux I__1492 (
            .O(N__17495),
            .I(N__17490));
    LocalMux I__1491 (
            .O(N__17490),
            .I(neo_pixel_transmitter_t0_9));
    InMux I__1490 (
            .O(N__17487),
            .I(N__17484));
    LocalMux I__1489 (
            .O(N__17484),
            .I(neopxl_color_prev_12));
    CascadeMux I__1488 (
            .O(N__17481),
            .I(n24_adj_801_cascade_));
    InMux I__1487 (
            .O(N__17478),
            .I(N__17475));
    LocalMux I__1486 (
            .O(N__17475),
            .I(n12414));
    InMux I__1485 (
            .O(N__17472),
            .I(N__17469));
    LocalMux I__1484 (
            .O(N__17469),
            .I(N__17466));
    Odrv4 I__1483 (
            .O(N__17466),
            .I(neopxl_color_prev_6));
    InMux I__1482 (
            .O(N__17463),
            .I(N__17457));
    InMux I__1481 (
            .O(N__17462),
            .I(N__17457));
    LocalMux I__1480 (
            .O(N__17457),
            .I(neo_pixel_transmitter_t0_21));
    InMux I__1479 (
            .O(N__17454),
            .I(N__17448));
    InMux I__1478 (
            .O(N__17453),
            .I(N__17448));
    LocalMux I__1477 (
            .O(N__17448),
            .I(neo_pixel_transmitter_t0_7));
    InMux I__1476 (
            .O(N__17445),
            .I(N__17439));
    InMux I__1475 (
            .O(N__17444),
            .I(N__17439));
    LocalMux I__1474 (
            .O(N__17439),
            .I(neo_pixel_transmitter_t0_12));
    InMux I__1473 (
            .O(N__17436),
            .I(N__17430));
    InMux I__1472 (
            .O(N__17435),
            .I(N__17430));
    LocalMux I__1471 (
            .O(N__17430),
            .I(neo_pixel_transmitter_t0_4));
    InMux I__1470 (
            .O(N__17427),
            .I(N__17421));
    InMux I__1469 (
            .O(N__17426),
            .I(N__17421));
    LocalMux I__1468 (
            .O(N__17421),
            .I(neo_pixel_transmitter_t0_0));
    IoInMux I__1467 (
            .O(N__17418),
            .I(N__17415));
    LocalMux I__1466 (
            .O(N__17415),
            .I(N__17412));
    IoSpan4Mux I__1465 (
            .O(N__17412),
            .I(N__17409));
    IoSpan4Mux I__1464 (
            .O(N__17409),
            .I(N__17406));
    IoSpan4Mux I__1463 (
            .O(N__17406),
            .I(N__17403));
    Odrv4 I__1462 (
            .O(N__17403),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_2_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_19_0_));
    defparam IN_MUX_bfv_2_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_20_0_ (
            .carryinitin(\nx.n10676 ),
            .carryinitout(bfn_2_20_0_));
    defparam IN_MUX_bfv_2_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_21_0_ (
            .carryinitin(\nx.n10683_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_2_21_0_));
    defparam IN_MUX_bfv_2_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_22_0_ (
            .carryinitin(\nx.n10689_THRU_CRY_1_THRU_CO ),
            .carryinitout(bfn_2_22_0_));
    defparam IN_MUX_bfv_2_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_23_0_ (
            .carryinitin(\nx.n10695_THRU_CRY_1_THRU_CO ),
            .carryinitout(bfn_2_23_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(\nx.n10714 ),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\nx.n10722 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_3_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_21_0_ (
            .carryinitin(\nx.n10730 ),
            .carryinitout(bfn_3_21_0_));
    defparam IN_MUX_bfv_4_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_23_0_));
    defparam IN_MUX_bfv_4_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_24_0_ (
            .carryinitin(\nx.n10771 ),
            .carryinitout(bfn_4_24_0_));
    defparam IN_MUX_bfv_5_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_22_0_));
    defparam IN_MUX_bfv_5_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_23_0_ (
            .carryinitin(\nx.n10763 ),
            .carryinitout(bfn_5_23_0_));
    defparam IN_MUX_bfv_5_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_21_0_));
    defparam IN_MUX_bfv_6_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_20_0_));
    defparam IN_MUX_bfv_7_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_22_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\nx.n11086 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(\nx.n11094 ),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(\nx.n11102 ),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\nx.n11060 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\nx.n11068 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(\nx.n11076 ),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\nx.n11035 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\nx.n11043 ),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\nx.n11051 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(\nx.n11011 ),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(\nx.n11019 ),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\nx.n11027 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(\nx.n10988 ),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_10_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_25_0_ (
            .carryinitin(\nx.n10996 ),
            .carryinitout(bfn_10_25_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(\nx.n10966 ),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(\nx.n10974 ),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_16_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_25_0_ (
            .carryinitin(\nx.n10945 ),
            .carryinitout(bfn_16_25_0_));
    defparam IN_MUX_bfv_16_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_26_0_ (
            .carryinitin(\nx.n10953 ),
            .carryinitout(bfn_16_26_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(\nx.n10925 ),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(\nx.n10933 ),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_13_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_27_0_ (
            .carryinitin(\nx.n10906 ),
            .carryinitout(bfn_13_27_0_));
    defparam IN_MUX_bfv_13_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_28_0_ (
            .carryinitin(\nx.n10914 ),
            .carryinitout(bfn_13_28_0_));
    defparam IN_MUX_bfv_11_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_25_0_));
    defparam IN_MUX_bfv_11_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_26_0_ (
            .carryinitin(\nx.n10888 ),
            .carryinitout(bfn_11_26_0_));
    defparam IN_MUX_bfv_11_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_27_0_ (
            .carryinitin(\nx.n10896 ),
            .carryinitout(bfn_11_27_0_));
    defparam IN_MUX_bfv_11_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_29_0_));
    defparam IN_MUX_bfv_11_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_30_0_ (
            .carryinitin(\nx.n10871 ),
            .carryinitout(bfn_11_30_0_));
    defparam IN_MUX_bfv_11_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_31_0_ (
            .carryinitin(\nx.n10879 ),
            .carryinitout(bfn_11_31_0_));
    defparam IN_MUX_bfv_9_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_26_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(\nx.n10855 ),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\nx.n10863 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_7_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_27_0_));
    defparam IN_MUX_bfv_7_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_28_0_ (
            .carryinitin(\nx.n10840 ),
            .carryinitout(bfn_7_28_0_));
    defparam IN_MUX_bfv_6_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_27_0_));
    defparam IN_MUX_bfv_6_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_28_0_ (
            .carryinitin(\nx.n10826 ),
            .carryinitout(bfn_6_28_0_));
    defparam IN_MUX_bfv_5_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_27_0_));
    defparam IN_MUX_bfv_5_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_28_0_ (
            .carryinitin(\nx.n10813 ),
            .carryinitout(bfn_5_28_0_));
    defparam IN_MUX_bfv_5_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_25_0_));
    defparam IN_MUX_bfv_5_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_26_0_ (
            .carryinitin(\nx.n10801 ),
            .carryinitout(bfn_5_26_0_));
    defparam IN_MUX_bfv_4_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_26_0_));
    defparam IN_MUX_bfv_4_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_27_0_ (
            .carryinitin(\nx.n10790 ),
            .carryinitout(bfn_4_27_0_));
    defparam IN_MUX_bfv_2_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_25_0_));
    defparam IN_MUX_bfv_2_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_26_0_ (
            .carryinitin(\nx.n10780 ),
            .carryinitout(bfn_2_26_0_));
    defparam IN_MUX_bfv_6_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_23_0_));
    defparam IN_MUX_bfv_6_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_24_0_ (
            .carryinitin(\nx.n10620 ),
            .carryinitout(bfn_6_24_0_));
    defparam IN_MUX_bfv_6_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_25_0_ (
            .carryinitin(\nx.n10628 ),
            .carryinitout(bfn_6_25_0_));
    defparam IN_MUX_bfv_6_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_26_0_ (
            .carryinitin(\nx.n10636 ),
            .carryinitout(bfn_6_26_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_1_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_23_0_ (
            .carryinitin(n10589),
            .carryinitout(bfn_1_23_0_));
    defparam IN_MUX_bfv_1_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_24_0_ (
            .carryinitin(n10597),
            .carryinitout(bfn_1_24_0_));
    defparam IN_MUX_bfv_1_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_25_0_ (
            .carryinitin(n10605),
            .carryinitout(bfn_1_25_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_9_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_29_0_));
    defparam IN_MUX_bfv_9_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_30_0_ (
            .carryinitin(n10651),
            .carryinitout(bfn_9_30_0_));
    defparam IN_MUX_bfv_9_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_31_0_ (
            .carryinitin(n10659),
            .carryinitout(bfn_9_31_0_));
    defparam IN_MUX_bfv_9_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_32_0_ (
            .carryinitin(n10667),
            .carryinitout(bfn_9_32_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_17_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__17418),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i0_LC_1_17_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i0_LC_1_17_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i0_LC_1_17_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i0_LC_1_17_0  (
            .in0(N__18624),
            .in1(N__17427),
            .in2(_gnd_net_),
            .in3(N__25224),
            .lcout(neo_pixel_transmitter_t0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46839),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i22_1_lut_LC_1_17_1 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i22_1_lut_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i22_1_lut_LC_1_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i22_1_lut_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17462),
            .lcout(\nx.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i1_1_lut_LC_1_17_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i1_1_lut_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i1_1_lut_LC_1_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i1_1_lut_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17426),
            .lcout(\nx.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i21_LC_1_17_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i21_LC_1_17_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i21_LC_1_17_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i21_LC_1_17_7  (
            .in0(N__25225),
            .in1(N__18906),
            .in2(_gnd_net_),
            .in3(N__17463),
            .lcout(neo_pixel_transmitter_t0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46839),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i12_LC_1_18_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i12_LC_1_18_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i12_LC_1_18_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i12_LC_1_18_0  (
            .in0(N__25230),
            .in1(N__18714),
            .in2(_gnd_net_),
            .in3(N__17445),
            .lcout(neo_pixel_transmitter_t0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46841),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i8_1_lut_LC_1_18_2 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i8_1_lut_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i8_1_lut_LC_1_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i8_1_lut_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17453),
            .lcout(\nx.n26_adj_722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i5_1_lut_LC_1_18_3 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i5_1_lut_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i5_1_lut_LC_1_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i5_1_lut_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17435),
            .lcout(\nx.n29_adj_714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i7_LC_1_18_4 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i7_LC_1_18_4 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i7_LC_1_18_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i7_LC_1_18_4  (
            .in0(N__25232),
            .in1(N__18510),
            .in2(_gnd_net_),
            .in3(N__17454),
            .lcout(neo_pixel_transmitter_t0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46841),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i7_1_lut_LC_1_18_5 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i7_1_lut_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i7_1_lut_LC_1_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i7_1_lut_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17945),
            .lcout(\nx.n27_adj_720 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i13_1_lut_LC_1_18_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i13_1_lut_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i13_1_lut_LC_1_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i13_1_lut_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17444),
            .lcout(\nx.n21_adj_737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i4_LC_1_18_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i4_LC_1_18_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i4_LC_1_18_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i4_LC_1_18_7  (
            .in0(N__18564),
            .in1(N__17436),
            .in2(_gnd_net_),
            .in3(N__25231),
            .lcout(neo_pixel_transmitter_t0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46841),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i20_LC_1_19_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i20_LC_1_19_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i20_LC_1_19_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i20_LC_1_19_0  (
            .in0(N__25234),
            .in1(N__18933),
            .in2(_gnd_net_),
            .in3(N__17556),
            .lcout(neo_pixel_transmitter_t0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46843),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i9_LC_1_19_1 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i9_LC_1_19_1 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i9_LC_1_19_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i9_LC_1_19_1  (
            .in0(N__17496),
            .in1(N__18768),
            .in2(_gnd_net_),
            .in3(N__25235),
            .lcout(neo_pixel_transmitter_t0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46843),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_169_LC_1_19_3.C_ON=1'b0;
    defparam i4_4_lut_adj_169_LC_1_19_3.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_169_LC_1_19_3.LUT_INIT=16'b0111101111011110;
    LogicCell40 i4_4_lut_adj_169_LC_1_19_3 (
            .in0(N__17472),
            .in1(N__26606),
            .in2(N__26220),
            .in3(N__17487),
            .lcout(n12_adj_844),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i10_1_lut_LC_1_19_4 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i10_1_lut_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i10_1_lut_LC_1_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i10_1_lut_LC_1_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17495),
            .lcout(\nx.n24_adj_734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i12_LC_1_19_5.C_ON=1'b0;
    defparam neopxl_color_prev_i12_LC_1_19_5.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i12_LC_1_19_5.LUT_INIT=16'b1100110011001100;
    LogicCell40 neopxl_color_prev_i12_LC_1_19_5 (
            .in0(_gnd_net_),
            .in1(N__26607),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(neopxl_color_prev_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46843),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i30_1_lut_LC_1_19_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i30_1_lut_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i30_1_lut_LC_1_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i30_1_lut_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20157),
            .lcout(\nx.n4_adj_710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i18_LC_1_19_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i18_LC_1_19_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i18_LC_1_19_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i18_LC_1_19_7  (
            .in0(N__18966),
            .in1(N__17568),
            .in2(_gnd_net_),
            .in3(N__25233),
            .lcout(neo_pixel_transmitter_t0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46843),
            .ce(),
            .sr(_gnd_net_));
    defparam i820_4_lut_LC_1_20_0.C_ON=1'b0;
    defparam i820_4_lut_LC_1_20_0.SEQ_MODE=4'b0000;
    defparam i820_4_lut_LC_1_20_0.LUT_INIT=16'b1100100010001000;
    LogicCell40 i820_4_lut_LC_1_20_0 (
            .in0(N__17799),
            .in1(N__17781),
            .in2(N__17820),
            .in3(N__17478),
            .lcout(),
            .ltout(n24_adj_801_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_1_20_1.C_ON=1'b0;
    defparam i2_4_lut_LC_1_20_1.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_1_20_1.LUT_INIT=16'b1010100000000000;
    LogicCell40 i2_4_lut_LC_1_20_1 (
            .in0(N__17745),
            .in1(N__17763),
            .in2(N__17481),
            .in3(N__17727),
            .lcout(n12382),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_LC_1_20_3.C_ON=1'b0;
    defparam i8_4_lut_LC_1_20_3.SEQ_MODE=4'b0000;
    defparam i8_4_lut_LC_1_20_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i8_4_lut_LC_1_20_3 (
            .in0(N__17514),
            .in1(N__17520),
            .in2(N__17607),
            .in3(N__17526),
            .lcout(n12414),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i6_LC_1_20_4.C_ON=1'b0;
    defparam neopxl_color_prev_i6_LC_1_20_4.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i6_LC_1_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 neopxl_color_prev_i6_LC_1_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26219),
            .lcout(neopxl_color_prev_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46845),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i19_1_lut_LC_1_20_5 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i19_1_lut_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i19_1_lut_LC_1_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i19_1_lut_LC_1_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17567),
            .lcout(\nx.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i21_1_lut_LC_1_20_7 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i21_1_lut_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i21_1_lut_LC_1_20_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \nx.sub_14_inv_0_i21_1_lut_LC_1_20_7  (
            .in0(_gnd_net_),
            .in1(N__17555),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\nx.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i31_LC_1_21_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i31_LC_1_21_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i31_LC_1_21_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i31_LC_1_21_0  (
            .in0(N__19047),
            .in1(N__17535),
            .in2(_gnd_net_),
            .in3(N__25237),
            .lcout(neo_pixel_transmitter_t0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46848),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i24_LC_1_21_1 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i24_LC_1_21_1 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i24_LC_1_21_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i24_LC_1_21_1  (
            .in0(N__25236),
            .in1(N__18819),
            .in2(_gnd_net_),
            .in3(N__17544),
            .lcout(neo_pixel_transmitter_t0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46848),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_1_21_2.C_ON=1'b0;
    defparam i7_4_lut_LC_1_21_2.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_1_21_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i7_4_lut_LC_1_21_2 (
            .in0(N__17841),
            .in1(N__17925),
            .in2(N__17865),
            .in3(N__17901),
            .lcout(n18_adj_815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i25_1_lut_LC_1_21_3 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i25_1_lut_LC_1_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i25_1_lut_LC_1_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i25_1_lut_LC_1_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17543),
            .lcout(\nx.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i32_1_lut_LC_1_21_4 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i32_1_lut_LC_1_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i32_1_lut_LC_1_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i32_1_lut_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17534),
            .lcout(\nx.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_1_21_5.C_ON=1'b0;
    defparam i6_4_lut_LC_1_21_5.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_1_21_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_LC_1_21_5 (
            .in0(N__17699),
            .in1(N__17621),
            .in2(N__17685),
            .in3(N__17586),
            .lcout(n15_adj_841),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_3_lut_LC_1_21_6.C_ON=1'b0;
    defparam i5_3_lut_LC_1_21_6.SEQ_MODE=4'b0000;
    defparam i5_3_lut_LC_1_21_6.LUT_INIT=16'b1111111111101110;
    LogicCell40 i5_3_lut_LC_1_21_6 (
            .in0(N__17651),
            .in1(N__17636),
            .in2(_gnd_net_),
            .in3(N__17666),
            .lcout(n14_adj_842),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_counter_634__i0_LC_1_22_0.C_ON=1'b1;
    defparam delay_counter_634__i0_LC_1_22_0.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i0_LC_1_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i0_LC_1_22_0 (
            .in0(_gnd_net_),
            .in1(N__17513),
            .in2(_gnd_net_),
            .in3(N__17499),
            .lcout(delay_counter_0),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(n10582),
            .clk(N__46852),
            .ce(N__22314),
            .sr(N__43506));
    defparam delay_counter_634__i1_LC_1_22_1.C_ON=1'b1;
    defparam delay_counter_634__i1_LC_1_22_1.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i1_LC_1_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i1_LC_1_22_1 (
            .in0(_gnd_net_),
            .in1(N__17700),
            .in2(_gnd_net_),
            .in3(N__17688),
            .lcout(delay_counter_1),
            .ltout(),
            .carryin(n10582),
            .carryout(n10583),
            .clk(N__46852),
            .ce(N__22314),
            .sr(N__43506));
    defparam delay_counter_634__i2_LC_1_22_2.C_ON=1'b1;
    defparam delay_counter_634__i2_LC_1_22_2.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i2_LC_1_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i2_LC_1_22_2 (
            .in0(_gnd_net_),
            .in1(N__17684),
            .in2(_gnd_net_),
            .in3(N__17670),
            .lcout(delay_counter_2),
            .ltout(),
            .carryin(n10583),
            .carryout(n10584),
            .clk(N__46852),
            .ce(N__22314),
            .sr(N__43506));
    defparam delay_counter_634__i3_LC_1_22_3.C_ON=1'b1;
    defparam delay_counter_634__i3_LC_1_22_3.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i3_LC_1_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i3_LC_1_22_3 (
            .in0(_gnd_net_),
            .in1(N__17667),
            .in2(_gnd_net_),
            .in3(N__17655),
            .lcout(delay_counter_3),
            .ltout(),
            .carryin(n10584),
            .carryout(n10585),
            .clk(N__46852),
            .ce(N__22314),
            .sr(N__43506));
    defparam delay_counter_634__i4_LC_1_22_4.C_ON=1'b1;
    defparam delay_counter_634__i4_LC_1_22_4.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i4_LC_1_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i4_LC_1_22_4 (
            .in0(_gnd_net_),
            .in1(N__17652),
            .in2(_gnd_net_),
            .in3(N__17640),
            .lcout(delay_counter_4),
            .ltout(),
            .carryin(n10585),
            .carryout(n10586),
            .clk(N__46852),
            .ce(N__22314),
            .sr(N__43506));
    defparam delay_counter_634__i5_LC_1_22_5.C_ON=1'b1;
    defparam delay_counter_634__i5_LC_1_22_5.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i5_LC_1_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i5_LC_1_22_5 (
            .in0(_gnd_net_),
            .in1(N__17637),
            .in2(_gnd_net_),
            .in3(N__17625),
            .lcout(delay_counter_5),
            .ltout(),
            .carryin(n10586),
            .carryout(n10587),
            .clk(N__46852),
            .ce(N__22314),
            .sr(N__43506));
    defparam delay_counter_634__i6_LC_1_22_6.C_ON=1'b1;
    defparam delay_counter_634__i6_LC_1_22_6.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i6_LC_1_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i6_LC_1_22_6 (
            .in0(_gnd_net_),
            .in1(N__17622),
            .in2(_gnd_net_),
            .in3(N__17610),
            .lcout(delay_counter_6),
            .ltout(),
            .carryin(n10587),
            .carryout(n10588),
            .clk(N__46852),
            .ce(N__22314),
            .sr(N__43506));
    defparam delay_counter_634__i7_LC_1_22_7.C_ON=1'b1;
    defparam delay_counter_634__i7_LC_1_22_7.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i7_LC_1_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i7_LC_1_22_7 (
            .in0(_gnd_net_),
            .in1(N__17603),
            .in2(_gnd_net_),
            .in3(N__17589),
            .lcout(delay_counter_7),
            .ltout(),
            .carryin(n10588),
            .carryout(n10589),
            .clk(N__46852),
            .ce(N__22314),
            .sr(N__43506));
    defparam delay_counter_634__i8_LC_1_23_0.C_ON=1'b1;
    defparam delay_counter_634__i8_LC_1_23_0.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i8_LC_1_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i8_LC_1_23_0 (
            .in0(_gnd_net_),
            .in1(N__17585),
            .in2(_gnd_net_),
            .in3(N__17571),
            .lcout(delay_counter_8),
            .ltout(),
            .carryin(bfn_1_23_0_),
            .carryout(n10590),
            .clk(N__46858),
            .ce(N__22303),
            .sr(N__43491));
    defparam delay_counter_634__i9_LC_1_23_1.C_ON=1'b1;
    defparam delay_counter_634__i9_LC_1_23_1.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i9_LC_1_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i9_LC_1_23_1 (
            .in0(_gnd_net_),
            .in1(N__17816),
            .in2(_gnd_net_),
            .in3(N__17802),
            .lcout(delay_counter_9),
            .ltout(),
            .carryin(n10590),
            .carryout(n10591),
            .clk(N__46858),
            .ce(N__22303),
            .sr(N__43491));
    defparam delay_counter_634__i10_LC_1_23_2.C_ON=1'b1;
    defparam delay_counter_634__i10_LC_1_23_2.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i10_LC_1_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i10_LC_1_23_2 (
            .in0(_gnd_net_),
            .in1(N__17798),
            .in2(_gnd_net_),
            .in3(N__17784),
            .lcout(delay_counter_10),
            .ltout(),
            .carryin(n10591),
            .carryout(n10592),
            .clk(N__46858),
            .ce(N__22303),
            .sr(N__43491));
    defparam delay_counter_634__i11_LC_1_23_3.C_ON=1'b1;
    defparam delay_counter_634__i11_LC_1_23_3.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i11_LC_1_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i11_LC_1_23_3 (
            .in0(_gnd_net_),
            .in1(N__17780),
            .in2(_gnd_net_),
            .in3(N__17766),
            .lcout(delay_counter_11),
            .ltout(),
            .carryin(n10592),
            .carryout(n10593),
            .clk(N__46858),
            .ce(N__22303),
            .sr(N__43491));
    defparam delay_counter_634__i12_LC_1_23_4.C_ON=1'b1;
    defparam delay_counter_634__i12_LC_1_23_4.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i12_LC_1_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i12_LC_1_23_4 (
            .in0(_gnd_net_),
            .in1(N__17762),
            .in2(_gnd_net_),
            .in3(N__17748),
            .lcout(delay_counter_12),
            .ltout(),
            .carryin(n10593),
            .carryout(n10594),
            .clk(N__46858),
            .ce(N__22303),
            .sr(N__43491));
    defparam delay_counter_634__i13_LC_1_23_5.C_ON=1'b1;
    defparam delay_counter_634__i13_LC_1_23_5.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i13_LC_1_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i13_LC_1_23_5 (
            .in0(_gnd_net_),
            .in1(N__17744),
            .in2(_gnd_net_),
            .in3(N__17730),
            .lcout(delay_counter_13),
            .ltout(),
            .carryin(n10594),
            .carryout(n10595),
            .clk(N__46858),
            .ce(N__22303),
            .sr(N__43491));
    defparam delay_counter_634__i14_LC_1_23_6.C_ON=1'b1;
    defparam delay_counter_634__i14_LC_1_23_6.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i14_LC_1_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i14_LC_1_23_6 (
            .in0(_gnd_net_),
            .in1(N__17726),
            .in2(_gnd_net_),
            .in3(N__17712),
            .lcout(delay_counter_14),
            .ltout(),
            .carryin(n10595),
            .carryout(n10596),
            .clk(N__46858),
            .ce(N__22303),
            .sr(N__43491));
    defparam delay_counter_634__i15_LC_1_23_7.C_ON=1'b1;
    defparam delay_counter_634__i15_LC_1_23_7.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i15_LC_1_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i15_LC_1_23_7 (
            .in0(_gnd_net_),
            .in1(N__19196),
            .in2(_gnd_net_),
            .in3(N__17709),
            .lcout(delay_counter_15),
            .ltout(),
            .carryin(n10596),
            .carryout(n10597),
            .clk(N__46858),
            .ce(N__22303),
            .sr(N__43491));
    defparam delay_counter_634__i16_LC_1_24_0.C_ON=1'b1;
    defparam delay_counter_634__i16_LC_1_24_0.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i16_LC_1_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i16_LC_1_24_0 (
            .in0(_gnd_net_),
            .in1(N__20597),
            .in2(_gnd_net_),
            .in3(N__17706),
            .lcout(delay_counter_16),
            .ltout(),
            .carryin(bfn_1_24_0_),
            .carryout(n10598),
            .clk(N__46863),
            .ce(N__22302),
            .sr(N__43505));
    defparam delay_counter_634__i17_LC_1_24_1.C_ON=1'b1;
    defparam delay_counter_634__i17_LC_1_24_1.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i17_LC_1_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i17_LC_1_24_1 (
            .in0(_gnd_net_),
            .in1(N__19217),
            .in2(_gnd_net_),
            .in3(N__17703),
            .lcout(delay_counter_17),
            .ltout(),
            .carryin(n10598),
            .carryout(n10599),
            .clk(N__46863),
            .ce(N__22302),
            .sr(N__43505));
    defparam delay_counter_634__i18_LC_1_24_2.C_ON=1'b1;
    defparam delay_counter_634__i18_LC_1_24_2.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i18_LC_1_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i18_LC_1_24_2 (
            .in0(_gnd_net_),
            .in1(N__20612),
            .in2(_gnd_net_),
            .in3(N__17880),
            .lcout(delay_counter_18),
            .ltout(),
            .carryin(n10599),
            .carryout(n10600),
            .clk(N__46863),
            .ce(N__22302),
            .sr(N__43505));
    defparam delay_counter_634__i19_LC_1_24_3.C_ON=1'b1;
    defparam delay_counter_634__i19_LC_1_24_3.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i19_LC_1_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i19_LC_1_24_3 (
            .in0(_gnd_net_),
            .in1(N__22040),
            .in2(_gnd_net_),
            .in3(N__17877),
            .lcout(delay_counter_19),
            .ltout(),
            .carryin(n10600),
            .carryout(n10601),
            .clk(N__46863),
            .ce(N__22302),
            .sr(N__43505));
    defparam delay_counter_634__i20_LC_1_24_4.C_ON=1'b1;
    defparam delay_counter_634__i20_LC_1_24_4.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i20_LC_1_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i20_LC_1_24_4 (
            .in0(_gnd_net_),
            .in1(N__22022),
            .in2(_gnd_net_),
            .in3(N__17874),
            .lcout(delay_counter_20),
            .ltout(),
            .carryin(n10601),
            .carryout(n10602),
            .clk(N__46863),
            .ce(N__22302),
            .sr(N__43505));
    defparam delay_counter_634__i21_LC_1_24_5.C_ON=1'b1;
    defparam delay_counter_634__i21_LC_1_24_5.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i21_LC_1_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i21_LC_1_24_5 (
            .in0(_gnd_net_),
            .in1(N__19298),
            .in2(_gnd_net_),
            .in3(N__17871),
            .lcout(delay_counter_21),
            .ltout(),
            .carryin(n10602),
            .carryout(n10603),
            .clk(N__46863),
            .ce(N__22302),
            .sr(N__43505));
    defparam delay_counter_634__i22_LC_1_24_6.C_ON=1'b1;
    defparam delay_counter_634__i22_LC_1_24_6.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i22_LC_1_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i22_LC_1_24_6 (
            .in0(_gnd_net_),
            .in1(N__20756),
            .in2(_gnd_net_),
            .in3(N__17868),
            .lcout(delay_counter_22),
            .ltout(),
            .carryin(n10603),
            .carryout(n10604),
            .clk(N__46863),
            .ce(N__22302),
            .sr(N__43505));
    defparam delay_counter_634__i23_LC_1_24_7.C_ON=1'b1;
    defparam delay_counter_634__i23_LC_1_24_7.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i23_LC_1_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i23_LC_1_24_7 (
            .in0(_gnd_net_),
            .in1(N__17861),
            .in2(_gnd_net_),
            .in3(N__17847),
            .lcout(delay_counter_23),
            .ltout(),
            .carryin(n10604),
            .carryout(n10605),
            .clk(N__46863),
            .ce(N__22302),
            .sr(N__43505));
    defparam delay_counter_634__i24_LC_1_25_0.C_ON=1'b1;
    defparam delay_counter_634__i24_LC_1_25_0.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i24_LC_1_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i24_LC_1_25_0 (
            .in0(_gnd_net_),
            .in1(N__20777),
            .in2(_gnd_net_),
            .in3(N__17844),
            .lcout(delay_counter_24),
            .ltout(),
            .carryin(bfn_1_25_0_),
            .carryout(n10606),
            .clk(N__46870),
            .ce(N__22310),
            .sr(N__43492));
    defparam delay_counter_634__i25_LC_1_25_1.C_ON=1'b1;
    defparam delay_counter_634__i25_LC_1_25_1.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i25_LC_1_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i25_LC_1_25_1 (
            .in0(_gnd_net_),
            .in1(N__17840),
            .in2(_gnd_net_),
            .in3(N__17826),
            .lcout(delay_counter_25),
            .ltout(),
            .carryin(n10606),
            .carryout(n10607),
            .clk(N__46870),
            .ce(N__22310),
            .sr(N__43492));
    defparam delay_counter_634__i26_LC_1_25_2.C_ON=1'b1;
    defparam delay_counter_634__i26_LC_1_25_2.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i26_LC_1_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i26_LC_1_25_2 (
            .in0(_gnd_net_),
            .in1(N__20741),
            .in2(_gnd_net_),
            .in3(N__17823),
            .lcout(delay_counter_26),
            .ltout(),
            .carryin(n10607),
            .carryout(n10608),
            .clk(N__46870),
            .ce(N__22310),
            .sr(N__43492));
    defparam delay_counter_634__i27_LC_1_25_3.C_ON=1'b1;
    defparam delay_counter_634__i27_LC_1_25_3.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i27_LC_1_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i27_LC_1_25_3 (
            .in0(_gnd_net_),
            .in1(N__17924),
            .in2(_gnd_net_),
            .in3(N__17910),
            .lcout(delay_counter_27),
            .ltout(),
            .carryin(n10608),
            .carryout(n10609),
            .clk(N__46870),
            .ce(N__22310),
            .sr(N__43492));
    defparam delay_counter_634__i28_LC_1_25_4.C_ON=1'b1;
    defparam delay_counter_634__i28_LC_1_25_4.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i28_LC_1_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i28_LC_1_25_4 (
            .in0(_gnd_net_),
            .in1(N__20792),
            .in2(_gnd_net_),
            .in3(N__17907),
            .lcout(delay_counter_28),
            .ltout(),
            .carryin(n10609),
            .carryout(n10610),
            .clk(N__46870),
            .ce(N__22310),
            .sr(N__43492));
    defparam delay_counter_634__i29_LC_1_25_5.C_ON=1'b1;
    defparam delay_counter_634__i29_LC_1_25_5.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i29_LC_1_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i29_LC_1_25_5 (
            .in0(_gnd_net_),
            .in1(N__19277),
            .in2(_gnd_net_),
            .in3(N__17904),
            .lcout(delay_counter_29),
            .ltout(),
            .carryin(n10610),
            .carryout(n10611),
            .clk(N__46870),
            .ce(N__22310),
            .sr(N__43492));
    defparam delay_counter_634__i30_LC_1_25_6.C_ON=1'b1;
    defparam delay_counter_634__i30_LC_1_25_6.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i30_LC_1_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i30_LC_1_25_6 (
            .in0(_gnd_net_),
            .in1(N__17900),
            .in2(_gnd_net_),
            .in3(N__17886),
            .lcout(delay_counter_30),
            .ltout(),
            .carryin(n10611),
            .carryout(n10612),
            .clk(N__46870),
            .ce(N__22310),
            .sr(N__43492));
    defparam delay_counter_634__i31_LC_1_25_7.C_ON=1'b0;
    defparam delay_counter_634__i31_LC_1_25_7.SEQ_MODE=4'b1000;
    defparam delay_counter_634__i31_LC_1_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_634__i31_LC_1_25_7 (
            .in0(_gnd_net_),
            .in1(N__23711),
            .in2(_gnd_net_),
            .in3(N__17883),
            .lcout(delay_counter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46870),
            .ce(N__22310),
            .sr(N__43492));
    defparam \nx.sub_14_inv_0_i9_1_lut_LC_2_17_0 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i9_1_lut_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i9_1_lut_LC_2_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i9_1_lut_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17963),
            .lcout(\nx.n25_adj_724 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i3_1_lut_LC_2_17_1 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i3_1_lut_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i3_1_lut_LC_2_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i3_1_lut_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17954),
            .lcout(\nx.n31_adj_711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i15_LC_2_17_2 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i15_LC_2_17_2 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i15_LC_2_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i15_LC_2_17_2  (
            .in0(N__17973),
            .in1(N__18654),
            .in2(_gnd_net_),
            .in3(N__25176),
            .lcout(neo_pixel_transmitter_t0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46840),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i24_1_lut_LC_2_17_3 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i24_1_lut_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i24_1_lut_LC_2_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i24_1_lut_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17981),
            .lcout(\nx.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_4 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_4 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_4  (
            .in0(N__17982),
            .in1(N__18846),
            .in2(_gnd_net_),
            .in3(N__25177),
            .lcout(neo_pixel_transmitter_t0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46840),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i16_1_lut_LC_2_17_5 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i16_1_lut_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i16_1_lut_LC_2_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i16_1_lut_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17972),
            .lcout(\nx.n18_adj_723 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i8_LC_2_17_6 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i8_LC_2_17_6 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i8_LC_2_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i8_LC_2_17_6  (
            .in0(N__18792),
            .in1(N__17964),
            .in2(_gnd_net_),
            .in3(N__25179),
            .lcout(neo_pixel_transmitter_t0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46840),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i2_LC_2_17_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i2_LC_2_17_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i2_LC_2_17_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i2_LC_2_17_7  (
            .in0(N__25178),
            .in1(N__18590),
            .in2(_gnd_net_),
            .in3(N__17955),
            .lcout(neo_pixel_transmitter_t0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46840),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_18_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_18_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_18_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_18_0  (
            .in0(N__25229),
            .in1(N__18533),
            .in2(_gnd_net_),
            .in3(N__17946),
            .lcout(neo_pixel_transmitter_t0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46844),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i23_1_lut_LC_2_18_1 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i23_1_lut_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i23_1_lut_LC_2_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i23_1_lut_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18047),
            .lcout(\nx.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i17_LC_2_18_2 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i17_LC_2_18_2 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i17_LC_2_18_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i17_LC_2_18_2  (
            .in0(N__25227),
            .in1(N__18993),
            .in2(_gnd_net_),
            .in3(N__17934),
            .lcout(neo_pixel_transmitter_t0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46844),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i10_LC_2_18_3 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i10_LC_2_18_3 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i10_LC_2_18_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i10_LC_2_18_3  (
            .in0(N__18744),
            .in1(N__18039),
            .in2(_gnd_net_),
            .in3(N__25226),
            .lcout(neo_pixel_transmitter_t0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46844),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i18_1_lut_LC_2_18_4 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i18_1_lut_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i18_1_lut_LC_2_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i18_1_lut_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17933),
            .lcout(\nx.n16_adj_672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i22_LC_2_18_5 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i22_LC_2_18_5 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i22_LC_2_18_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i22_LC_2_18_5  (
            .in0(N__18876),
            .in1(N__18048),
            .in2(_gnd_net_),
            .in3(N__25228),
            .lcout(neo_pixel_transmitter_t0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46844),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i11_1_lut_LC_2_18_7 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i11_1_lut_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i11_1_lut_LC_2_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i11_1_lut_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18038),
            .lcout(\nx.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_2_LC_2_19_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_2_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_2_LC_2_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_2_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__18030),
            .in2(N__18620),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_19_0_),
            .carryout(\nx.n10669 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_3_lut_LC_2_19_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_3_lut_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_3_lut_LC_2_19_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \nx.sub_14_add_2_3_lut_LC_2_19_1  (
            .in0(N__21375),
            .in1(N__19803),
            .in2(N__19743),
            .in3(N__18021),
            .lcout(\nx.n4_adj_771 ),
            .ltout(),
            .carryin(\nx.n10669 ),
            .carryout(\nx.n10670 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_4_lut_LC_2_19_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_4_lut_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_4_lut_LC_2_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_4_lut_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(N__18018),
            .in2(N__18591),
            .in3(N__18009),
            .lcout(\nx.one_wire_N_599_2 ),
            .ltout(),
            .carryin(\nx.n10670 ),
            .carryout(\nx.n10671 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_5_lut_LC_2_19_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_5_lut_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_5_lut_LC_2_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_5_lut_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(N__19815),
            .in2(N__19710),
            .in3(N__18006),
            .lcout(\nx.one_wire_N_599_3 ),
            .ltout(),
            .carryin(\nx.n10671 ),
            .carryout(\nx.n10672 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_6_lut_LC_2_19_4 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_6_lut_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_6_lut_LC_2_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_6_lut_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__18003),
            .in2(N__18563),
            .in3(N__17997),
            .lcout(\nx.one_wire_N_599_4 ),
            .ltout(),
            .carryin(\nx.n10672 ),
            .carryout(\nx.n10673 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_7_lut_LC_2_19_5 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_7_lut_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_7_lut_LC_2_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_7_lut_LC_2_19_5  (
            .in0(_gnd_net_),
            .in1(N__19771),
            .in2(N__19791),
            .in3(N__17994),
            .lcout(\nx.one_wire_N_599_5 ),
            .ltout(),
            .carryin(\nx.n10673 ),
            .carryout(\nx.n10674 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_8_lut_LC_2_19_6 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_8_lut_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_8_lut_LC_2_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_8_lut_LC_2_19_6  (
            .in0(_gnd_net_),
            .in1(N__17991),
            .in2(N__18534),
            .in3(N__17985),
            .lcout(\nx.one_wire_N_599_6 ),
            .ltout(),
            .carryin(\nx.n10674 ),
            .carryout(\nx.n10675 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_9_lut_LC_2_19_7 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_9_lut_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_9_lut_LC_2_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_9_lut_LC_2_19_7  (
            .in0(_gnd_net_),
            .in1(N__18138),
            .in2(N__18509),
            .in3(N__18132),
            .lcout(\nx.one_wire_N_599_7 ),
            .ltout(),
            .carryin(\nx.n10675 ),
            .carryout(\nx.n10676 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_10_lut_LC_2_20_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_10_lut_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_10_lut_LC_2_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_10_lut_LC_2_20_0  (
            .in0(_gnd_net_),
            .in1(N__18787),
            .in2(N__18129),
            .in3(N__18117),
            .lcout(\nx.one_wire_N_599_8 ),
            .ltout(),
            .carryin(bfn_2_20_0_),
            .carryout(\nx.n10677 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_11_lut_LC_2_20_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_11_lut_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_11_lut_LC_2_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_11_lut_LC_2_20_1  (
            .in0(_gnd_net_),
            .in1(N__18763),
            .in2(N__18114),
            .in3(N__18105),
            .lcout(\nx.one_wire_N_599_9 ),
            .ltout(),
            .carryin(\nx.n10677 ),
            .carryout(\nx.n10678 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_12_lut_LC_2_20_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_12_lut_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_12_lut_LC_2_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_12_lut_LC_2_20_2  (
            .in0(_gnd_net_),
            .in1(N__18102),
            .in2(N__18743),
            .in3(N__18093),
            .lcout(\nx.one_wire_N_599_10 ),
            .ltout(),
            .carryin(\nx.n10678 ),
            .carryout(\nx.n10679 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_13_lut_LC_2_20_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_13_lut_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_13_lut_LC_2_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.sub_14_add_2_13_lut_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(N__21426),
            .in2(N__21560),
            .in3(N__18090),
            .lcout(\nx.one_wire_N_599_11 ),
            .ltout(),
            .carryin(\nx.n10679 ),
            .carryout(\nx.n10680 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_14_lut_LC_2_20_4 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_14_lut_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_14_lut_LC_2_20_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_14_lut_LC_2_20_4  (
            .in0(N__18087),
            .in1(N__18081),
            .in2(N__18710),
            .in3(N__18069),
            .lcout(\nx.n13173 ),
            .ltout(),
            .carryin(\nx.n10680 ),
            .carryout(\nx.n10681 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_15_lut_LC_2_20_5 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_15_lut_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_15_lut_LC_2_20_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_15_lut_LC_2_20_5  (
            .in0(N__18066),
            .in1(N__19944),
            .in2(N__19932),
            .in3(N__18060),
            .lcout(\nx.n13175 ),
            .ltout(),
            .carryin(\nx.n10681 ),
            .carryout(\nx.n10682 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_16_lut_LC_2_20_6 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_16_lut_LC_2_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_16_lut_LC_2_20_6 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_16_lut_LC_2_20_6  (
            .in0(N__18057),
            .in1(N__18459),
            .in2(N__18680),
            .in3(N__18051),
            .lcout(\nx.n13177 ),
            .ltout(),
            .carryin(\nx.n10682 ),
            .carryout(\nx.n10683 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_16_THRU_CRY_0_LC_2_20_7 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_16_THRU_CRY_0_LC_2_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_16_THRU_CRY_0_LC_2_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_16_THRU_CRY_0_LC_2_20_7  (
            .in0(_gnd_net_),
            .in1(N__42223),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10683 ),
            .carryout(\nx.n10683_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_17_lut_LC_2_21_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_17_lut_LC_2_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_17_lut_LC_2_21_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_17_lut_LC_2_21_0  (
            .in0(N__18234),
            .in1(N__18650),
            .in2(N__18228),
            .in3(N__18216),
            .lcout(\nx.n13179 ),
            .ltout(),
            .carryin(bfn_2_21_0_),
            .carryout(\nx.n10684 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_18_lut_LC_2_21_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_18_lut_LC_2_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_18_lut_LC_2_21_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_18_lut_LC_2_21_1  (
            .in0(N__18213),
            .in1(N__19138),
            .in2(N__19110),
            .in3(N__18207),
            .lcout(\nx.n13181 ),
            .ltout(),
            .carryin(\nx.n10684 ),
            .carryout(\nx.n10685 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_19_lut_LC_2_21_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_19_lut_LC_2_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_19_lut_LC_2_21_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_19_lut_LC_2_21_2  (
            .in0(N__18204),
            .in1(N__18198),
            .in2(N__18992),
            .in3(N__18189),
            .lcout(\nx.n13183 ),
            .ltout(),
            .carryin(\nx.n10685 ),
            .carryout(\nx.n10686 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_20_lut_LC_2_21_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_20_lut_LC_2_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_20_lut_LC_2_21_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_20_lut_LC_2_21_3  (
            .in0(N__18186),
            .in1(N__18177),
            .in2(N__18965),
            .in3(N__18171),
            .lcout(\nx.n13185 ),
            .ltout(),
            .carryin(\nx.n10686 ),
            .carryout(\nx.n10687 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_21_lut_LC_2_21_4 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_21_lut_LC_2_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_21_lut_LC_2_21_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_21_lut_LC_2_21_4  (
            .in0(N__18168),
            .in1(N__21402),
            .in2(N__19881),
            .in3(N__18162),
            .lcout(\nx.n13187 ),
            .ltout(),
            .carryin(\nx.n10687 ),
            .carryout(\nx.n10688 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_22_lut_LC_2_21_5 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_22_lut_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_22_lut_LC_2_21_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_22_lut_LC_2_21_5  (
            .in0(N__18159),
            .in1(N__18925),
            .in2(N__18150),
            .in3(N__18141),
            .lcout(\nx.n13189 ),
            .ltout(),
            .carryin(\nx.n10688 ),
            .carryout(\nx.n10689 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_22_THRU_CRY_0_LC_2_21_6 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_22_THRU_CRY_0_LC_2_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_22_THRU_CRY_0_LC_2_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_22_THRU_CRY_0_LC_2_21_6  (
            .in0(_gnd_net_),
            .in1(N__42225),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10689 ),
            .carryout(\nx.n10689_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_22_THRU_CRY_1_LC_2_21_7 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_22_THRU_CRY_1_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_22_THRU_CRY_1_LC_2_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_22_THRU_CRY_1_LC_2_21_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__42281),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10689_THRU_CRY_0_THRU_CO ),
            .carryout(\nx.n10689_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_23_lut_LC_2_22_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_23_lut_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_23_lut_LC_2_22_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_23_lut_LC_2_22_0  (
            .in0(N__18339),
            .in1(N__18902),
            .in2(N__18333),
            .in3(N__18318),
            .lcout(\nx.n13191 ),
            .ltout(),
            .carryin(bfn_2_22_0_),
            .carryout(\nx.n10690 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_24_lut_LC_2_22_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_24_lut_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_24_lut_LC_2_22_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_24_lut_LC_2_22_1  (
            .in0(N__18315),
            .in1(N__18309),
            .in2(N__18875),
            .in3(N__18300),
            .lcout(\nx.n13193 ),
            .ltout(),
            .carryin(\nx.n10690 ),
            .carryout(\nx.n10691 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_25_lut_LC_2_22_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_25_lut_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_25_lut_LC_2_22_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_25_lut_LC_2_22_2  (
            .in0(N__18297),
            .in1(N__18842),
            .in2(N__18291),
            .in3(N__18279),
            .lcout(\nx.n13195 ),
            .ltout(),
            .carryin(\nx.n10691 ),
            .carryout(\nx.n10692 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_26_lut_LC_2_22_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_26_lut_LC_2_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_26_lut_LC_2_22_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_26_lut_LC_2_22_3  (
            .in0(N__18276),
            .in1(N__18267),
            .in2(N__18818),
            .in3(N__18261),
            .lcout(\nx.n13197 ),
            .ltout(),
            .carryin(\nx.n10692 ),
            .carryout(\nx.n10693 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_27_lut_LC_2_22_4 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_27_lut_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_27_lut_LC_2_22_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_27_lut_LC_2_22_4  (
            .in0(N__18258),
            .in1(N__19897),
            .in2(N__20127),
            .in3(N__18249),
            .lcout(\nx.n13199 ),
            .ltout(),
            .carryin(\nx.n10693 ),
            .carryout(\nx.n10694 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_28_lut_LC_2_22_5 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_28_lut_LC_2_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_28_lut_LC_2_22_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_28_lut_LC_2_22_5  (
            .in0(N__18246),
            .in1(N__23295),
            .in2(N__23327),
            .in3(N__18237),
            .lcout(\nx.n13201 ),
            .ltout(),
            .carryin(\nx.n10694 ),
            .carryout(\nx.n10695 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_28_THRU_CRY_0_LC_2_22_6 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_28_THRU_CRY_0_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_28_THRU_CRY_0_LC_2_22_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_28_THRU_CRY_0_LC_2_22_6  (
            .in0(_gnd_net_),
            .in1(N__42229),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10695 ),
            .carryout(\nx.n10695_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_28_THRU_CRY_1_LC_2_22_7 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_28_THRU_CRY_1_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_28_THRU_CRY_1_LC_2_22_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \nx.sub_14_add_2_28_THRU_CRY_1_LC_2_22_7  (
            .in0(_gnd_net_),
            .in1(N__42224),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\nx.n10695_THRU_CRY_0_THRU_CO ),
            .carryout(\nx.n10695_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_29_lut_LC_2_23_0 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_29_lut_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_29_lut_LC_2_23_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_29_lut_LC_2_23_0  (
            .in0(N__18423),
            .in1(N__18354),
            .in2(N__19089),
            .in3(N__18417),
            .lcout(\nx.n13203 ),
            .ltout(),
            .carryin(bfn_2_23_0_),
            .carryout(\nx.n10696 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_30_lut_LC_2_23_1 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_30_lut_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_30_lut_LC_2_23_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_30_lut_LC_2_23_1  (
            .in0(N__18414),
            .in1(N__23664),
            .in2(N__25268),
            .in3(N__18408),
            .lcout(\nx.n13205 ),
            .ltout(),
            .carryin(\nx.n10696 ),
            .carryout(\nx.n10697 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_31_lut_LC_2_23_2 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_31_lut_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_31_lut_LC_2_23_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_31_lut_LC_2_23_2  (
            .in0(N__18405),
            .in1(N__18399),
            .in2(N__20184),
            .in3(N__18387),
            .lcout(\nx.n13207 ),
            .ltout(),
            .carryin(\nx.n10697 ),
            .carryout(\nx.n10698 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_32_lut_LC_2_23_3 .C_ON=1'b1;
    defparam \nx.sub_14_add_2_32_lut_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_32_lut_LC_2_23_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \nx.sub_14_add_2_32_lut_LC_2_23_3  (
            .in0(N__18384),
            .in1(N__19641),
            .in2(N__21119),
            .in3(N__18378),
            .lcout(\nx.n13209 ),
            .ltout(),
            .carryin(\nx.n10698 ),
            .carryout(\nx.n10699 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_add_2_33_lut_LC_2_23_4 .C_ON=1'b0;
    defparam \nx.sub_14_add_2_33_lut_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_add_2_33_lut_LC_2_23_4 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \nx.sub_14_add_2_33_lut_LC_2_23_4  (
            .in0(N__18375),
            .in1(N__19046),
            .in2(N__18366),
            .in3(N__18357),
            .lcout(\nx.n7608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i28_1_lut_LC_2_23_5 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i28_1_lut_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i28_1_lut_LC_2_23_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i28_1_lut_LC_2_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18347),
            .lcout(\nx.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i27_LC_2_23_6 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i27_LC_2_23_6 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i27_LC_2_23_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i27_LC_2_23_6  (
            .in0(N__18348),
            .in1(N__19088),
            .in2(_gnd_net_),
            .in3(N__25239),
            .lcout(neo_pixel_transmitter_t0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46864),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i6_LC_2_24_0.C_ON=1'b0;
    defparam neopxl_color_i6_LC_2_24_0.SEQ_MODE=4'b1001;
    defparam neopxl_color_i6_LC_2_24_0.LUT_INIT=16'b0101010101000000;
    LogicCell40 neopxl_color_i6_LC_2_24_0 (
            .in0(N__43675),
            .in1(N__43955),
            .in2(N__47697),
            .in3(N__26207),
            .lcout(neopxl_color_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46871),
            .ce(),
            .sr(N__20406));
    defparam \nx.mod_5_i946_3_lut_LC_2_24_6 .C_ON=1'b0;
    defparam \nx.mod_5_i946_3_lut_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i946_3_lut_LC_2_24_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i946_3_lut_LC_2_24_6  (
            .in0(_gnd_net_),
            .in1(N__20367),
            .in2(N__20481),
            .in3(N__20381),
            .lcout(\nx.n1407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i948_3_lut_LC_2_24_7 .C_ON=1'b0;
    defparam \nx.mod_5_i948_3_lut_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i948_3_lut_LC_2_24_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i948_3_lut_LC_2_24_7  (
            .in0(N__20226),
            .in1(N__25482),
            .in2(_gnd_net_),
            .in3(N__20476),
            .lcout(\nx.n1409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_2_lut_LC_2_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_2_lut_LC_2_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_2_lut_LC_2_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_2_lut_LC_2_25_0  (
            .in0(_gnd_net_),
            .in1(N__24096),
            .in2(_gnd_net_),
            .in3(N__18447),
            .lcout(\nx.n1477 ),
            .ltout(),
            .carryin(bfn_2_25_0_),
            .carryout(\nx.n10773 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_3_lut_LC_2_25_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_3_lut_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_3_lut_LC_2_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_3_lut_LC_2_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19608),
            .in3(N__18444),
            .lcout(\nx.n1476 ),
            .ltout(),
            .carryin(\nx.n10773 ),
            .carryout(\nx.n10774 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_4_lut_LC_2_25_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_4_lut_LC_2_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_4_lut_LC_2_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_4_lut_LC_2_25_2  (
            .in0(_gnd_net_),
            .in1(N__42282),
            .in2(N__19571),
            .in3(N__18441),
            .lcout(\nx.n1475 ),
            .ltout(),
            .carryin(\nx.n10774 ),
            .carryout(\nx.n10775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_5_lut_LC_2_25_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_5_lut_LC_2_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_5_lut_LC_2_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_5_lut_LC_2_25_3  (
            .in0(_gnd_net_),
            .in1(N__42288),
            .in2(N__19322),
            .in3(N__18438),
            .lcout(\nx.n1474 ),
            .ltout(),
            .carryin(\nx.n10775 ),
            .carryout(\nx.n10776 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_6_lut_LC_2_25_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_6_lut_LC_2_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_6_lut_LC_2_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_6_lut_LC_2_25_4  (
            .in0(_gnd_net_),
            .in1(N__42283),
            .in2(N__19443),
            .in3(N__18435),
            .lcout(\nx.n1473 ),
            .ltout(),
            .carryin(\nx.n10776 ),
            .carryout(\nx.n10777 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_7_lut_LC_2_25_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_7_lut_LC_2_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_7_lut_LC_2_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_7_lut_LC_2_25_5  (
            .in0(_gnd_net_),
            .in1(N__19388),
            .in2(N__42299),
            .in3(N__18432),
            .lcout(\nx.n1472 ),
            .ltout(),
            .carryin(\nx.n10777 ),
            .carryout(\nx.n10778 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_8_lut_LC_2_25_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_8_lut_LC_2_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_8_lut_LC_2_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_8_lut_LC_2_25_6  (
            .in0(_gnd_net_),
            .in1(N__42287),
            .in2(N__19422),
            .in3(N__18429),
            .lcout(\nx.n1471 ),
            .ltout(),
            .carryin(\nx.n10778 ),
            .carryout(\nx.n10779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_9_lut_LC_2_25_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_9_lut_LC_2_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_9_lut_LC_2_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_9_lut_LC_2_25_7  (
            .in0(_gnd_net_),
            .in1(N__42289),
            .in2(N__19349),
            .in3(N__18426),
            .lcout(\nx.n1470 ),
            .ltout(),
            .carryin(\nx.n10779 ),
            .carryout(\nx.n10780 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_10_lut_LC_2_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_10_lut_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_10_lut_LC_2_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_10_lut_LC_2_26_0  (
            .in0(_gnd_net_),
            .in1(N__19238),
            .in2(N__42300),
            .in3(N__18483),
            .lcout(\nx.n1469 ),
            .ltout(),
            .carryin(bfn_2_26_0_),
            .carryout(\nx.n10781 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_11_lut_LC_2_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1004_11_lut_LC_2_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_11_lut_LC_2_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1004_11_lut_LC_2_26_1  (
            .in0(_gnd_net_),
            .in1(N__42293),
            .in2(N__20436),
            .in3(N__18480),
            .lcout(\nx.n1468 ),
            .ltout(),
            .carryin(\nx.n10781 ),
            .carryout(\nx.n10782 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1004_12_lut_LC_2_26_2 .C_ON=1'b0;
    defparam \nx.mod_5_add_1004_12_lut_LC_2_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1004_12_lut_LC_2_26_2 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1004_12_lut_LC_2_26_2  (
            .in0(N__42294),
            .in1(N__20259),
            .in2(N__19521),
            .in3(N__18477),
            .lcout(\nx.n1499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_134_LC_2_26_4 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_134_LC_2_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_134_LC_2_26_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_134_LC_2_26_4  (
            .in0(N__24105),
            .in1(N__23829),
            .in2(N__30534),
            .in3(N__36060),
            .lcout(\nx.n46_adj_779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1008_3_lut_LC_2_26_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1008_3_lut_LC_2_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1008_3_lut_LC_2_26_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1008_3_lut_LC_2_26_7  (
            .in0(_gnd_net_),
            .in1(N__18474),
            .in2(N__19242),
            .in3(N__19514),
            .lcout(\nx.n1501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i14_LC_3_16_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i14_LC_3_16_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i14_LC_3_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i14_LC_3_16_0  (
            .in0(N__18681),
            .in1(N__18468),
            .in2(_gnd_net_),
            .in3(N__25156),
            .lcout(neo_pixel_transmitter_t0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46846),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i15_1_lut_LC_3_16_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i15_1_lut_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i15_1_lut_LC_3_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i15_1_lut_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18467),
            .lcout(\nx.n19_adj_725 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_done_104_LC_3_17_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_done_104_LC_3_17_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_done_104_LC_3_17_0 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \nx.neo_pixel_transmitter_done_104_LC_3_17_0  (
            .in0(N__24908),
            .in1(N__23250),
            .in2(_gnd_net_),
            .in3(N__23493),
            .lcout(\nx.neo_pixel_transmitter_done ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46842),
            .ce(N__20079),
            .sr(_gnd_net_));
    defparam \nx.i9152_2_lut_LC_3_17_1 .C_ON=1'b0;
    defparam \nx.i9152_2_lut_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9152_2_lut_LC_3_17_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \nx.i9152_2_lut_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__26800),
            .in2(_gnd_net_),
            .in3(N__24907),
            .lcout(),
            .ltout(\nx.n11834_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_151_LC_3_17_2 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_151_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_151_LC_3_17_2 .LUT_INIT=16'b0101000111110001;
    LogicCell40 \nx.i1_4_lut_adj_151_LC_3_17_2  (
            .in0(N__21327),
            .in1(N__21382),
            .in2(N__18627),
            .in3(N__21296),
            .lcout(\nx.n103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i0_LC_3_18_0 .C_ON=1'b1;
    defparam \nx.timer_632__i0_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i0_LC_3_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i0_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__18616),
            .in2(_gnd_net_),
            .in3(N__18597),
            .lcout(timer_0),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\nx.n10707 ),
            .clk(N__46847),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i1_LC_3_18_1 .C_ON=1'b1;
    defparam \nx.timer_632__i1_LC_3_18_1 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i1_LC_3_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i1_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__19741),
            .in2(_gnd_net_),
            .in3(N__18594),
            .lcout(timer_1),
            .ltout(),
            .carryin(\nx.n10707 ),
            .carryout(\nx.n10708 ),
            .clk(N__46847),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i2_LC_3_18_2 .C_ON=1'b1;
    defparam \nx.timer_632__i2_LC_3_18_2 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i2_LC_3_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i2_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(N__18589),
            .in2(_gnd_net_),
            .in3(N__18570),
            .lcout(timer_2),
            .ltout(),
            .carryin(\nx.n10708 ),
            .carryout(\nx.n10709 ),
            .clk(N__46847),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i3_LC_3_18_3 .C_ON=1'b1;
    defparam \nx.timer_632__i3_LC_3_18_3 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i3_LC_3_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i3_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__19708),
            .in2(_gnd_net_),
            .in3(N__18567),
            .lcout(timer_3),
            .ltout(),
            .carryin(\nx.n10709 ),
            .carryout(\nx.n10710 ),
            .clk(N__46847),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i4_LC_3_18_4 .C_ON=1'b1;
    defparam \nx.timer_632__i4_LC_3_18_4 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i4_LC_3_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i4_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(N__18559),
            .in2(_gnd_net_),
            .in3(N__18540),
            .lcout(timer_4),
            .ltout(),
            .carryin(\nx.n10710 ),
            .carryout(\nx.n10711 ),
            .clk(N__46847),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i5_LC_3_18_5 .C_ON=1'b1;
    defparam \nx.timer_632__i5_LC_3_18_5 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i5_LC_3_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i5_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(N__19772),
            .in2(_gnd_net_),
            .in3(N__18537),
            .lcout(timer_5),
            .ltout(),
            .carryin(\nx.n10711 ),
            .carryout(\nx.n10712 ),
            .clk(N__46847),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i6_LC_3_18_6 .C_ON=1'b1;
    defparam \nx.timer_632__i6_LC_3_18_6 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i6_LC_3_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i6_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__18532),
            .in2(_gnd_net_),
            .in3(N__18513),
            .lcout(timer_6),
            .ltout(),
            .carryin(\nx.n10712 ),
            .carryout(\nx.n10713 ),
            .clk(N__46847),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i7_LC_3_18_7 .C_ON=1'b1;
    defparam \nx.timer_632__i7_LC_3_18_7 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i7_LC_3_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i7_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__18505),
            .in2(_gnd_net_),
            .in3(N__18486),
            .lcout(timer_7),
            .ltout(),
            .carryin(\nx.n10713 ),
            .carryout(\nx.n10714 ),
            .clk(N__46847),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i8_LC_3_19_0 .C_ON=1'b1;
    defparam \nx.timer_632__i8_LC_3_19_0 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i8_LC_3_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i8_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__18788),
            .in2(_gnd_net_),
            .in3(N__18771),
            .lcout(timer_8),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\nx.n10715 ),
            .clk(N__46849),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i9_LC_3_19_1 .C_ON=1'b1;
    defparam \nx.timer_632__i9_LC_3_19_1 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i9_LC_3_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i9_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__18764),
            .in2(_gnd_net_),
            .in3(N__18747),
            .lcout(timer_9),
            .ltout(),
            .carryin(\nx.n10715 ),
            .carryout(\nx.n10716 ),
            .clk(N__46849),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i10_LC_3_19_2 .C_ON=1'b1;
    defparam \nx.timer_632__i10_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i10_LC_3_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i10_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__18739),
            .in2(_gnd_net_),
            .in3(N__18720),
            .lcout(timer_10),
            .ltout(),
            .carryin(\nx.n10716 ),
            .carryout(\nx.n10717 ),
            .clk(N__46849),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i11_LC_3_19_3 .C_ON=1'b1;
    defparam \nx.timer_632__i11_LC_3_19_3 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i11_LC_3_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i11_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__21556),
            .in2(_gnd_net_),
            .in3(N__18717),
            .lcout(timer_11),
            .ltout(),
            .carryin(\nx.n10717 ),
            .carryout(\nx.n10718 ),
            .clk(N__46849),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i12_LC_3_19_4 .C_ON=1'b1;
    defparam \nx.timer_632__i12_LC_3_19_4 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i12_LC_3_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i12_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__18706),
            .in2(_gnd_net_),
            .in3(N__18687),
            .lcout(timer_12),
            .ltout(),
            .carryin(\nx.n10718 ),
            .carryout(\nx.n10719 ),
            .clk(N__46849),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i13_LC_3_19_5 .C_ON=1'b1;
    defparam \nx.timer_632__i13_LC_3_19_5 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i13_LC_3_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i13_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__19927),
            .in2(_gnd_net_),
            .in3(N__18684),
            .lcout(timer_13),
            .ltout(),
            .carryin(\nx.n10719 ),
            .carryout(\nx.n10720 ),
            .clk(N__46849),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i14_LC_3_19_6 .C_ON=1'b1;
    defparam \nx.timer_632__i14_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i14_LC_3_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i14_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__18676),
            .in2(_gnd_net_),
            .in3(N__18657),
            .lcout(timer_14),
            .ltout(),
            .carryin(\nx.n10720 ),
            .carryout(\nx.n10721 ),
            .clk(N__46849),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i15_LC_3_19_7 .C_ON=1'b1;
    defparam \nx.timer_632__i15_LC_3_19_7 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i15_LC_3_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i15_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__18649),
            .in2(_gnd_net_),
            .in3(N__18630),
            .lcout(timer_15),
            .ltout(),
            .carryin(\nx.n10721 ),
            .carryout(\nx.n10722 ),
            .clk(N__46849),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i16_LC_3_20_0 .C_ON=1'b1;
    defparam \nx.timer_632__i16_LC_3_20_0 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i16_LC_3_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i16_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__19139),
            .in2(_gnd_net_),
            .in3(N__18996),
            .lcout(timer_16),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\nx.n10723 ),
            .clk(N__46853),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i17_LC_3_20_1 .C_ON=1'b1;
    defparam \nx.timer_632__i17_LC_3_20_1 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i17_LC_3_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i17_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__18988),
            .in2(_gnd_net_),
            .in3(N__18969),
            .lcout(timer_17),
            .ltout(),
            .carryin(\nx.n10723 ),
            .carryout(\nx.n10724 ),
            .clk(N__46853),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i18_LC_3_20_2 .C_ON=1'b1;
    defparam \nx.timer_632__i18_LC_3_20_2 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i18_LC_3_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i18_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__18958),
            .in2(_gnd_net_),
            .in3(N__18939),
            .lcout(timer_18),
            .ltout(),
            .carryin(\nx.n10724 ),
            .carryout(\nx.n10725 ),
            .clk(N__46853),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i19_LC_3_20_3 .C_ON=1'b1;
    defparam \nx.timer_632__i19_LC_3_20_3 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i19_LC_3_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i19_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__19879),
            .in2(_gnd_net_),
            .in3(N__18936),
            .lcout(timer_19),
            .ltout(),
            .carryin(\nx.n10725 ),
            .carryout(\nx.n10726 ),
            .clk(N__46853),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i20_LC_3_20_4 .C_ON=1'b1;
    defparam \nx.timer_632__i20_LC_3_20_4 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i20_LC_3_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i20_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__18926),
            .in2(_gnd_net_),
            .in3(N__18909),
            .lcout(timer_20),
            .ltout(),
            .carryin(\nx.n10726 ),
            .carryout(\nx.n10727 ),
            .clk(N__46853),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i21_LC_3_20_5 .C_ON=1'b1;
    defparam \nx.timer_632__i21_LC_3_20_5 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i21_LC_3_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i21_LC_3_20_5  (
            .in0(_gnd_net_),
            .in1(N__18898),
            .in2(_gnd_net_),
            .in3(N__18879),
            .lcout(timer_21),
            .ltout(),
            .carryin(\nx.n10727 ),
            .carryout(\nx.n10728 ),
            .clk(N__46853),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i22_LC_3_20_6 .C_ON=1'b1;
    defparam \nx.timer_632__i22_LC_3_20_6 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i22_LC_3_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i22_LC_3_20_6  (
            .in0(_gnd_net_),
            .in1(N__18868),
            .in2(_gnd_net_),
            .in3(N__18849),
            .lcout(timer_22),
            .ltout(),
            .carryin(\nx.n10728 ),
            .carryout(\nx.n10729 ),
            .clk(N__46853),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i23_LC_3_20_7 .C_ON=1'b1;
    defparam \nx.timer_632__i23_LC_3_20_7 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i23_LC_3_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i23_LC_3_20_7  (
            .in0(_gnd_net_),
            .in1(N__18841),
            .in2(_gnd_net_),
            .in3(N__18822),
            .lcout(timer_23),
            .ltout(),
            .carryin(\nx.n10729 ),
            .carryout(\nx.n10730 ),
            .clk(N__46853),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i24_LC_3_21_0 .C_ON=1'b1;
    defparam \nx.timer_632__i24_LC_3_21_0 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i24_LC_3_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i24_LC_3_21_0  (
            .in0(_gnd_net_),
            .in1(N__18814),
            .in2(_gnd_net_),
            .in3(N__18795),
            .lcout(timer_24),
            .ltout(),
            .carryin(bfn_3_21_0_),
            .carryout(\nx.n10731 ),
            .clk(N__46859),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i25_LC_3_21_1 .C_ON=1'b1;
    defparam \nx.timer_632__i25_LC_3_21_1 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i25_LC_3_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i25_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(N__19898),
            .in2(_gnd_net_),
            .in3(N__19095),
            .lcout(timer_25),
            .ltout(),
            .carryin(\nx.n10731 ),
            .carryout(\nx.n10732 ),
            .clk(N__46859),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i26_LC_3_21_2 .C_ON=1'b1;
    defparam \nx.timer_632__i26_LC_3_21_2 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i26_LC_3_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i26_LC_3_21_2  (
            .in0(_gnd_net_),
            .in1(N__23323),
            .in2(_gnd_net_),
            .in3(N__19092),
            .lcout(timer_26),
            .ltout(),
            .carryin(\nx.n10732 ),
            .carryout(\nx.n10733 ),
            .clk(N__46859),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i27_LC_3_21_3 .C_ON=1'b1;
    defparam \nx.timer_632__i27_LC_3_21_3 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i27_LC_3_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i27_LC_3_21_3  (
            .in0(_gnd_net_),
            .in1(N__19084),
            .in2(_gnd_net_),
            .in3(N__19062),
            .lcout(timer_27),
            .ltout(),
            .carryin(\nx.n10733 ),
            .carryout(\nx.n10734 ),
            .clk(N__46859),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i28_LC_3_21_4 .C_ON=1'b1;
    defparam \nx.timer_632__i28_LC_3_21_4 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i28_LC_3_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i28_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(N__25258),
            .in2(_gnd_net_),
            .in3(N__19059),
            .lcout(timer_28),
            .ltout(),
            .carryin(\nx.n10734 ),
            .carryout(\nx.n10735 ),
            .clk(N__46859),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i29_LC_3_21_5 .C_ON=1'b1;
    defparam \nx.timer_632__i29_LC_3_21_5 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i29_LC_3_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i29_LC_3_21_5  (
            .in0(_gnd_net_),
            .in1(N__20176),
            .in2(_gnd_net_),
            .in3(N__19056),
            .lcout(timer_29),
            .ltout(),
            .carryin(\nx.n10735 ),
            .carryout(\nx.n10736 ),
            .clk(N__46859),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i30_LC_3_21_6 .C_ON=1'b1;
    defparam \nx.timer_632__i30_LC_3_21_6 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i30_LC_3_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i30_LC_3_21_6  (
            .in0(_gnd_net_),
            .in1(N__21109),
            .in2(_gnd_net_),
            .in3(N__19053),
            .lcout(timer_30),
            .ltout(),
            .carryin(\nx.n10736 ),
            .carryout(\nx.n10737 ),
            .clk(N__46859),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.timer_632__i31_LC_3_21_7 .C_ON=1'b0;
    defparam \nx.timer_632__i31_LC_3_21_7 .SEQ_MODE=4'b1000;
    defparam \nx.timer_632__i31_LC_3_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.timer_632__i31_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(N__19045),
            .in2(_gnd_net_),
            .in3(N__19050),
            .lcout(timer_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46859),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_184_LC_3_22_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_184_LC_3_22_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_184_LC_3_22_0.LUT_INIT=16'b1100110011001000;
    LogicCell40 i1_2_lut_3_lut_4_lut_4_lut_adj_184_LC_3_22_0 (
            .in0(N__45020),
            .in1(N__47667),
            .in2(N__45695),
            .in3(N__42639),
            .lcout(),
            .ltout(n11826_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i1_LC_3_22_1.C_ON=1'b0;
    defparam pin_output_enable__i1_LC_3_22_1.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i1_LC_3_22_1.LUT_INIT=16'b1100111011000100;
    LogicCell40 pin_output_enable__i1_LC_3_22_1 (
            .in0(N__47125),
            .in1(N__19007),
            .in2(N__19023),
            .in3(N__47672),
            .lcout(pin_oe_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46865),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_3_22_2.C_ON=1'b0;
    defparam i4_4_lut_LC_3_22_2.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_3_22_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i4_4_lut_LC_3_22_2 (
            .in0(N__19221),
            .in1(N__20583),
            .in2(N__19203),
            .in3(N__19182),
            .lcout(n12379),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_187_LC_3_22_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_187_LC_3_22_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_187_LC_3_22_3.LUT_INIT=16'b1010101010001010;
    LogicCell40 i1_2_lut_3_lut_4_lut_4_lut_adj_187_LC_3_22_3 (
            .in0(N__47666),
            .in1(N__42635),
            .in2(N__45696),
            .in3(N__45021),
            .lcout(),
            .ltout(n11828_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i5_LC_3_22_4.C_ON=1'b0;
    defparam pin_output_enable__i5_LC_3_22_4.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i5_LC_3_22_4.LUT_INIT=16'b1010110010101010;
    LogicCell40 pin_output_enable__i5_LC_3_22_4 (
            .in0(N__19154),
            .in1(N__47668),
            .in2(N__19170),
            .in3(N__47126),
            .lcout(pin_oe_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46865),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i16_LC_3_22_5 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i16_LC_3_22_5 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i16_LC_3_22_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i16_LC_3_22_5  (
            .in0(N__19143),
            .in1(N__19122),
            .in2(_gnd_net_),
            .in3(N__25220),
            .lcout(neo_pixel_transmitter_t0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46865),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i874_3_lut_LC_3_22_7 .C_ON=1'b0;
    defparam \nx.mod_5_i874_3_lut_LC_3_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i874_3_lut_LC_3_22_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i874_3_lut_LC_3_22_7  (
            .in0(_gnd_net_),
            .in1(N__22095),
            .in2(N__22119),
            .in3(N__21980),
            .lcout(\nx.n1303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i944_3_lut_LC_3_23_0 .C_ON=1'b0;
    defparam \nx.mod_5_i944_3_lut_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i944_3_lut_LC_3_23_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i944_3_lut_LC_3_23_0  (
            .in0(N__20342),
            .in1(_gnd_net_),
            .in2(N__20325),
            .in3(N__20467),
            .lcout(\nx.n1405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i17_1_lut_LC_3_23_1 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i17_1_lut_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i17_1_lut_LC_3_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i17_1_lut_LC_3_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19121),
            .lcout(\nx.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i880_3_lut_LC_3_23_2 .C_ON=1'b0;
    defparam \nx.mod_5_i880_3_lut_LC_3_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i880_3_lut_LC_3_23_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i880_3_lut_LC_3_23_2  (
            .in0(N__21777),
            .in1(N__24053),
            .in2(_gnd_net_),
            .in3(N__21965),
            .lcout(\nx.n1309 ),
            .ltout(\nx.n1309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_3_lut_LC_3_23_3 .C_ON=1'b0;
    defparam \nx.i3_3_lut_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.i3_3_lut_LC_3_23_3 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \nx.i3_3_lut_LC_3_23_3  (
            .in0(_gnd_net_),
            .in1(N__25477),
            .in2(N__19098),
            .in3(N__20341),
            .lcout(\nx.n12_adj_669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_158_LC_3_23_4.C_ON=1'b0;
    defparam i6_4_lut_adj_158_LC_3_23_4.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_158_LC_3_23_4.LUT_INIT=16'b1111111011111010;
    LogicCell40 i6_4_lut_adj_158_LC_3_23_4 (
            .in0(N__19302),
            .in1(N__22008),
            .in2(N__19284),
            .in3(N__19263),
            .lcout(n17_adj_816),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i879_3_lut_LC_3_23_5 .C_ON=1'b0;
    defparam \nx.mod_5_i879_3_lut_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i879_3_lut_LC_3_23_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i879_3_lut_LC_3_23_5  (
            .in0(_gnd_net_),
            .in1(N__21761),
            .in2(N__21981),
            .in3(N__21741),
            .lcout(\nx.n1308 ),
            .ltout(\nx.n1308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8_4_lut_LC_3_23_6 .C_ON=1'b0;
    defparam \nx.i8_4_lut_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.i8_4_lut_LC_3_23_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i8_4_lut_LC_3_23_6  (
            .in0(N__19257),
            .in1(N__20290),
            .in2(N__19251),
            .in3(N__20496),
            .lcout(\nx.n1334 ),
            .ltout(\nx.n1334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i941_3_lut_LC_3_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i941_3_lut_LC_3_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i941_3_lut_LC_3_23_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i941_3_lut_LC_3_23_7  (
            .in0(N__20291),
            .in1(_gnd_net_),
            .in2(N__19248),
            .in3(N__20274),
            .lcout(\nx.n1402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9149_3_lut_LC_3_24_1 .C_ON=1'b0;
    defparam \nx.i9149_3_lut_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9149_3_lut_LC_3_24_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.i9149_3_lut_LC_3_24_1  (
            .in0(_gnd_net_),
            .in1(N__20313),
            .in2(N__20550),
            .in3(N__20475),
            .lcout(\nx.n1404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i945_3_lut_LC_3_24_2 .C_ON=1'b0;
    defparam \nx.mod_5_i945_3_lut_LC_3_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i945_3_lut_LC_3_24_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i945_3_lut_LC_3_24_2  (
            .in0(_gnd_net_),
            .in1(N__20352),
            .in2(N__20480),
            .in3(N__20519),
            .lcout(\nx.n1406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i942_3_lut_LC_3_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i942_3_lut_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i942_3_lut_LC_3_24_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i942_3_lut_LC_3_24_3  (
            .in0(_gnd_net_),
            .in1(N__20573),
            .in2(N__20304),
            .in3(N__20474),
            .lcout(\nx.n1403 ),
            .ltout(\nx.n1403_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_3_lut_adj_72_LC_3_24_4 .C_ON=1'b0;
    defparam \nx.i3_3_lut_adj_72_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.i3_3_lut_adj_72_LC_3_24_4 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i3_3_lut_adj_72_LC_3_24_4  (
            .in0(_gnd_net_),
            .in1(N__24103),
            .in2(N__19245),
            .in3(N__19603),
            .lcout(\nx.n13_adj_729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_4_lut_adj_71_LC_3_24_5 .C_ON=1'b0;
    defparam \nx.i6_4_lut_adj_71_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.i6_4_lut_adj_71_LC_3_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i6_4_lut_adj_71_LC_3_24_5  (
            .in0(N__20252),
            .in1(N__19232),
            .in2(N__19387),
            .in3(N__20422),
            .lcout(),
            .ltout(\nx.n16_adj_727_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8_3_lut_LC_3_24_6 .C_ON=1'b0;
    defparam \nx.i8_3_lut_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.i8_3_lut_LC_3_24_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \nx.i8_3_lut_LC_3_24_6  (
            .in0(_gnd_net_),
            .in1(N__19438),
            .in2(N__19461),
            .in3(N__19564),
            .lcout(\nx.n18_adj_728 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i947_3_lut_LC_3_24_7 .C_ON=1'b0;
    defparam \nx.mod_5_i947_3_lut_LC_3_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i947_3_lut_LC_3_24_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i947_3_lut_LC_3_24_7  (
            .in0(_gnd_net_),
            .in1(N__20210),
            .in2(N__20196),
            .in3(N__20470),
            .lcout(\nx.n1408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1010_3_lut_LC_3_25_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1010_3_lut_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1010_3_lut_LC_3_25_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1010_3_lut_LC_3_25_0  (
            .in0(_gnd_net_),
            .in1(N__19418),
            .in2(N__19458),
            .in3(N__19505),
            .lcout(\nx.n1503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1012_3_lut_LC_3_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1012_3_lut_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1012_3_lut_LC_3_25_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1012_3_lut_LC_3_25_1  (
            .in0(N__19449),
            .in1(_gnd_net_),
            .in2(N__19520),
            .in3(N__19442),
            .lcout(\nx.n1505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_73_LC_3_25_2 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_73_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_73_LC_3_25_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_adj_73_LC_3_25_2  (
            .in0(N__19318),
            .in1(N__19417),
            .in2(N__19404),
            .in3(N__19395),
            .lcout(\nx.n1433 ),
            .ltout(\nx.n1433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1011_3_lut_LC_3_25_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1011_3_lut_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1011_3_lut_LC_3_25_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1011_3_lut_LC_3_25_3  (
            .in0(_gnd_net_),
            .in1(N__19389),
            .in2(N__19365),
            .in3(N__19362),
            .lcout(\nx.n1504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1009_3_lut_LC_3_25_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1009_3_lut_LC_3_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1009_3_lut_LC_3_25_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1009_3_lut_LC_3_25_4  (
            .in0(_gnd_net_),
            .in1(N__19356),
            .in2(N__19350),
            .in3(N__19509),
            .lcout(\nx.n1502 ),
            .ltout(\nx.n1502_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_2_lut_LC_3_25_5 .C_ON=1'b0;
    defparam \nx.i5_2_lut_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.i5_2_lut_LC_3_25_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i5_2_lut_LC_3_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19332),
            .in3(N__21007),
            .lcout(\nx.n16_adj_732 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1013_3_lut_LC_3_25_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1013_3_lut_LC_3_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1013_3_lut_LC_3_25_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1013_3_lut_LC_3_25_6  (
            .in0(_gnd_net_),
            .in1(N__19329),
            .in2(N__19323),
            .in3(N__19513),
            .lcout(\nx.n1506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1015_3_lut_LC_3_25_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1015_3_lut_LC_3_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1015_3_lut_LC_3_25_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1015_3_lut_LC_3_25_7  (
            .in0(_gnd_net_),
            .in1(N__19614),
            .in2(N__19519),
            .in3(N__19607),
            .lcout(\nx.n1508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1007_3_lut_LC_3_26_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1007_3_lut_LC_3_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1007_3_lut_LC_3_26_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1007_3_lut_LC_3_26_0  (
            .in0(_gnd_net_),
            .in1(N__20432),
            .in2(N__19587),
            .in3(N__19501),
            .lcout(\nx.n1500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1014_3_lut_LC_3_26_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1014_3_lut_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1014_3_lut_LC_3_26_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1014_3_lut_LC_3_26_1  (
            .in0(_gnd_net_),
            .in1(N__19578),
            .in2(N__19518),
            .in3(N__19572),
            .lcout(\nx.n1507 ),
            .ltout(\nx.n1507_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_4_lut_adj_75_LC_3_26_2 .C_ON=1'b0;
    defparam \nx.i7_4_lut_adj_75_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.i7_4_lut_adj_75_LC_3_26_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i7_4_lut_adj_75_LC_3_26_2  (
            .in0(N__21028),
            .in1(N__20689),
            .in2(N__19548),
            .in3(N__19467),
            .lcout(),
            .ltout(\nx.n18_adj_731_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_76_LC_3_26_3 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_76_LC_3_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_76_LC_3_26_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_adj_76_LC_3_26_3  (
            .in0(N__20632),
            .in1(N__20957),
            .in2(N__19545),
            .in3(N__20941),
            .lcout(),
            .ltout(\nx.n20_adj_733_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_77_LC_3_26_4 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_77_LC_3_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_77_LC_3_26_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_77_LC_3_26_4  (
            .in0(N__20909),
            .in1(N__20653),
            .in2(N__19542),
            .in3(N__19539),
            .lcout(\nx.n1532 ),
            .ltout(\nx.n1532_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9208_1_lut_LC_3_26_5 .C_ON=1'b0;
    defparam \nx.i9208_1_lut_LC_3_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9208_1_lut_LC_3_26_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \nx.i9208_1_lut_LC_3_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19533),
            .in3(_gnd_net_),
            .lcout(\nx.n13604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1016_3_lut_LC_3_26_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1016_3_lut_LC_3_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1016_3_lut_LC_3_26_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1016_3_lut_LC_3_26_6  (
            .in0(N__19530),
            .in1(N__24104),
            .in2(_gnd_net_),
            .in3(N__19500),
            .lcout(\nx.n1509 ),
            .ltout(\nx.n1509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5936_2_lut_LC_3_26_7 .C_ON=1'b0;
    defparam \nx.i5936_2_lut_LC_3_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.i5936_2_lut_LC_3_26_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \nx.i5936_2_lut_LC_3_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19470),
            .in3(N__23826),
            .lcout(\nx.n9729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i26_4_lut_adj_139_LC_3_27_7 .C_ON=1'b0;
    defparam \nx.i26_4_lut_adj_139_LC_3_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.i26_4_lut_adj_139_LC_3_27_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i26_4_lut_adj_139_LC_3_27_7  (
            .in0(N__20808),
            .in1(N__19647),
            .in2(N__24717),
            .in3(N__20823),
            .lcout(\nx.n54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.start_103_LC_4_16_0 .C_ON=1'b0;
    defparam \nx.start_103_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \nx.start_103_LC_4_16_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \nx.start_103_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__23249),
            .in2(_gnd_net_),
            .in3(N__23492),
            .lcout(\nx.start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46850),
            .ce(N__19620),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i31_1_lut_LC_4_16_1 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i31_1_lut_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i31_1_lut_LC_4_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i31_1_lut_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21089),
            .lcout(\nx.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_adj_116_LC_4_17_0 .C_ON=1'b0;
    defparam \nx.i20_4_lut_adj_116_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_adj_116_LC_4_17_0 .LUT_INIT=16'b1100111011001111;
    LogicCell40 \nx.i20_4_lut_adj_116_LC_4_17_0  (
            .in0(N__24945),
            .in1(N__23470),
            .in2(N__23259),
            .in3(N__21078),
            .lcout(),
            .ltout(\nx.n7_adj_764_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_118_LC_4_17_1 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_118_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_118_LC_4_17_1 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \nx.i1_4_lut_adj_118_LC_4_17_1  (
            .in0(N__21348),
            .in1(N__22872),
            .in2(N__19626),
            .in3(N__23479),
            .lcout(n11353),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7535_3_lut_LC_4_17_2 .C_ON=1'b0;
    defparam \nx.i7535_3_lut_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \nx.i7535_3_lut_LC_4_17_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \nx.i7535_3_lut_LC_4_17_2  (
            .in0(N__23248),
            .in1(N__24933),
            .in2(_gnd_net_),
            .in3(N__21347),
            .lcout(),
            .ltout(\nx.n11864_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_150_LC_4_17_3 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_150_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_150_LC_4_17_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \nx.i15_4_lut_adj_150_LC_4_17_3  (
            .in0(N__21390),
            .in1(N__23480),
            .in2(N__19623),
            .in3(N__21269),
            .lcout(\nx.n7_adj_667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7561_2_lut_LC_4_17_4 .C_ON=1'b0;
    defparam \nx.i7561_2_lut_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \nx.i7561_2_lut_LC_4_17_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \nx.i7561_2_lut_LC_4_17_4  (
            .in0(N__23243),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23469),
            .lcout(\nx.n11892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9093_2_lut_3_lut_LC_4_17_6 .C_ON=1'b0;
    defparam \nx.i9093_2_lut_3_lut_LC_4_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9093_2_lut_3_lut_LC_4_17_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \nx.i9093_2_lut_3_lut_LC_4_17_6  (
            .in0(N__23244),
            .in1(N__21333),
            .in2(_gnd_net_),
            .in3(N__21384),
            .lcout(\nx.n13445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_4_lut_adj_152_LC_4_18_0 .C_ON=1'b0;
    defparam \nx.i6_4_lut_adj_152_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.i6_4_lut_adj_152_LC_4_18_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \nx.i6_4_lut_adj_152_LC_4_18_0  (
            .in0(N__19989),
            .in1(N__19830),
            .in2(N__19824),
            .in3(N__20067),
            .lcout(\nx.n16_adj_785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i4_1_lut_LC_4_18_1 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i4_1_lut_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i4_1_lut_LC_4_18_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \nx.sub_14_inv_0_i4_1_lut_LC_4_18_1  (
            .in0(_gnd_net_),
            .in1(N__19688),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\nx.n30_adj_712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i2_1_lut_LC_4_18_3 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i2_1_lut_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i2_1_lut_LC_4_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i2_1_lut_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19718),
            .lcout(\nx.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i6_1_lut_LC_4_18_4 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i6_1_lut_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i6_1_lut_LC_4_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i6_1_lut_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19751),
            .lcout(\nx.n28_adj_715 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i5_LC_4_18_5 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i5_LC_4_18_5 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i5_LC_4_18_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i5_LC_4_18_5  (
            .in0(N__25117),
            .in1(_gnd_net_),
            .in2(N__19755),
            .in3(N__19773),
            .lcout(neo_pixel_transmitter_t0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46851),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i1_LC_4_18_6 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i1_LC_4_18_6 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i1_LC_4_18_6 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i1_LC_4_18_6  (
            .in0(N__19742),
            .in1(N__25116),
            .in2(N__19722),
            .in3(_gnd_net_),
            .lcout(neo_pixel_transmitter_t0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46851),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_147_LC_4_18_7 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_147_LC_4_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_147_LC_4_18_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \nx.i1_2_lut_adj_147_LC_4_18_7  (
            .in0(_gnd_net_),
            .in1(N__19670),
            .in2(_gnd_net_),
            .in3(N__20100),
            .lcout(\nx.n13211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i3_LC_4_19_0 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i3_LC_4_19_0 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i3_LC_4_19_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i3_LC_4_19_0  (
            .in0(N__25166),
            .in1(N__19709),
            .in2(_gnd_net_),
            .in3(N__19689),
            .lcout(neo_pixel_transmitter_t0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46854),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_153_LC_4_19_1 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_153_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_153_LC_4_19_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \nx.i1_4_lut_adj_153_LC_4_19_1  (
            .in0(N__20049),
            .in1(N__19677),
            .in2(N__19671),
            .in3(N__19962),
            .lcout(),
            .ltout(\nx.n6_adj_786_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_4_lut_adj_154_LC_4_19_2 .C_ON=1'b0;
    defparam \nx.i4_4_lut_adj_154_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.i4_4_lut_adj_154_LC_4_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i4_4_lut_adj_154_LC_4_19_2  (
            .in0(N__20030),
            .in1(N__20009),
            .in2(N__20103),
            .in3(N__20099),
            .lcout(\nx.n13659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5953_4_lut_LC_4_19_3 .C_ON=1'b0;
    defparam \nx.i5953_4_lut_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.i5953_4_lut_LC_4_19_3 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \nx.i5953_4_lut_LC_4_19_3  (
            .in0(N__20048),
            .in1(N__19988),
            .in2(N__20010),
            .in3(N__19961),
            .lcout(\nx.n9747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_148_LC_4_19_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_148_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_148_LC_4_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_148_LC_4_19_4  (
            .in0(N__20063),
            .in1(N__20047),
            .in2(N__20031),
            .in3(N__20016),
            .lcout(),
            .ltout(\nx.n13217_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_149_LC_4_19_5 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_149_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_149_LC_4_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_149_LC_4_19_5  (
            .in0(N__20005),
            .in1(N__19987),
            .in2(N__19965),
            .in3(N__19960),
            .lcout(\nx.n7564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i14_1_lut_LC_4_19_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i14_1_lut_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i14_1_lut_LC_4_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i14_1_lut_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19907),
            .lcout(\nx.n20_adj_726 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_7  (
            .in0(N__19908),
            .in1(N__19928),
            .in2(_gnd_net_),
            .in3(N__25165),
            .lcout(neo_pixel_transmitter_t0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46854),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_1 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_1 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_1  (
            .in0(N__19899),
            .in1(N__20139),
            .in2(_gnd_net_),
            .in3(N__25217),
            .lcout(neo_pixel_transmitter_t0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46860),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i19_LC_4_20_3 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i19_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i19_LC_4_20_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i19_LC_4_20_3  (
            .in0(N__19880),
            .in1(N__21414),
            .in2(_gnd_net_),
            .in3(N__25216),
            .lcout(neo_pixel_transmitter_t0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46860),
            .ce(),
            .sr(_gnd_net_));
    defparam i8987_3_lut_LC_4_20_4.C_ON=1'b0;
    defparam i8987_3_lut_LC_4_20_4.SEQ_MODE=4'b0000;
    defparam i8987_3_lut_LC_4_20_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 i8987_3_lut_LC_4_20_4 (
            .in0(N__19860),
            .in1(N__19842),
            .in2(_gnd_net_),
            .in3(N__46410),
            .lcout(n13382),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_20_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_20_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_20_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_20_7  (
            .in0(N__20177),
            .in1(N__20153),
            .in2(_gnd_net_),
            .in3(N__25218),
            .lcout(neo_pixel_transmitter_t0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46860),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i809_rep_49_3_lut_LC_4_21_0 .C_ON=1'b0;
    defparam \nx.mod_5_i809_rep_49_3_lut_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i809_rep_49_3_lut_LC_4_21_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i809_rep_49_3_lut_LC_4_21_0  (
            .in0(_gnd_net_),
            .in1(N__23628),
            .in2(N__21576),
            .in3(N__21816),
            .lcout(\nx.n1206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i26_1_lut_LC_4_21_2 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i26_1_lut_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i26_1_lut_LC_4_21_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \nx.sub_14_inv_0_i26_1_lut_LC_4_21_2  (
            .in0(_gnd_net_),
            .in1(N__20138),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\nx.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i808_3_lut_LC_4_21_3 .C_ON=1'b0;
    defparam \nx.mod_5_i808_3_lut_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i808_3_lut_LC_4_21_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i808_3_lut_LC_4_21_3  (
            .in0(_gnd_net_),
            .in1(N__21899),
            .in2(N__21827),
            .in3(N__21879),
            .lcout(\nx.n1205 ),
            .ltout(\nx.n1205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_3_lut_adj_18_LC_4_21_4 .C_ON=1'b0;
    defparam \nx.i3_3_lut_adj_18_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.i3_3_lut_adj_18_LC_4_21_4 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i3_3_lut_adj_18_LC_4_21_4  (
            .in0(_gnd_net_),
            .in1(N__24054),
            .in2(N__20112),
            .in3(N__21760),
            .lcout(\nx.n11_adj_674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i810_3_lut_LC_4_21_5 .C_ON=1'b0;
    defparam \nx.mod_5_i810_3_lut_LC_4_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i810_3_lut_LC_4_21_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i810_3_lut_LC_4_21_5  (
            .in0(_gnd_net_),
            .in1(N__21605),
            .in2(N__21826),
            .in3(N__21585),
            .lcout(\nx.n1207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i811_3_lut_LC_4_21_6 .C_ON=1'b0;
    defparam \nx.mod_5_i811_3_lut_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i811_3_lut_LC_4_21_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i811_3_lut_LC_4_21_6  (
            .in0(_gnd_net_),
            .in1(N__21632),
            .in2(N__21618),
            .in3(N__21809),
            .lcout(\nx.n1208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i807_3_lut_LC_4_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_i807_3_lut_LC_4_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i807_3_lut_LC_4_21_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i807_3_lut_LC_4_21_7  (
            .in0(_gnd_net_),
            .in1(N__23517),
            .in2(N__21825),
            .in3(N__21870),
            .lcout(\nx.n1204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_4_lut_adj_20_LC_4_22_0 .C_ON=1'b0;
    defparam \nx.i7_4_lut_adj_20_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.i7_4_lut_adj_20_LC_4_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i7_4_lut_adj_20_LC_4_22_0  (
            .in0(N__21670),
            .in1(N__21697),
            .in2(N__20235),
            .in3(N__20109),
            .lcout(\nx.n1235 ),
            .ltout(\nx.n1235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i875_3_lut_LC_4_22_1 .C_ON=1'b0;
    defparam \nx.mod_5_i875_3_lut_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i875_3_lut_LC_4_22_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i875_3_lut_LC_4_22_1  (
            .in0(_gnd_net_),
            .in1(N__22142),
            .in2(N__20241),
            .in3(N__22128),
            .lcout(\nx.n1304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i812_3_lut_LC_4_22_2 .C_ON=1'b0;
    defparam \nx.mod_5_i812_3_lut_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i812_3_lut_LC_4_22_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i812_3_lut_LC_4_22_2  (
            .in0(N__21645),
            .in1(N__24000),
            .in2(_gnd_net_),
            .in3(N__21821),
            .lcout(\nx.n1209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i806_3_lut_LC_4_22_3 .C_ON=1'b0;
    defparam \nx.mod_5_i806_3_lut_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i806_3_lut_LC_4_22_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i806_3_lut_LC_4_22_3  (
            .in0(_gnd_net_),
            .in1(N__21861),
            .in2(N__21828),
            .in3(N__21837),
            .lcout(\nx.n1203 ),
            .ltout(\nx.n1203_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_4_lut_adj_19_LC_4_22_4 .C_ON=1'b0;
    defparam \nx.i5_4_lut_adj_19_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.i5_4_lut_adj_19_LC_4_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i5_4_lut_adj_19_LC_4_22_4  (
            .in0(N__22073),
            .in1(N__21724),
            .in2(N__20238),
            .in3(N__22111),
            .lcout(\nx.n13_adj_675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i878_3_lut_LC_4_22_5 .C_ON=1'b0;
    defparam \nx.mod_5_i878_3_lut_LC_4_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i878_3_lut_LC_4_22_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i878_3_lut_LC_4_22_5  (
            .in0(N__21725),
            .in1(_gnd_net_),
            .in2(N__21983),
            .in3(N__21708),
            .lcout(\nx.n1307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i876_3_lut_LC_4_22_6 .C_ON=1'b0;
    defparam \nx.mod_5_i876_3_lut_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i876_3_lut_LC_4_22_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i876_3_lut_LC_4_22_6  (
            .in0(N__21671),
            .in1(_gnd_net_),
            .in2(N__22155),
            .in3(N__21973),
            .lcout(\nx.n1305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i877_3_lut_LC_4_22_7 .C_ON=1'b0;
    defparam \nx.mod_5_i877_3_lut_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i877_3_lut_LC_4_22_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i877_3_lut_LC_4_22_7  (
            .in0(N__21698),
            .in1(_gnd_net_),
            .in2(N__21984),
            .in3(N__21681),
            .lcout(\nx.n1306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_2_lut_LC_4_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_2_lut_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_2_lut_LC_4_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_2_lut_LC_4_23_0  (
            .in0(_gnd_net_),
            .in1(N__25476),
            .in2(_gnd_net_),
            .in3(N__20214),
            .lcout(\nx.n1377 ),
            .ltout(),
            .carryin(bfn_4_23_0_),
            .carryout(\nx.n10764 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_3_lut_LC_4_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_3_lut_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_3_lut_LC_4_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_3_lut_LC_4_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20211),
            .in3(N__20187),
            .lcout(\nx.n1376 ),
            .ltout(),
            .carryin(\nx.n10764 ),
            .carryout(\nx.n10765 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_4_lut_LC_4_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_4_lut_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_4_lut_LC_4_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_4_lut_LC_4_23_2  (
            .in0(_gnd_net_),
            .in1(N__41610),
            .in2(N__20382),
            .in3(N__20355),
            .lcout(\nx.n1375 ),
            .ltout(),
            .carryin(\nx.n10765 ),
            .carryout(\nx.n10766 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_5_lut_LC_4_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_5_lut_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_5_lut_LC_4_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_5_lut_LC_4_23_3  (
            .in0(_gnd_net_),
            .in1(N__41613),
            .in2(N__20520),
            .in3(N__20346),
            .lcout(\nx.n1374 ),
            .ltout(),
            .carryin(\nx.n10766 ),
            .carryout(\nx.n10767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_6_lut_LC_4_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_6_lut_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_6_lut_LC_4_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_6_lut_LC_4_23_4  (
            .in0(_gnd_net_),
            .in1(N__41611),
            .in2(N__20343),
            .in3(N__20316),
            .lcout(\nx.n1373 ),
            .ltout(),
            .carryin(\nx.n10767 ),
            .carryout(\nx.n10768 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_7_lut_LC_4_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_7_lut_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_7_lut_LC_4_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_7_lut_LC_4_23_5  (
            .in0(_gnd_net_),
            .in1(N__41614),
            .in2(N__20549),
            .in3(N__20307),
            .lcout(\nx.n1372 ),
            .ltout(),
            .carryin(\nx.n10768 ),
            .carryout(\nx.n10769 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_8_lut_LC_4_23_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_8_lut_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_8_lut_LC_4_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_8_lut_LC_4_23_6  (
            .in0(_gnd_net_),
            .in1(N__41612),
            .in2(N__20574),
            .in3(N__20295),
            .lcout(\nx.n1371 ),
            .ltout(),
            .carryin(\nx.n10769 ),
            .carryout(\nx.n10770 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_9_lut_LC_4_23_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_9_lut_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_9_lut_LC_4_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_9_lut_LC_4_23_7  (
            .in0(_gnd_net_),
            .in1(N__41615),
            .in2(N__20292),
            .in3(N__20268),
            .lcout(\nx.n1370 ),
            .ltout(),
            .carryin(\nx.n10770 ),
            .carryout(\nx.n10771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_10_lut_LC_4_24_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_937_10_lut_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_10_lut_LC_4_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_937_10_lut_LC_4_24_0  (
            .in0(_gnd_net_),
            .in1(N__42279),
            .in2(N__21930),
            .in3(N__20265),
            .lcout(\nx.n1369 ),
            .ltout(),
            .carryin(bfn_4_24_0_),
            .carryout(\nx.n10772 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_937_11_lut_LC_4_24_1 .C_ON=1'b0;
    defparam \nx.mod_5_add_937_11_lut_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_937_11_lut_LC_4_24_1 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_937_11_lut_LC_4_24_1  (
            .in0(N__42280),
            .in1(N__20469),
            .in2(N__22059),
            .in3(N__20262),
            .lcout(\nx.n1400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_156_LC_4_24_2.C_ON=1'b0;
    defparam i1_2_lut_adj_156_LC_4_24_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_156_LC_4_24_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_156_LC_4_24_2 (
            .in0(_gnd_net_),
            .in1(N__20613),
            .in2(_gnd_net_),
            .in3(N__20598),
            .lcout(n6_adj_843),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_LC_4_24_3 .C_ON=1'b0;
    defparam \nx.i1_2_lut_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_LC_4_24_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i1_2_lut_LC_4_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22058),
            .in3(N__21925),
            .lcout(),
            .ltout(\nx.n10_adj_668_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_4_lut_LC_4_24_4 .C_ON=1'b0;
    defparam \nx.i7_4_lut_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.i7_4_lut_LC_4_24_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i7_4_lut_LC_4_24_4  (
            .in0(N__20572),
            .in1(N__20545),
            .in2(N__20523),
            .in3(N__20518),
            .lcout(\nx.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i940_3_lut_LC_4_24_5 .C_ON=1'b0;
    defparam \nx.mod_5_i940_3_lut_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i940_3_lut_LC_4_24_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i940_3_lut_LC_4_24_5  (
            .in0(_gnd_net_),
            .in1(N__21929),
            .in2(N__20490),
            .in3(N__20468),
            .lcout(\nx.n1401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_185_LC_4_24_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_185_LC_4_24_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_185_LC_4_24_7.LUT_INIT=16'b1111101000000000;
    LogicCell40 i1_2_lut_3_lut_adj_185_LC_4_24_7 (
            .in0(N__47665),
            .in1(_gnd_net_),
            .in2(N__43940),
            .in3(N__26209),
            .lcout(n22_adj_795),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_LC_4_25_1 .C_ON=1'b0;
    defparam \nx.i11_4_lut_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_LC_4_25_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_LC_4_25_1  (
            .in0(N__22216),
            .in1(N__20799),
            .in2(N__22536),
            .in3(N__20388),
            .lcout(\nx.n1631 ),
            .ltout(\nx.n1631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9206_1_lut_LC_4_25_2 .C_ON=1'b0;
    defparam \nx.i9206_1_lut_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9206_1_lut_LC_4_25_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \nx.i9206_1_lut_LC_4_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20394),
            .in3(_gnd_net_),
            .lcout(\nx.n13602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_3_lut_adj_21_LC_4_25_3 .C_ON=1'b0;
    defparam \nx.i3_3_lut_adj_21_LC_4_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.i3_3_lut_adj_21_LC_4_25_3 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \nx.i3_3_lut_adj_21_LC_4_25_3  (
            .in0(_gnd_net_),
            .in1(N__23866),
            .in2(N__22260),
            .in3(N__22174),
            .lcout(),
            .ltout(\nx.n15_adj_676_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_LC_4_25_4 .C_ON=1'b0;
    defparam \nx.i10_4_lut_LC_4_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_LC_4_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_LC_4_25_4  (
            .in0(N__22555),
            .in1(N__22416),
            .in2(N__20391),
            .in3(N__20817),
            .lcout(\nx.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_135_LC_4_25_5 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_135_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_135_LC_4_25_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_135_LC_4_25_5  (
            .in0(N__30146),
            .in1(N__24052),
            .in2(N__25332),
            .in3(N__28213),
            .lcout(\nx.n47_adj_780 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_2_lut_LC_4_25_6 .C_ON=1'b0;
    defparam \nx.i6_2_lut_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.i6_2_lut_LC_4_25_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i6_2_lut_LC_4_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22512),
            .in3(N__22576),
            .lcout(\nx.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_adj_159_LC_4_25_7.C_ON=1'b0;
    defparam i8_4_lut_adj_159_LC_4_25_7.SEQ_MODE=4'b0000;
    defparam i8_4_lut_adj_159_LC_4_25_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i8_4_lut_adj_159_LC_4_25_7 (
            .in0(N__20793),
            .in1(N__20778),
            .in2(N__20763),
            .in3(N__20742),
            .lcout(n19_adj_814),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_2_lut_LC_4_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_2_lut_LC_4_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_2_lut_LC_4_26_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1071_2_lut_LC_4_26_0  (
            .in0(N__23828),
            .in1(N__23827),
            .in2(N__20711),
            .in3(N__20727),
            .lcout(\nx.n1609 ),
            .ltout(),
            .carryin(bfn_4_26_0_),
            .carryout(\nx.n10783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_3_lut_LC_4_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_3_lut_LC_4_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_3_lut_LC_4_26_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1071_3_lut_LC_4_26_1  (
            .in0(N__20724),
            .in1(N__20723),
            .in2(N__20712),
            .in3(N__20694),
            .lcout(\nx.n1608 ),
            .ltout(),
            .carryin(\nx.n10783 ),
            .carryout(\nx.n10784 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_4_lut_LC_4_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_4_lut_LC_4_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_4_lut_LC_4_26_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_4_lut_LC_4_26_2  (
            .in0(N__20691),
            .in1(N__20690),
            .in2(N__20889),
            .in3(N__20673),
            .lcout(\nx.n1607 ),
            .ltout(),
            .carryin(\nx.n10784 ),
            .carryout(\nx.n10785 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_5_lut_LC_4_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_5_lut_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_5_lut_LC_4_26_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_5_lut_LC_4_26_3  (
            .in0(N__20670),
            .in1(N__20669),
            .in2(N__20892),
            .in3(N__20658),
            .lcout(\nx.n1606 ),
            .ltout(),
            .carryin(\nx.n10785 ),
            .carryout(\nx.n10786 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_6_lut_LC_4_26_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_6_lut_LC_4_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_6_lut_LC_4_26_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_6_lut_LC_4_26_4  (
            .in0(N__20655),
            .in1(N__20654),
            .in2(N__20890),
            .in3(N__20637),
            .lcout(\nx.n1605 ),
            .ltout(),
            .carryin(\nx.n10786 ),
            .carryout(\nx.n10787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_7_lut_LC_4_26_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_7_lut_LC_4_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_7_lut_LC_4_26_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_7_lut_LC_4_26_5  (
            .in0(N__20634),
            .in1(N__20633),
            .in2(N__20893),
            .in3(N__20616),
            .lcout(\nx.n1604 ),
            .ltout(),
            .carryin(\nx.n10787 ),
            .carryout(\nx.n10788 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_8_lut_LC_4_26_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_8_lut_LC_4_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_8_lut_LC_4_26_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_8_lut_LC_4_26_6  (
            .in0(N__21030),
            .in1(N__21029),
            .in2(N__20891),
            .in3(N__21012),
            .lcout(\nx.n1603 ),
            .ltout(),
            .carryin(\nx.n10788 ),
            .carryout(\nx.n10789 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_9_lut_LC_4_26_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_9_lut_LC_4_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_9_lut_LC_4_26_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_9_lut_LC_4_26_7  (
            .in0(N__21009),
            .in1(N__21008),
            .in2(N__20894),
            .in3(N__20991),
            .lcout(\nx.n1602 ),
            .ltout(),
            .carryin(\nx.n10789 ),
            .carryout(\nx.n10790 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_10_lut_LC_4_27_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_10_lut_LC_4_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_10_lut_LC_4_27_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_10_lut_LC_4_27_0  (
            .in0(N__20988),
            .in1(N__20987),
            .in2(N__20895),
            .in3(N__20973),
            .lcout(\nx.n1601 ),
            .ltout(),
            .carryin(bfn_4_27_0_),
            .carryout(\nx.n10791 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_11_lut_LC_4_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_11_lut_LC_4_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_11_lut_LC_4_27_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_11_lut_LC_4_27_1  (
            .in0(N__20970),
            .in1(N__20969),
            .in2(N__20897),
            .in3(N__20946),
            .lcout(\nx.n1600 ),
            .ltout(),
            .carryin(\nx.n10791 ),
            .carryout(\nx.n10792 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_12_lut_LC_4_27_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1071_12_lut_LC_4_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_12_lut_LC_4_27_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_12_lut_LC_4_27_2  (
            .in0(N__20942),
            .in1(N__20943),
            .in2(N__20896),
            .in3(N__20925),
            .lcout(\nx.n1599 ),
            .ltout(),
            .carryin(\nx.n10792 ),
            .carryout(\nx.n10793 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1071_13_lut_LC_4_27_3 .C_ON=1'b0;
    defparam \nx.mod_5_add_1071_13_lut_LC_4_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1071_13_lut_LC_4_27_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1071_13_lut_LC_4_27_3  (
            .in0(N__20922),
            .in1(N__20921),
            .in2(N__20898),
            .in3(N__20826),
            .lcout(\nx.n1598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_136_LC_4_27_5 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_136_LC_4_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_136_LC_4_27_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_136_LC_4_27_5  (
            .in0(N__28936),
            .in1(N__23952),
            .in2(N__26034),
            .in3(N__34340),
            .lcout(\nx.n45_adj_781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_4_lut_adj_22_LC_4_27_7 .C_ON=1'b0;
    defparam \nx.i7_4_lut_adj_22_LC_4_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.i7_4_lut_adj_22_LC_4_27_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i7_4_lut_adj_22_LC_4_27_7  (
            .in0(N__22195),
            .in1(N__22483),
            .in2(N__22462),
            .in3(N__22435),
            .lcout(\nx.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_0__bdd_4_lut_LC_5_14_7.C_ON=1'b0;
    defparam current_pin_0__bdd_4_lut_LC_5_14_7.SEQ_MODE=4'b0000;
    defparam current_pin_0__bdd_4_lut_LC_5_14_7.LUT_INIT=16'b1111001110001000;
    LogicCell40 current_pin_0__bdd_4_lut_LC_5_14_7 (
            .in0(N__21234),
            .in1(N__46545),
            .in2(N__21216),
            .in3(N__46405),
            .lcout(n13649),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i6_LC_5_15_0.C_ON=1'b0;
    defparam pin_output_enable__i6_LC_5_15_0.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i6_LC_5_15_0.LUT_INIT=16'b1101100011001100;
    LogicCell40 pin_output_enable__i6_LC_5_15_0 (
            .in0(N__22893),
            .in1(N__21176),
            .in2(N__47675),
            .in3(N__47121),
            .lcout(pin_oe_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46861),
            .ce(),
            .sr(_gnd_net_));
    defparam n13649_bdd_4_lut_LC_5_15_1.C_ON=1'b0;
    defparam n13649_bdd_4_lut_LC_5_15_1.SEQ_MODE=4'b0000;
    defparam n13649_bdd_4_lut_LC_5_15_1.LUT_INIT=16'b1110111000110000;
    LogicCell40 n13649_bdd_4_lut_LC_5_15_1 (
            .in0(N__21165),
            .in1(N__46566),
            .in2(N__21147),
            .in3(N__21126),
            .lcout(n13652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i30_LC_5_16_3 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i30_LC_5_16_3 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i30_LC_5_16_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i30_LC_5_16_3  (
            .in0(N__21120),
            .in1(N__21090),
            .in2(_gnd_net_),
            .in3(N__25157),
            .lcout(neo_pixel_transmitter_t0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46855),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7610_4_lut_LC_5_17_0 .C_ON=1'b0;
    defparam \nx.i7610_4_lut_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.i7610_4_lut_LC_5_17_0 .LUT_INIT=16'b1111111111001010;
    LogicCell40 \nx.i7610_4_lut_LC_5_17_0  (
            .in0(N__23203),
            .in1(N__22855),
            .in2(N__26805),
            .in3(N__23183),
            .lcout(\nx.n11946 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i53_4_lut_LC_5_17_2 .C_ON=1'b0;
    defparam \nx.i53_4_lut_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \nx.i53_4_lut_LC_5_17_2 .LUT_INIT=16'b1100110011111010;
    LogicCell40 \nx.i53_4_lut_LC_5_17_2  (
            .in0(N__21072),
            .in1(N__21268),
            .in2(N__23187),
            .in3(N__23481),
            .lcout(),
            .ltout(\nx.n11948_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i52_4_lut_LC_5_17_3 .C_ON=1'b0;
    defparam \nx.i52_4_lut_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.i52_4_lut_LC_5_17_3 .LUT_INIT=16'b0000000111101111;
    LogicCell40 \nx.i52_4_lut_LC_5_17_3  (
            .in0(N__24943),
            .in1(N__26795),
            .in2(N__21066),
            .in3(N__22887),
            .lcout(\nx.n11988 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8984_3_lut_LC_5_17_4.C_ON=1'b0;
    defparam i8984_3_lut_LC_5_17_4.SEQ_MODE=4'b0000;
    defparam i8984_3_lut_LC_5_17_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i8984_3_lut_LC_5_17_4 (
            .in0(N__21063),
            .in1(N__21048),
            .in2(_gnd_net_),
            .in3(N__46396),
            .lcout(),
            .ltout(n13379_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13613_bdd_4_lut_LC_5_17_5.C_ON=1'b0;
    defparam n13613_bdd_4_lut_LC_5_17_5.SEQ_MODE=4'b0000;
    defparam n13613_bdd_4_lut_LC_5_17_5.LUT_INIT=16'b1111110000100010;
    LogicCell40 n13613_bdd_4_lut_LC_5_17_5 (
            .in0(N__21507),
            .in1(N__45645),
            .in2(N__21033),
            .in3(N__21447),
            .lcout(n13616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_4_lut_4_lut_LC_5_17_6 .C_ON=1'b0;
    defparam \nx.i3_4_lut_4_lut_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.i3_4_lut_4_lut_LC_5_17_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \nx.i3_4_lut_4_lut_LC_5_17_6  (
            .in0(N__26796),
            .in1(N__23482),
            .in2(N__21276),
            .in3(N__24944),
            .lcout(\nx.n12451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9091_2_lut_LC_5_17_7 .C_ON=1'b0;
    defparam \nx.i9091_2_lut_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \nx.i9091_2_lut_LC_5_17_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \nx.i9091_2_lut_LC_5_17_7  (
            .in0(N__24942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26794),
            .lcout(\nx.n13438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i15_LC_5_18_0.C_ON=1'b0;
    defparam neopxl_color_i15_LC_5_18_0.SEQ_MODE=4'b1000;
    defparam neopxl_color_i15_LC_5_18_0.LUT_INIT=16'b1111011100010000;
    LogicCell40 neopxl_color_i15_LC_5_18_0 (
            .in0(N__47673),
            .in1(N__43939),
            .in2(N__43701),
            .in3(N__25757),
            .lcout(neopxl_color_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46856),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_145_LC_5_18_1 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_145_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_145_LC_5_18_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \nx.i1_2_lut_adj_145_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(N__21331),
            .in2(_gnd_net_),
            .in3(N__21383),
            .lcout(\nx.n11908 ),
            .ltout(\nx.n11908_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7592_4_lut_LC_5_18_2 .C_ON=1'b0;
    defparam \nx.i7592_4_lut_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.i7592_4_lut_LC_5_18_2 .LUT_INIT=16'b1111111111100100;
    LogicCell40 \nx.i7592_4_lut_LC_5_18_2  (
            .in0(N__26802),
            .in1(N__22854),
            .in2(N__21351),
            .in3(N__23168),
            .lcout(\nx.n11926 ),
            .ltout(\nx.n11926_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_127_LC_5_18_3 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_127_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_127_LC_5_18_3 .LUT_INIT=16'b1011101000000000;
    LogicCell40 \nx.i1_4_lut_adj_127_LC_5_18_3  (
            .in0(N__23472),
            .in1(N__22868),
            .in2(N__21339),
            .in3(N__21240),
            .lcout(n7671),
            .ltout(n7671_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.state_i1_LC_5_18_4 .C_ON=1'b0;
    defparam \nx.state_i1_LC_5_18_4 .SEQ_MODE=4'b1000;
    defparam \nx.state_i1_LC_5_18_4 .LUT_INIT=16'b1101111111110000;
    LogicCell40 \nx.state_i1_LC_5_18_4  (
            .in0(N__26803),
            .in1(N__26855),
            .in2(N__21336),
            .in3(N__23473),
            .lcout(state_1_adj_791),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46856),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2_2_lut_adj_146_LC_5_18_5 .C_ON=1'b0;
    defparam \nx.i2_2_lut_adj_146_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.i2_2_lut_adj_146_LC_5_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \nx.i2_2_lut_adj_146_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(N__21332),
            .in2(_gnd_net_),
            .in3(N__21297),
            .lcout(\nx.n11113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_3_lut_4_lut_LC_5_18_6 .C_ON=1'b0;
    defparam \nx.i1_3_lut_4_lut_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.i1_3_lut_4_lut_LC_5_18_6 .LUT_INIT=16'b1011111110111011;
    LogicCell40 \nx.i1_3_lut_4_lut_LC_5_18_6  (
            .in0(N__26801),
            .in1(N__23471),
            .in2(N__24957),
            .in3(N__21258),
            .lcout(\nx.n12381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i11_LC_5_18_7 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i11_LC_5_18_7 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i11_LC_5_18_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i11_LC_5_18_7  (
            .in0(N__21564),
            .in1(N__21438),
            .in2(_gnd_net_),
            .in3(N__25155),
            .lcout(neo_pixel_transmitter_t0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46856),
            .ce(),
            .sr(_gnd_net_));
    defparam i8983_3_lut_LC_5_19_0.C_ON=1'b0;
    defparam i8983_3_lut_LC_5_19_0.SEQ_MODE=4'b0000;
    defparam i8983_3_lut_LC_5_19_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 i8983_3_lut_LC_5_19_0 (
            .in0(N__21537),
            .in1(N__21522),
            .in2(_gnd_net_),
            .in3(N__46407),
            .lcout(n13378),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8986_3_lut_LC_5_19_2.C_ON=1'b0;
    defparam i8986_3_lut_LC_5_19_2.SEQ_MODE=4'b0000;
    defparam i8986_3_lut_LC_5_19_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 i8986_3_lut_LC_5_19_2 (
            .in0(N__21498),
            .in1(N__21477),
            .in2(_gnd_net_),
            .in3(N__46406),
            .lcout(),
            .ltout(n13381_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_1__bdd_4_lut_9226_LC_5_19_3.C_ON=1'b0;
    defparam current_pin_1__bdd_4_lut_9226_LC_5_19_3.SEQ_MODE=4'b0000;
    defparam current_pin_1__bdd_4_lut_9226_LC_5_19_3.LUT_INIT=16'b1101110110100000;
    LogicCell40 current_pin_1__bdd_4_lut_9226_LC_5_19_3 (
            .in0(N__45644),
            .in1(N__21456),
            .in2(N__21450),
            .in3(N__46565),
            .lcout(n13613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i12_1_lut_LC_5_19_7 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i12_1_lut_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i12_1_lut_LC_5_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i12_1_lut_LC_5_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21437),
            .lcout(\nx.n22_adj_749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i739_3_lut_LC_5_20_0 .C_ON=1'b0;
    defparam \nx.mod_5_i739_3_lut_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i739_3_lut_LC_5_20_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i739_3_lut_LC_5_20_0  (
            .in0(N__23553),
            .in1(_gnd_net_),
            .in2(N__23604),
            .in3(N__23361),
            .lcout(\nx.n1104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i743_3_lut_LC_5_20_1 .C_ON=1'b0;
    defparam \nx.mod_5_i743_3_lut_LC_5_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i743_3_lut_LC_5_20_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i743_3_lut_LC_5_20_1  (
            .in0(_gnd_net_),
            .in1(N__23582),
            .in2(N__23388),
            .in3(N__23552),
            .lcout(\nx.n1108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i20_1_lut_LC_5_20_2 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i20_1_lut_LC_5_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i20_1_lut_LC_5_20_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \nx.sub_14_inv_0_i20_1_lut_LC_5_20_2  (
            .in0(N__21413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\nx.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i741_3_lut_LC_5_20_3 .C_ON=1'b0;
    defparam \nx.mod_5_i741_3_lut_LC_5_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i741_3_lut_LC_5_20_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i741_3_lut_LC_5_20_3  (
            .in0(_gnd_net_),
            .in1(N__23548),
            .in2(N__23652),
            .in3(N__23373),
            .lcout(\nx.n1106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i744_3_lut_LC_5_20_4 .C_ON=1'b0;
    defparam \nx.mod_5_i744_3_lut_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i744_3_lut_LC_5_20_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i744_3_lut_LC_5_20_4  (
            .in0(_gnd_net_),
            .in1(N__23397),
            .in2(N__23558),
            .in3(N__23951),
            .lcout(\nx.n1109 ),
            .ltout(\nx.n1109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5944_2_lut_LC_5_20_5 .C_ON=1'b0;
    defparam \nx.i5944_2_lut_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.i5944_2_lut_LC_5_20_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \nx.i5944_2_lut_LC_5_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21654),
            .in3(N__23998),
            .lcout(),
            .ltout(\nx.n9737_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_4_lut_LC_5_20_6 .C_ON=1'b0;
    defparam \nx.i5_4_lut_LC_5_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.i5_4_lut_LC_5_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i5_4_lut_LC_5_20_6  (
            .in0(N__21601),
            .in1(N__21895),
            .in2(N__21651),
            .in3(N__23509),
            .lcout(),
            .ltout(\nx.n12_adj_673_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_4_lut_LC_5_20_7 .C_ON=1'b0;
    defparam \nx.i6_4_lut_LC_5_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.i6_4_lut_LC_5_20_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i6_4_lut_LC_5_20_7  (
            .in0(N__23623),
            .in1(N__23348),
            .in2(N__21648),
            .in3(N__21853),
            .lcout(\nx.n1136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_2_lut_LC_5_21_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_2_lut_LC_5_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_2_lut_LC_5_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_2_lut_LC_5_21_0  (
            .in0(_gnd_net_),
            .in1(N__23999),
            .in2(_gnd_net_),
            .in3(N__21636),
            .lcout(\nx.n1177 ),
            .ltout(),
            .carryin(bfn_5_21_0_),
            .carryout(\nx.n10749 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_3_lut_LC_5_21_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_3_lut_LC_5_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_3_lut_LC_5_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_3_lut_LC_5_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21633),
            .in3(N__21609),
            .lcout(\nx.n1176 ),
            .ltout(),
            .carryin(\nx.n10749 ),
            .carryout(\nx.n10750 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_4_lut_LC_5_21_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_4_lut_LC_5_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_4_lut_LC_5_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_4_lut_LC_5_21_2  (
            .in0(_gnd_net_),
            .in1(N__42219),
            .in2(N__21606),
            .in3(N__21579),
            .lcout(\nx.n1175 ),
            .ltout(),
            .carryin(\nx.n10750 ),
            .carryout(\nx.n10751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_5_lut_LC_5_21_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_5_lut_LC_5_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_5_lut_LC_5_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_5_lut_LC_5_21_3  (
            .in0(_gnd_net_),
            .in1(N__42193),
            .in2(N__23627),
            .in3(N__21567),
            .lcout(\nx.n1174 ),
            .ltout(),
            .carryin(\nx.n10751 ),
            .carryout(\nx.n10752 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_6_lut_LC_5_21_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_6_lut_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_6_lut_LC_5_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_6_lut_LC_5_21_4  (
            .in0(_gnd_net_),
            .in1(N__42220),
            .in2(N__21900),
            .in3(N__21873),
            .lcout(\nx.n1173 ),
            .ltout(),
            .carryin(\nx.n10752 ),
            .carryout(\nx.n10753 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_7_lut_LC_5_21_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_7_lut_LC_5_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_7_lut_LC_5_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_7_lut_LC_5_21_5  (
            .in0(_gnd_net_),
            .in1(N__42194),
            .in2(N__23516),
            .in3(N__21864),
            .lcout(\nx.n1172 ),
            .ltout(),
            .carryin(\nx.n10753 ),
            .carryout(\nx.n10754 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_8_lut_LC_5_21_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_803_8_lut_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_8_lut_LC_5_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_803_8_lut_LC_5_21_6  (
            .in0(_gnd_net_),
            .in1(N__42221),
            .in2(N__21860),
            .in3(N__21831),
            .lcout(\nx.n1171 ),
            .ltout(),
            .carryin(\nx.n10754 ),
            .carryout(\nx.n10755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_803_9_lut_LC_5_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_add_803_9_lut_LC_5_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_803_9_lut_LC_5_21_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_803_9_lut_LC_5_21_7  (
            .in0(N__42222),
            .in1(N__21820),
            .in2(N__23349),
            .in3(N__21780),
            .lcout(\nx.n1202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_2_lut_LC_5_22_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_2_lut_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_2_lut_LC_5_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_2_lut_LC_5_22_0  (
            .in0(_gnd_net_),
            .in1(N__24048),
            .in2(_gnd_net_),
            .in3(N__21765),
            .lcout(\nx.n1277 ),
            .ltout(),
            .carryin(bfn_5_22_0_),
            .carryout(\nx.n10756 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_3_lut_LC_5_22_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_3_lut_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_3_lut_LC_5_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_3_lut_LC_5_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21762),
            .in3(N__21729),
            .lcout(\nx.n1276 ),
            .ltout(),
            .carryin(\nx.n10756 ),
            .carryout(\nx.n10757 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_4_lut_LC_5_22_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_4_lut_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_4_lut_LC_5_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_4_lut_LC_5_22_2  (
            .in0(_gnd_net_),
            .in1(N__42096),
            .in2(N__21726),
            .in3(N__21702),
            .lcout(\nx.n1275 ),
            .ltout(),
            .carryin(\nx.n10757 ),
            .carryout(\nx.n10758 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_5_lut_LC_5_22_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_5_lut_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_5_lut_LC_5_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_5_lut_LC_5_22_3  (
            .in0(_gnd_net_),
            .in1(N__42195),
            .in2(N__21699),
            .in3(N__21675),
            .lcout(\nx.n1274 ),
            .ltout(),
            .carryin(\nx.n10758 ),
            .carryout(\nx.n10759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_6_lut_LC_5_22_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_6_lut_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_6_lut_LC_5_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_6_lut_LC_5_22_4  (
            .in0(_gnd_net_),
            .in1(N__42097),
            .in2(N__21672),
            .in3(N__22146),
            .lcout(\nx.n1273 ),
            .ltout(),
            .carryin(\nx.n10759 ),
            .carryout(\nx.n10760 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_7_lut_LC_5_22_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_7_lut_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_7_lut_LC_5_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_7_lut_LC_5_22_5  (
            .in0(_gnd_net_),
            .in1(N__42196),
            .in2(N__22143),
            .in3(N__22122),
            .lcout(\nx.n1272 ),
            .ltout(),
            .carryin(\nx.n10760 ),
            .carryout(\nx.n10761 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_8_lut_LC_5_22_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_8_lut_LC_5_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_8_lut_LC_5_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_8_lut_LC_5_22_6  (
            .in0(_gnd_net_),
            .in1(N__42098),
            .in2(N__22118),
            .in3(N__22086),
            .lcout(\nx.n1271 ),
            .ltout(),
            .carryin(\nx.n10761 ),
            .carryout(\nx.n10762 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_9_lut_LC_5_22_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_870_9_lut_LC_5_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_9_lut_LC_5_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_870_9_lut_LC_5_22_7  (
            .in0(_gnd_net_),
            .in1(N__42197),
            .in2(N__21999),
            .in3(N__22083),
            .lcout(\nx.n1270 ),
            .ltout(),
            .carryin(\nx.n10762 ),
            .carryout(\nx.n10763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_870_10_lut_LC_5_23_0 .C_ON=1'b0;
    defparam \nx.mod_5_add_870_10_lut_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_870_10_lut_LC_5_23_0 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_870_10_lut_LC_5_23_0  (
            .in0(N__42198),
            .in1(N__21972),
            .in2(N__22080),
            .in3(N__22062),
            .lcout(\nx.n1301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_157_LC_5_23_5.C_ON=1'b0;
    defparam i1_2_lut_adj_157_LC_5_23_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_157_LC_5_23_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_157_LC_5_23_5 (
            .in0(_gnd_net_),
            .in1(N__22044),
            .in2(_gnd_net_),
            .in3(N__22026),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i873_3_lut_LC_5_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i873_3_lut_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i873_3_lut_LC_5_23_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i873_3_lut_LC_5_23_7  (
            .in0(_gnd_net_),
            .in1(N__21998),
            .in2(N__21982),
            .in3(N__21936),
            .lcout(\nx.n1302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i21_4_lut_adj_140_LC_5_24_1 .C_ON=1'b0;
    defparam \nx.i21_4_lut_adj_140_LC_5_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.i21_4_lut_adj_140_LC_5_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i21_4_lut_adj_140_LC_5_24_1  (
            .in0(N__31778),
            .in1(N__23864),
            .in2(N__26082),
            .in3(N__38912),
            .lcout(),
            .ltout(\nx.n49_adj_784_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i27_4_lut_LC_5_24_2 .C_ON=1'b0;
    defparam \nx.i27_4_lut_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.i27_4_lut_LC_5_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i27_4_lut_LC_5_24_2  (
            .in0(N__25434),
            .in1(N__22269),
            .in2(N__21915),
            .in3(N__21912),
            .lcout(state_3_N_448_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9167_2_lut_3_lut_LC_5_24_4.C_ON=1'b0;
    defparam i9167_2_lut_3_lut_LC_5_24_4.SEQ_MODE=4'b0000;
    defparam i9167_2_lut_3_lut_LC_5_24_4.LUT_INIT=16'b0100010000000000;
    LogicCell40 i9167_2_lut_3_lut_LC_5_24_4 (
            .in0(N__43652),
            .in1(N__43947),
            .in2(_gnd_net_),
            .in3(N__47664),
            .lcout(n7664),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2_2_lut_adj_132_LC_5_24_5 .C_ON=1'b0;
    defparam \nx.i2_2_lut_adj_132_LC_5_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.i2_2_lut_adj_132_LC_5_24_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \nx.i2_2_lut_adj_132_LC_5_24_5  (
            .in0(N__26353),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25899),
            .lcout(),
            .ltout(\nx.n30_adj_777_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_138_LC_5_24_6 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_138_LC_5_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_138_LC_5_24_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \nx.i15_4_lut_adj_138_LC_5_24_6  (
            .in0(N__30791),
            .in1(N__32391),
            .in2(N__22272),
            .in3(N__23997),
            .lcout(\nx.n43_adj_783 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_2_lut_LC_5_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_2_lut_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_2_lut_LC_5_25_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1138_2_lut_LC_5_25_0  (
            .in0(N__23868),
            .in1(N__23867),
            .in2(N__22238),
            .in3(N__22263),
            .lcout(\nx.n1709 ),
            .ltout(),
            .carryin(bfn_5_25_0_),
            .carryout(\nx.n10794 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_3_lut_LC_5_25_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_3_lut_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_3_lut_LC_5_25_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1138_3_lut_LC_5_25_1  (
            .in0(N__22259),
            .in1(N__22258),
            .in2(N__22239),
            .in3(N__22221),
            .lcout(\nx.n1708 ),
            .ltout(),
            .carryin(\nx.n10794 ),
            .carryout(\nx.n10795 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_4_lut_LC_5_25_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_4_lut_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_4_lut_LC_5_25_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_4_lut_LC_5_25_2  (
            .in0(N__22218),
            .in1(N__22217),
            .in2(N__22385),
            .in3(N__22200),
            .lcout(\nx.n1707 ),
            .ltout(),
            .carryin(\nx.n10795 ),
            .carryout(\nx.n10796 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_5_lut_LC_5_25_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_5_lut_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_5_lut_LC_5_25_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_5_lut_LC_5_25_3  (
            .in0(N__22197),
            .in1(N__22196),
            .in2(N__22388),
            .in3(N__22179),
            .lcout(\nx.n1706 ),
            .ltout(),
            .carryin(\nx.n10796 ),
            .carryout(\nx.n10797 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_6_lut_LC_5_25_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_6_lut_LC_5_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_6_lut_LC_5_25_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_6_lut_LC_5_25_4  (
            .in0(N__22176),
            .in1(N__22175),
            .in2(N__22386),
            .in3(N__22158),
            .lcout(\nx.n1705 ),
            .ltout(),
            .carryin(\nx.n10797 ),
            .carryout(\nx.n10798 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_7_lut_LC_5_25_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_7_lut_LC_5_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_7_lut_LC_5_25_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_7_lut_LC_5_25_5  (
            .in0(N__22578),
            .in1(N__22577),
            .in2(N__22389),
            .in3(N__22560),
            .lcout(\nx.n1704 ),
            .ltout(),
            .carryin(\nx.n10798 ),
            .carryout(\nx.n10799 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_8_lut_LC_5_25_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_8_lut_LC_5_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_8_lut_LC_5_25_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_8_lut_LC_5_25_6  (
            .in0(N__22557),
            .in1(N__22556),
            .in2(N__22387),
            .in3(N__22539),
            .lcout(\nx.n1703 ),
            .ltout(),
            .carryin(\nx.n10799 ),
            .carryout(\nx.n10800 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_9_lut_LC_5_25_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_9_lut_LC_5_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_9_lut_LC_5_25_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_9_lut_LC_5_25_7  (
            .in0(N__22535),
            .in1(N__22534),
            .in2(N__22390),
            .in3(N__22515),
            .lcout(\nx.n1702 ),
            .ltout(),
            .carryin(\nx.n10800 ),
            .carryout(\nx.n10801 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_10_lut_LC_5_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_10_lut_LC_5_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_10_lut_LC_5_26_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_10_lut_LC_5_26_0  (
            .in0(N__22511),
            .in1(N__22510),
            .in2(N__22391),
            .in3(N__22491),
            .lcout(\nx.n1701 ),
            .ltout(),
            .carryin(bfn_5_26_0_),
            .carryout(\nx.n10802 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_11_lut_LC_5_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_11_lut_LC_5_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_11_lut_LC_5_26_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_11_lut_LC_5_26_1  (
            .in0(N__22487),
            .in1(N__22488),
            .in2(N__22394),
            .in3(N__22467),
            .lcout(\nx.n1700 ),
            .ltout(),
            .carryin(\nx.n10802 ),
            .carryout(\nx.n10803 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_12_lut_LC_5_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_12_lut_LC_5_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_12_lut_LC_5_26_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_12_lut_LC_5_26_2  (
            .in0(N__22464),
            .in1(N__22463),
            .in2(N__22392),
            .in3(N__22440),
            .lcout(\nx.n1699 ),
            .ltout(),
            .carryin(\nx.n10803 ),
            .carryout(\nx.n10804 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_13_lut_LC_5_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1138_13_lut_LC_5_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_13_lut_LC_5_26_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_13_lut_LC_5_26_3  (
            .in0(N__22437),
            .in1(N__22436),
            .in2(N__22395),
            .in3(N__22419),
            .lcout(\nx.n1698 ),
            .ltout(),
            .carryin(\nx.n10804 ),
            .carryout(\nx.n10805 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1138_14_lut_LC_5_26_4 .C_ON=1'b0;
    defparam \nx.mod_5_add_1138_14_lut_LC_5_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1138_14_lut_LC_5_26_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1138_14_lut_LC_5_26_4  (
            .in0(N__22414),
            .in1(N__22415),
            .in2(N__22393),
            .in3(N__22317),
            .lcout(\nx.n1697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_3_lut_adj_130_LC_5_26_5 .C_ON=1'b0;
    defparam \nx.i7_3_lut_adj_130_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.i7_3_lut_adj_130_LC_5_26_5 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \nx.i7_3_lut_adj_130_LC_5_26_5  (
            .in0(_gnd_net_),
            .in1(N__22654),
            .in2(N__22606),
            .in3(N__22822),
            .lcout(\nx.n20_adj_775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_3_lut_adj_119_LC_5_26_7 .C_ON=1'b0;
    defparam \nx.i3_3_lut_adj_119_LC_5_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.i3_3_lut_adj_119_LC_5_26_7 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \nx.i3_3_lut_adj_119_LC_5_26_7  (
            .in0(N__24743),
            .in1(_gnd_net_),
            .in2(N__22690),
            .in3(N__22630),
            .lcout(\nx.n16_adj_766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_2_lut_LC_5_27_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_2_lut_LC_5_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_2_lut_LC_5_27_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1205_2_lut_LC_5_27_0  (
            .in0(N__24764),
            .in1(N__24763),
            .in2(N__22913),
            .in3(N__22695),
            .lcout(\nx.n1809 ),
            .ltout(),
            .carryin(bfn_5_27_0_),
            .carryout(\nx.n10806 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_3_lut_LC_5_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_3_lut_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_3_lut_LC_5_27_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1205_3_lut_LC_5_27_1  (
            .in0(N__22692),
            .in1(N__22691),
            .in2(N__22914),
            .in3(N__22668),
            .lcout(\nx.n1808 ),
            .ltout(),
            .carryin(\nx.n10806 ),
            .carryout(\nx.n10807 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_4_lut_LC_5_27_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_4_lut_LC_5_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_4_lut_LC_5_27_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_4_lut_LC_5_27_2  (
            .in0(N__22665),
            .in1(N__22661),
            .in2(N__22999),
            .in3(N__22641),
            .lcout(\nx.n1807 ),
            .ltout(),
            .carryin(\nx.n10807 ),
            .carryout(\nx.n10808 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_5_lut_LC_5_27_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_5_lut_LC_5_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_5_lut_LC_5_27_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_5_lut_LC_5_27_3  (
            .in0(N__22638),
            .in1(N__22637),
            .in2(N__23002),
            .in3(N__22617),
            .lcout(\nx.n1806 ),
            .ltout(),
            .carryin(\nx.n10808 ),
            .carryout(\nx.n10809 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_6_lut_LC_5_27_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_6_lut_LC_5_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_6_lut_LC_5_27_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_6_lut_LC_5_27_4  (
            .in0(N__22764),
            .in1(N__22763),
            .in2(N__23000),
            .in3(N__22614),
            .lcout(\nx.n1805 ),
            .ltout(),
            .carryin(\nx.n10809 ),
            .carryout(\nx.n10810 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_7_lut_LC_5_27_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_7_lut_LC_5_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_7_lut_LC_5_27_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_7_lut_LC_5_27_5  (
            .in0(N__22742),
            .in1(N__22741),
            .in2(N__23003),
            .in3(N__22611),
            .lcout(\nx.n1804 ),
            .ltout(),
            .carryin(\nx.n10810 ),
            .carryout(\nx.n10811 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_8_lut_LC_5_27_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_8_lut_LC_5_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_8_lut_LC_5_27_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_8_lut_LC_5_27_6  (
            .in0(N__22608),
            .in1(N__22607),
            .in2(N__23001),
            .in3(N__22584),
            .lcout(\nx.n1803 ),
            .ltout(),
            .carryin(\nx.n10811 ),
            .carryout(\nx.n10812 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_9_lut_LC_5_27_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_9_lut_LC_5_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_9_lut_LC_5_27_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_9_lut_LC_5_27_7  (
            .in0(N__22794),
            .in1(N__22787),
            .in2(N__23004),
            .in3(N__22581),
            .lcout(\nx.n1802 ),
            .ltout(),
            .carryin(\nx.n10812 ),
            .carryout(\nx.n10813 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_10_lut_LC_5_28_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_10_lut_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_10_lut_LC_5_28_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_10_lut_LC_5_28_0  (
            .in0(N__23112),
            .in1(N__23111),
            .in2(N__22993),
            .in3(N__22833),
            .lcout(\nx.n1801 ),
            .ltout(),
            .carryin(bfn_5_28_0_),
            .carryout(\nx.n10814 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_11_lut_LC_5_28_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_11_lut_LC_5_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_11_lut_LC_5_28_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_11_lut_LC_5_28_1  (
            .in0(N__22830),
            .in1(N__22829),
            .in2(N__22996),
            .in3(N__22809),
            .lcout(\nx.n1800 ),
            .ltout(),
            .carryin(\nx.n10814 ),
            .carryout(\nx.n10815 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_12_lut_LC_5_28_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_12_lut_LC_5_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_12_lut_LC_5_28_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_12_lut_LC_5_28_2  (
            .in0(N__22716),
            .in1(N__22715),
            .in2(N__22994),
            .in3(N__22806),
            .lcout(\nx.n1799 ),
            .ltout(),
            .carryin(\nx.n10815 ),
            .carryout(\nx.n10816 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_13_lut_LC_5_28_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_13_lut_LC_5_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_13_lut_LC_5_28_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_13_lut_LC_5_28_3  (
            .in0(N__23064),
            .in1(N__23063),
            .in2(N__22997),
            .in3(N__22803),
            .lcout(\nx.n1798 ),
            .ltout(),
            .carryin(\nx.n10816 ),
            .carryout(\nx.n10817 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_14_lut_LC_5_28_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1205_14_lut_LC_5_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_14_lut_LC_5_28_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_14_lut_LC_5_28_4  (
            .in0(N__23088),
            .in1(N__23087),
            .in2(N__22995),
            .in3(N__22800),
            .lcout(\nx.n1797 ),
            .ltout(),
            .carryin(\nx.n10817 ),
            .carryout(\nx.n10818 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1205_15_lut_LC_5_28_5 .C_ON=1'b0;
    defparam \nx.mod_5_add_1205_15_lut_LC_5_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1205_15_lut_LC_5_28_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1205_15_lut_LC_5_28_5  (
            .in0(N__23042),
            .in1(N__23043),
            .in2(N__22998),
            .in3(N__22797),
            .lcout(\nx.n1796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_2_lut_LC_5_28_6 .C_ON=1'b0;
    defparam \nx.i4_2_lut_LC_5_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.i4_2_lut_LC_5_28_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i4_2_lut_LC_5_28_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24138),
            .in3(N__24157),
            .lcout(\nx.n18_adj_716 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_129_LC_5_29_1 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_129_LC_5_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_129_LC_5_29_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_adj_129_LC_5_29_1  (
            .in0(N__22786),
            .in1(N__22762),
            .in2(N__22743),
            .in3(N__22714),
            .lcout(),
            .ltout(\nx.n22_adj_774_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_131_LC_5_29_2 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_131_LC_5_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_131_LC_5_29_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_131_LC_5_29_2  (
            .in0(N__23121),
            .in1(N__23110),
            .in2(N__23091),
            .in3(N__23086),
            .lcout(),
            .ltout(\nx.n24_adj_776_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_143_LC_5_29_3 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_143_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_143_LC_5_29_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_143_LC_5_29_3  (
            .in0(N__23062),
            .in1(N__23041),
            .in2(N__23016),
            .in3(N__23013),
            .lcout(\nx.n1730 ),
            .ltout(\nx.n1730_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9205_1_lut_LC_5_29_4 .C_ON=1'b0;
    defparam \nx.i9205_1_lut_LC_5_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.i9205_1_lut_LC_5_29_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \nx.i9205_1_lut_LC_5_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22917),
            .in3(_gnd_net_),
            .lcout(\nx.n13601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_67_LC_5_29_6 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_67_LC_5_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_67_LC_5_29_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_67_LC_5_29_6  (
            .in0(N__24372),
            .in1(N__24345),
            .in2(N__24321),
            .in3(N__24286),
            .lcout(\nx.n24_adj_717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7635_2_lut_3_lut_4_lut_4_lut_LC_6_16_3.C_ON=1'b0;
    defparam i7635_2_lut_3_lut_4_lut_4_lut_LC_6_16_3.SEQ_MODE=4'b0000;
    defparam i7635_2_lut_3_lut_4_lut_4_lut_LC_6_16_3.LUT_INIT=16'b1111101100000000;
    LogicCell40 i7635_2_lut_3_lut_4_lut_4_lut_LC_6_16_3 (
            .in0(N__42628),
            .in1(N__45671),
            .in2(N__44439),
            .in3(N__47624),
            .lcout(n11972),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9118_3_lut_4_lut_LC_6_17_0 .C_ON=1'b0;
    defparam \nx.i9118_3_lut_4_lut_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.i9118_3_lut_4_lut_LC_6_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9118_3_lut_4_lut_LC_6_17_0  (
            .in0(N__23261),
            .in1(N__23478),
            .in2(N__22881),
            .in3(N__23182),
            .lcout(\nx.n13514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9133_4_lut_LC_6_17_4 .C_ON=1'b0;
    defparam \nx.i9133_4_lut_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \nx.i9133_4_lut_LC_6_17_4 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \nx.i9133_4_lut_LC_6_17_4  (
            .in0(N__24941),
            .in1(N__23205),
            .in2(N__26804),
            .in3(N__22856),
            .lcout(\nx.n13513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.equal_372_i8_2_lut_LC_6_17_5 .C_ON=1'b0;
    defparam \nx.equal_372_i8_2_lut_LC_6_17_5 .SEQ_MODE=4'b0000;
    defparam \nx.equal_372_i8_2_lut_LC_6_17_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \nx.equal_372_i8_2_lut_LC_6_17_5  (
            .in0(_gnd_net_),
            .in1(N__23260),
            .in2(_gnd_net_),
            .in3(N__24940),
            .lcout(\nx.n7598 ),
            .ltout(\nx.n7598_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9095_3_lut_LC_6_17_6 .C_ON=1'b0;
    defparam \nx.i9095_3_lut_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9095_3_lut_LC_6_17_6 .LUT_INIT=16'b1111000011110011;
    LogicCell40 \nx.i9095_3_lut_LC_6_17_6  (
            .in0(_gnd_net_),
            .in1(N__22857),
            .in2(N__22836),
            .in3(N__23181),
            .lcout(\nx.n13435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_4_lut_4_lut_LC_6_18_0 .C_ON=1'b0;
    defparam \nx.i4_4_lut_4_lut_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.i4_4_lut_4_lut_LC_6_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \nx.i4_4_lut_4_lut_LC_6_18_0  (
            .in0(N__23476),
            .in1(N__23142),
            .in2(N__26797),
            .in3(N__26854),
            .lcout(\nx.n10_adj_760 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i26_LC_6_18_1 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i26_LC_6_18_1 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i26_LC_6_18_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i26_LC_6_18_1  (
            .in0(N__23304),
            .in1(N__23331),
            .in2(_gnd_net_),
            .in3(N__25238),
            .lcout(neo_pixel_transmitter_t0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46862),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8969_3_lut_LC_6_18_3 .C_ON=1'b0;
    defparam \nx.i8969_3_lut_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.i8969_3_lut_LC_6_18_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \nx.i8969_3_lut_LC_6_18_3  (
            .in0(N__26174),
            .in1(N__25756),
            .in2(_gnd_net_),
            .in3(N__24984),
            .lcout(\nx.n13364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4191_3_lut_LC_6_18_4 .C_ON=1'b0;
    defparam \nx.i4191_3_lut_LC_6_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.i4191_3_lut_LC_6_18_4 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \nx.i4191_3_lut_LC_6_18_4  (
            .in0(N__23477),
            .in1(N__26777),
            .in2(_gnd_net_),
            .in3(N__26708),
            .lcout(\nx.n7983 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i27_1_lut_LC_6_18_6 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i27_1_lut_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i27_1_lut_LC_6_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i27_1_lut_LC_6_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23303),
            .lcout(\nx.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_3_lut_adj_142_LC_6_19_1 .C_ON=1'b0;
    defparam \nx.i5_3_lut_adj_142_LC_6_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.i5_3_lut_adj_142_LC_6_19_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \nx.i5_3_lut_adj_142_LC_6_19_1  (
            .in0(N__26798),
            .in1(N__23283),
            .in2(_gnd_net_),
            .in3(N__23127),
            .lcout(\nx.n7994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam update_color_126_LC_6_19_2.C_ON=1'b0;
    defparam update_color_126_LC_6_19_2.SEQ_MODE=4'b1001;
    defparam update_color_126_LC_6_19_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 update_color_126_LC_6_19_2 (
            .in0(N__25053),
            .in1(N__25788),
            .in2(N__23277),
            .in3(N__24996),
            .lcout(update_color),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46866),
            .ce(),
            .sr(N__25047));
    defparam \nx.i9076_3_lut_4_lut_LC_6_19_3 .C_ON=1'b0;
    defparam \nx.i9076_3_lut_4_lut_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9076_3_lut_4_lut_LC_6_19_3 .LUT_INIT=16'b1010111110111111;
    LogicCell40 \nx.i9076_3_lut_4_lut_LC_6_19_3  (
            .in0(N__23262),
            .in1(N__23204),
            .in2(N__24956),
            .in3(N__23169),
            .lcout(),
            .ltout(\nx.n13436_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i822_4_lut_LC_6_19_4 .C_ON=1'b0;
    defparam \nx.i822_4_lut_LC_6_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.i822_4_lut_LC_6_19_4 .LUT_INIT=16'b0111001011111010;
    LogicCell40 \nx.i822_4_lut_LC_6_19_4  (
            .in0(N__23474),
            .in1(N__23141),
            .in2(N__23130),
            .in3(N__26853),
            .lcout(\nx.n3901 ),
            .ltout(\nx.n3901_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9173_4_lut_4_lut_LC_6_19_5 .C_ON=1'b0;
    defparam \nx.i9173_4_lut_4_lut_LC_6_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9173_4_lut_4_lut_LC_6_19_5 .LUT_INIT=16'b0000101000011011;
    LogicCell40 \nx.i9173_4_lut_4_lut_LC_6_19_5  (
            .in0(N__26799),
            .in1(N__23475),
            .in2(N__23409),
            .in3(N__23406),
            .lcout(\nx.n7657 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_2_lut_LC_6_20_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_2_lut_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_2_lut_LC_6_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_2_lut_LC_6_20_0  (
            .in0(_gnd_net_),
            .in1(N__23940),
            .in2(_gnd_net_),
            .in3(N__23391),
            .lcout(\nx.n1077 ),
            .ltout(),
            .carryin(bfn_6_20_0_),
            .carryout(\nx.n10743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_3_lut_LC_6_20_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_3_lut_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_3_lut_LC_6_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_3_lut_LC_6_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23583),
            .in3(N__23379),
            .lcout(\nx.n1076 ),
            .ltout(),
            .carryin(\nx.n10743 ),
            .carryout(\nx.n10744 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_4_lut_LC_6_20_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_4_lut_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_4_lut_LC_6_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_4_lut_LC_6_20_2  (
            .in0(_gnd_net_),
            .in1(N__42217),
            .in2(N__25415),
            .in3(N__23376),
            .lcout(\nx.n1075 ),
            .ltout(),
            .carryin(\nx.n10744 ),
            .carryout(\nx.n10745 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_5_lut_LC_6_20_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_5_lut_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_5_lut_LC_6_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_5_lut_LC_6_20_3  (
            .in0(_gnd_net_),
            .in1(N__42093),
            .in2(N__23651),
            .in3(N__23367),
            .lcout(\nx.n1074 ),
            .ltout(),
            .carryin(\nx.n10745 ),
            .carryout(\nx.n10746 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_6_lut_LC_6_20_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_6_lut_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_6_lut_LC_6_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_6_lut_LC_6_20_4  (
            .in0(_gnd_net_),
            .in1(N__42218),
            .in2(N__25395),
            .in3(N__23364),
            .lcout(\nx.n1073 ),
            .ltout(),
            .carryin(\nx.n10746 ),
            .carryout(\nx.n10747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_7_lut_LC_6_20_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_736_7_lut_LC_6_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_7_lut_LC_6_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_736_7_lut_LC_6_20_5  (
            .in0(_gnd_net_),
            .in1(N__42094),
            .in2(N__23603),
            .in3(N__23355),
            .lcout(\nx.n1072 ),
            .ltout(),
            .carryin(\nx.n10747 ),
            .carryout(\nx.n10748 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_736_8_lut_LC_6_20_6 .C_ON=1'b0;
    defparam \nx.mod_5_add_736_8_lut_LC_6_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_736_8_lut_LC_6_20_6 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_736_8_lut_LC_6_20_6  (
            .in0(N__42095),
            .in1(N__25614),
            .in2(N__23559),
            .in3(N__23352),
            .lcout(\nx.n1103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i676_3_lut_LC_6_20_7 .C_ON=1'b0;
    defparam \nx.mod_5_i676_3_lut_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i676_3_lut_LC_6_20_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i676_3_lut_LC_6_20_7  (
            .in0(_gnd_net_),
            .in1(N__25328),
            .in2(N__25284),
            .in3(N__25357),
            .lcout(\nx.n1009 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.sub_14_inv_0_i29_1_lut_LC_6_21_0 .C_ON=1'b0;
    defparam \nx.sub_14_inv_0_i29_1_lut_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.sub_14_inv_0_i29_1_lut_LC_6_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.sub_14_inv_0_i29_1_lut_LC_6_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25068),
            .lcout(\nx.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9195_2_lut_LC_6_21_2 .C_ON=1'b0;
    defparam \nx.i9195_2_lut_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9195_2_lut_LC_6_21_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \nx.i9195_2_lut_LC_6_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25695),
            .in3(N__25365),
            .lcout(\nx.n1007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i742_3_lut_LC_6_21_3 .C_ON=1'b0;
    defparam \nx.mod_5_i742_3_lut_LC_6_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i742_3_lut_LC_6_21_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i742_3_lut_LC_6_21_3  (
            .in0(_gnd_net_),
            .in1(N__23634),
            .in2(N__25416),
            .in3(N__23554),
            .lcout(\nx.n1107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i672_3_lut_LC_6_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i672_3_lut_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i672_3_lut_LC_6_21_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i672_3_lut_LC_6_21_4  (
            .in0(_gnd_net_),
            .in1(N__25641),
            .in2(N__25665),
            .in3(N__25366),
            .lcout(\nx.n1005 ),
            .ltout(\nx.n1005_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2_3_lut_LC_6_21_5 .C_ON=1'b0;
    defparam \nx.i2_3_lut_LC_6_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.i2_3_lut_LC_6_21_5 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i2_3_lut_LC_6_21_5  (
            .in0(_gnd_net_),
            .in1(N__23950),
            .in2(N__23586),
            .in3(N__23581),
            .lcout(),
            .ltout(\nx.n7_adj_690_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_4_lut_LC_6_21_6 .C_ON=1'b0;
    defparam \nx.i4_4_lut_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.i4_4_lut_LC_6_21_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \nx.i4_4_lut_LC_6_21_6  (
            .in0(N__25610),
            .in1(N__25422),
            .in2(N__23562),
            .in3(N__25411),
            .lcout(\nx.n1037 ),
            .ltout(\nx.n1037_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i740_3_lut_LC_6_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_i740_3_lut_LC_6_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i740_3_lut_LC_6_21_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i740_3_lut_LC_6_21_7  (
            .in0(N__25394),
            .in1(_gnd_net_),
            .in2(N__23526),
            .in3(N__23523),
            .lcout(\nx.n1105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8903_4_lut_LC_6_22_0 .C_ON=1'b0;
    defparam \nx.i8903_4_lut_LC_6_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.i8903_4_lut_LC_6_22_0 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \nx.i8903_4_lut_LC_6_22_0  (
            .in0(N__25938),
            .in1(N__25898),
            .in2(N__23751),
            .in3(N__25559),
            .lcout(\nx.n7899 ),
            .ltout(\nx.n7899_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_3_lut_4_lut_adj_144_LC_6_22_1 .C_ON=1'b0;
    defparam \nx.i1_3_lut_4_lut_adj_144_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_3_lut_4_lut_adj_144_LC_6_22_1 .LUT_INIT=16'b0000011100001011;
    LogicCell40 \nx.i1_3_lut_4_lut_adj_144_LC_6_22_1  (
            .in0(N__25560),
            .in1(N__25326),
            .in2(N__23754),
            .in3(N__25940),
            .lcout(\nx.n12839 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_3_lut_LC_6_22_2 .C_ON=1'b0;
    defparam \nx.i1_3_lut_LC_6_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_3_lut_LC_6_22_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i1_3_lut_LC_6_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25856),
            .in3(N__25830),
            .lcout(\nx.n740 ),
            .ltout(\nx.n740_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8902_4_lut_LC_6_22_3 .C_ON=1'b0;
    defparam \nx.i8902_4_lut_LC_6_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.i8902_4_lut_LC_6_22_3 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \nx.i8902_4_lut_LC_6_22_3  (
            .in0(N__25897),
            .in1(N__25947),
            .in2(N__23742),
            .in3(N__26081),
            .lcout(\nx.n11866 ),
            .ltout(\nx.n11866_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_LC_6_22_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_LC_6_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_LC_6_22_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \nx.i1_4_lut_LC_6_22_4  (
            .in0(N__26088),
            .in1(_gnd_net_),
            .in2(N__23739),
            .in3(N__25594),
            .lcout(\nx.n838 ),
            .ltout(\nx.n838_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_43_LC_6_22_5 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_43_LC_6_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_43_LC_6_22_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \nx.i1_2_lut_adj_43_LC_6_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23736),
            .in3(N__25939),
            .lcout(\nx.n7497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_3_lut_LC_6_22_6 .C_ON=1'b0;
    defparam \nx.i12_3_lut_LC_6_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.i12_3_lut_LC_6_22_6 .LUT_INIT=16'b0011000000001100;
    LogicCell40 \nx.i12_3_lut_LC_6_22_6  (
            .in0(_gnd_net_),
            .in1(N__26025),
            .in2(N__25984),
            .in3(N__26069),
            .lcout(\nx.n708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5701_4_lut_LC_6_22_7.C_ON=1'b0;
    defparam i5701_4_lut_LC_6_22_7.SEQ_MODE=4'b0000;
    defparam i5701_4_lut_LC_6_22_7.LUT_INIT=16'b0011001100110010;
    LogicCell40 i5701_4_lut_LC_6_22_7 (
            .in0(N__23733),
            .in1(N__23718),
            .in2(N__23697),
            .in3(N__23682),
            .lcout(n1907),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.bit_ctr__i0_LC_6_23_0 .C_ON=1'b1;
    defparam \nx.bit_ctr__i0_LC_6_23_0 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i0_LC_6_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i0_LC_6_23_0  (
            .in0(_gnd_net_),
            .in1(N__26155),
            .in2(_gnd_net_),
            .in3(N__23670),
            .lcout(\nx.bit_ctr_0 ),
            .ltout(),
            .carryin(bfn_6_23_0_),
            .carryout(\nx.n10613 ),
            .clk(N__46875),
            .ce(N__24240),
            .sr(N__24208));
    defparam \nx.bit_ctr__i1_LC_6_23_1 .C_ON=1'b1;
    defparam \nx.bit_ctr__i1_LC_6_23_1 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i1_LC_6_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i1_LC_6_23_1  (
            .in0(_gnd_net_),
            .in1(N__24842),
            .in2(_gnd_net_),
            .in3(N__23667),
            .lcout(\nx.bit_ctr_1 ),
            .ltout(),
            .carryin(\nx.n10613 ),
            .carryout(\nx.n10614 ),
            .clk(N__46875),
            .ce(N__24240),
            .sr(N__24208));
    defparam \nx.bit_ctr__i2_LC_6_23_2 .C_ON=1'b1;
    defparam \nx.bit_ctr__i2_LC_6_23_2 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i2_LC_6_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i2_LC_6_23_2  (
            .in0(_gnd_net_),
            .in1(N__26870),
            .in2(_gnd_net_),
            .in3(N__23784),
            .lcout(\nx.bit_ctr_2 ),
            .ltout(),
            .carryin(\nx.n10614 ),
            .carryout(\nx.n10615 ),
            .clk(N__46875),
            .ce(N__24240),
            .sr(N__24208));
    defparam \nx.bit_ctr__i3_LC_6_23_3 .C_ON=1'b1;
    defparam \nx.bit_ctr__i3_LC_6_23_3 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i3_LC_6_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i3_LC_6_23_3  (
            .in0(_gnd_net_),
            .in1(N__30792),
            .in2(_gnd_net_),
            .in3(N__23781),
            .lcout(\nx.bit_ctr_3 ),
            .ltout(),
            .carryin(\nx.n10615 ),
            .carryout(\nx.n10616 ),
            .clk(N__46875),
            .ce(N__24240),
            .sr(N__24208));
    defparam \nx.bit_ctr__i4_LC_6_23_4 .C_ON=1'b1;
    defparam \nx.bit_ctr__i4_LC_6_23_4 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i4_LC_6_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i4_LC_6_23_4  (
            .in0(_gnd_net_),
            .in1(N__32392),
            .in2(_gnd_net_),
            .in3(N__23778),
            .lcout(\nx.bit_ctr_4 ),
            .ltout(),
            .carryin(\nx.n10616 ),
            .carryout(\nx.n10617 ),
            .clk(N__46875),
            .ce(N__24240),
            .sr(N__24208));
    defparam \nx.bit_ctr__i5_LC_6_23_5 .C_ON=1'b1;
    defparam \nx.bit_ctr__i5_LC_6_23_5 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i5_LC_6_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i5_LC_6_23_5  (
            .in0(_gnd_net_),
            .in1(N__29329),
            .in2(_gnd_net_),
            .in3(N__23775),
            .lcout(\nx.bit_ctr_5 ),
            .ltout(),
            .carryin(\nx.n10617 ),
            .carryout(\nx.n10618 ),
            .clk(N__46875),
            .ce(N__24240),
            .sr(N__24208));
    defparam \nx.bit_ctr__i6_LC_6_23_6 .C_ON=1'b1;
    defparam \nx.bit_ctr__i6_LC_6_23_6 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i6_LC_6_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i6_LC_6_23_6  (
            .in0(_gnd_net_),
            .in1(N__35233),
            .in2(_gnd_net_),
            .in3(N__23772),
            .lcout(\nx.bit_ctr_6 ),
            .ltout(),
            .carryin(\nx.n10618 ),
            .carryout(\nx.n10619 ),
            .clk(N__46875),
            .ce(N__24240),
            .sr(N__24208));
    defparam \nx.bit_ctr__i7_LC_6_23_7 .C_ON=1'b1;
    defparam \nx.bit_ctr__i7_LC_6_23_7 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i7_LC_6_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i7_LC_6_23_7  (
            .in0(_gnd_net_),
            .in1(N__28205),
            .in2(_gnd_net_),
            .in3(N__23769),
            .lcout(\nx.bit_ctr_7 ),
            .ltout(),
            .carryin(\nx.n10619 ),
            .carryout(\nx.n10620 ),
            .clk(N__46875),
            .ce(N__24240),
            .sr(N__24208));
    defparam \nx.bit_ctr__i8_LC_6_24_0 .C_ON=1'b1;
    defparam \nx.bit_ctr__i8_LC_6_24_0 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i8_LC_6_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i8_LC_6_24_0  (
            .in0(_gnd_net_),
            .in1(N__30123),
            .in2(_gnd_net_),
            .in3(N__23766),
            .lcout(\nx.bit_ctr_8 ),
            .ltout(),
            .carryin(bfn_6_24_0_),
            .carryout(\nx.n10621 ),
            .clk(N__46876),
            .ce(N__24250),
            .sr(N__24212));
    defparam \nx.bit_ctr__i9_LC_6_24_1 .C_ON=1'b1;
    defparam \nx.bit_ctr__i9_LC_6_24_1 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i9_LC_6_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i9_LC_6_24_1  (
            .in0(_gnd_net_),
            .in1(N__38913),
            .in2(_gnd_net_),
            .in3(N__23763),
            .lcout(\nx.bit_ctr_9 ),
            .ltout(),
            .carryin(\nx.n10621 ),
            .carryout(\nx.n10622 ),
            .clk(N__46876),
            .ce(N__24250),
            .sr(N__24212));
    defparam \nx.bit_ctr__i10_LC_6_24_2 .C_ON=1'b1;
    defparam \nx.bit_ctr__i10_LC_6_24_2 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i10_LC_6_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i10_LC_6_24_2  (
            .in0(_gnd_net_),
            .in1(N__39899),
            .in2(_gnd_net_),
            .in3(N__23760),
            .lcout(\nx.bit_ctr_10 ),
            .ltout(),
            .carryin(\nx.n10622 ),
            .carryout(\nx.n10623 ),
            .clk(N__46876),
            .ce(N__24250),
            .sr(N__24212));
    defparam \nx.bit_ctr__i11_LC_6_24_3 .C_ON=1'b1;
    defparam \nx.bit_ctr__i11_LC_6_24_3 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i11_LC_6_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i11_LC_6_24_3  (
            .in0(_gnd_net_),
            .in1(N__36045),
            .in2(_gnd_net_),
            .in3(N__23757),
            .lcout(\nx.bit_ctr_11 ),
            .ltout(),
            .carryin(\nx.n10623 ),
            .carryout(\nx.n10624 ),
            .clk(N__46876),
            .ce(N__24250),
            .sr(N__24212));
    defparam \nx.bit_ctr__i12_LC_6_24_4 .C_ON=1'b1;
    defparam \nx.bit_ctr__i12_LC_6_24_4 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i12_LC_6_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i12_LC_6_24_4  (
            .in0(_gnd_net_),
            .in1(N__34328),
            .in2(_gnd_net_),
            .in3(N__23889),
            .lcout(\nx.bit_ctr_12 ),
            .ltout(),
            .carryin(\nx.n10624 ),
            .carryout(\nx.n10625 ),
            .clk(N__46876),
            .ce(N__24250),
            .sr(N__24212));
    defparam \nx.bit_ctr__i13_LC_6_24_5 .C_ON=1'b1;
    defparam \nx.bit_ctr__i13_LC_6_24_5 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i13_LC_6_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i13_LC_6_24_5  (
            .in0(_gnd_net_),
            .in1(N__31779),
            .in2(_gnd_net_),
            .in3(N__23886),
            .lcout(\nx.bit_ctr_13 ),
            .ltout(),
            .carryin(\nx.n10625 ),
            .carryout(\nx.n10626 ),
            .clk(N__46876),
            .ce(N__24250),
            .sr(N__24212));
    defparam \nx.bit_ctr__i14_LC_6_24_6 .C_ON=1'b1;
    defparam \nx.bit_ctr__i14_LC_6_24_6 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i14_LC_6_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i14_LC_6_24_6  (
            .in0(_gnd_net_),
            .in1(N__30510),
            .in2(_gnd_net_),
            .in3(N__23883),
            .lcout(\nx.bit_ctr_14 ),
            .ltout(),
            .carryin(\nx.n10626 ),
            .carryout(\nx.n10627 ),
            .clk(N__46876),
            .ce(N__24250),
            .sr(N__24212));
    defparam \nx.bit_ctr__i15_LC_6_24_7 .C_ON=1'b1;
    defparam \nx.bit_ctr__i15_LC_6_24_7 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i15_LC_6_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i15_LC_6_24_7  (
            .in0(_gnd_net_),
            .in1(N__28917),
            .in2(_gnd_net_),
            .in3(N__23880),
            .lcout(\nx.bit_ctr_15 ),
            .ltout(),
            .carryin(\nx.n10627 ),
            .carryout(\nx.n10628 ),
            .clk(N__46876),
            .ce(N__24250),
            .sr(N__24212));
    defparam \nx.bit_ctr__i16_LC_6_25_0 .C_ON=1'b1;
    defparam \nx.bit_ctr__i16_LC_6_25_0 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i16_LC_6_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i16_LC_6_25_0  (
            .in0(_gnd_net_),
            .in1(N__26354),
            .in2(_gnd_net_),
            .in3(N__23877),
            .lcout(\nx.bit_ctr_16 ),
            .ltout(),
            .carryin(bfn_6_25_0_),
            .carryout(\nx.n10629 ),
            .clk(N__46878),
            .ce(N__24255),
            .sr(N__24213));
    defparam \nx.bit_ctr__i17_LC_6_25_1 .C_ON=1'b1;
    defparam \nx.bit_ctr__i17_LC_6_25_1 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i17_LC_6_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i17_LC_6_25_1  (
            .in0(_gnd_net_),
            .in1(N__25514),
            .in2(_gnd_net_),
            .in3(N__23874),
            .lcout(\nx.bit_ctr_17 ),
            .ltout(),
            .carryin(\nx.n10629 ),
            .carryout(\nx.n10630 ),
            .clk(N__46878),
            .ce(N__24255),
            .sr(N__24213));
    defparam \nx.bit_ctr__i18_LC_6_25_2 .C_ON=1'b1;
    defparam \nx.bit_ctr__i18_LC_6_25_2 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i18_LC_6_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i18_LC_6_25_2  (
            .in0(_gnd_net_),
            .in1(N__24753),
            .in2(_gnd_net_),
            .in3(N__23871),
            .lcout(\nx.bit_ctr_18 ),
            .ltout(),
            .carryin(\nx.n10630 ),
            .carryout(\nx.n10631 ),
            .clk(N__46878),
            .ce(N__24255),
            .sr(N__24213));
    defparam \nx.bit_ctr__i19_LC_6_25_3 .C_ON=1'b1;
    defparam \nx.bit_ctr__i19_LC_6_25_3 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i19_LC_6_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i19_LC_6_25_3  (
            .in0(_gnd_net_),
            .in1(N__23865),
            .in2(_gnd_net_),
            .in3(N__23832),
            .lcout(\nx.bit_ctr_19 ),
            .ltout(),
            .carryin(\nx.n10631 ),
            .carryout(\nx.n10632 ),
            .clk(N__46878),
            .ce(N__24255),
            .sr(N__24213));
    defparam \nx.bit_ctr__i20_LC_6_25_4 .C_ON=1'b1;
    defparam \nx.bit_ctr__i20_LC_6_25_4 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i20_LC_6_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i20_LC_6_25_4  (
            .in0(_gnd_net_),
            .in1(N__23813),
            .in2(_gnd_net_),
            .in3(N__24108),
            .lcout(\nx.bit_ctr_20 ),
            .ltout(),
            .carryin(\nx.n10632 ),
            .carryout(\nx.n10633 ),
            .clk(N__46878),
            .ce(N__24255),
            .sr(N__24213));
    defparam \nx.bit_ctr__i21_LC_6_25_5 .C_ON=1'b1;
    defparam \nx.bit_ctr__i21_LC_6_25_5 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i21_LC_6_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i21_LC_6_25_5  (
            .in0(_gnd_net_),
            .in1(N__24092),
            .in2(_gnd_net_),
            .in3(N__24060),
            .lcout(\nx.bit_ctr_21 ),
            .ltout(),
            .carryin(\nx.n10633 ),
            .carryout(\nx.n10634 ),
            .clk(N__46878),
            .ce(N__24255),
            .sr(N__24213));
    defparam \nx.bit_ctr__i22_LC_6_25_6 .C_ON=1'b1;
    defparam \nx.bit_ctr__i22_LC_6_25_6 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i22_LC_6_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i22_LC_6_25_6  (
            .in0(_gnd_net_),
            .in1(N__25463),
            .in2(_gnd_net_),
            .in3(N__24057),
            .lcout(\nx.bit_ctr_22 ),
            .ltout(),
            .carryin(\nx.n10634 ),
            .carryout(\nx.n10635 ),
            .clk(N__46878),
            .ce(N__24255),
            .sr(N__24213));
    defparam \nx.bit_ctr__i23_LC_6_25_7 .C_ON=1'b1;
    defparam \nx.bit_ctr__i23_LC_6_25_7 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i23_LC_6_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i23_LC_6_25_7  (
            .in0(_gnd_net_),
            .in1(N__24044),
            .in2(_gnd_net_),
            .in3(N__24003),
            .lcout(\nx.bit_ctr_23 ),
            .ltout(),
            .carryin(\nx.n10635 ),
            .carryout(\nx.n10636 ),
            .clk(N__46878),
            .ce(N__24255),
            .sr(N__24213));
    defparam \nx.bit_ctr__i24_LC_6_26_0 .C_ON=1'b1;
    defparam \nx.bit_ctr__i24_LC_6_26_0 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i24_LC_6_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i24_LC_6_26_0  (
            .in0(_gnd_net_),
            .in1(N__23987),
            .in2(_gnd_net_),
            .in3(N__23955),
            .lcout(\nx.bit_ctr_24 ),
            .ltout(),
            .carryin(bfn_6_26_0_),
            .carryout(\nx.n10637 ),
            .clk(N__46882),
            .ce(N__24254),
            .sr(N__24204));
    defparam \nx.bit_ctr__i25_LC_6_26_1 .C_ON=1'b1;
    defparam \nx.bit_ctr__i25_LC_6_26_1 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i25_LC_6_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i25_LC_6_26_1  (
            .in0(_gnd_net_),
            .in1(N__23939),
            .in2(_gnd_net_),
            .in3(N__23901),
            .lcout(\nx.bit_ctr_25 ),
            .ltout(),
            .carryin(\nx.n10637 ),
            .carryout(\nx.n10638 ),
            .clk(N__46882),
            .ce(N__24254),
            .sr(N__24204));
    defparam \nx.bit_ctr__i26_LC_6_26_2 .C_ON=1'b1;
    defparam \nx.bit_ctr__i26_LC_6_26_2 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i26_LC_6_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i26_LC_6_26_2  (
            .in0(_gnd_net_),
            .in1(N__25313),
            .in2(_gnd_net_),
            .in3(N__23898),
            .lcout(\nx.bit_ctr_26 ),
            .ltout(),
            .carryin(\nx.n10638 ),
            .carryout(\nx.n10639 ),
            .clk(N__46882),
            .ce(N__24254),
            .sr(N__24204));
    defparam \nx.bit_ctr__i27_LC_6_26_3 .C_ON=1'b1;
    defparam \nx.bit_ctr__i27_LC_6_26_3 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i27_LC_6_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i27_LC_6_26_3  (
            .in0(_gnd_net_),
            .in1(N__25925),
            .in2(_gnd_net_),
            .in3(N__23895),
            .lcout(\nx.bit_ctr_27 ),
            .ltout(),
            .carryin(\nx.n10639 ),
            .carryout(\nx.n10640 ),
            .clk(N__46882),
            .ce(N__24254),
            .sr(N__24204));
    defparam \nx.bit_ctr__i28_LC_6_26_4 .C_ON=1'b1;
    defparam \nx.bit_ctr__i28_LC_6_26_4 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i28_LC_6_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i28_LC_6_26_4  (
            .in0(_gnd_net_),
            .in1(N__25893),
            .in2(_gnd_net_),
            .in3(N__23892),
            .lcout(\nx.bit_ctr_28 ),
            .ltout(),
            .carryin(\nx.n10640 ),
            .carryout(\nx.n10641 ),
            .clk(N__46882),
            .ce(N__24254),
            .sr(N__24204));
    defparam \nx.bit_ctr__i29_LC_6_26_5 .C_ON=1'b1;
    defparam \nx.bit_ctr__i29_LC_6_26_5 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i29_LC_6_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i29_LC_6_26_5  (
            .in0(_gnd_net_),
            .in1(N__26068),
            .in2(_gnd_net_),
            .in3(N__24264),
            .lcout(\nx.bit_ctr_29 ),
            .ltout(),
            .carryin(\nx.n10641 ),
            .carryout(\nx.n10642 ),
            .clk(N__46882),
            .ce(N__24254),
            .sr(N__24204));
    defparam \nx.bit_ctr__i30_LC_6_26_6 .C_ON=1'b1;
    defparam \nx.bit_ctr__i30_LC_6_26_6 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i30_LC_6_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i30_LC_6_26_6  (
            .in0(_gnd_net_),
            .in1(N__26016),
            .in2(_gnd_net_),
            .in3(N__24261),
            .lcout(\nx.bit_ctr_30 ),
            .ltout(),
            .carryin(\nx.n10642 ),
            .carryout(\nx.n10643 ),
            .clk(N__46882),
            .ce(N__24254),
            .sr(N__24204));
    defparam \nx.bit_ctr__i31_LC_6_26_7 .C_ON=1'b0;
    defparam \nx.bit_ctr__i31_LC_6_26_7 .SEQ_MODE=4'b1000;
    defparam \nx.bit_ctr__i31_LC_6_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.bit_ctr__i31_LC_6_26_7  (
            .in0(_gnd_net_),
            .in1(N__25974),
            .in2(_gnd_net_),
            .in3(N__24258),
            .lcout(\nx.bit_ctr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46882),
            .ce(N__24254),
            .sr(N__24204));
    defparam \nx.mod_5_add_1272_2_lut_LC_6_27_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_2_lut_LC_6_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_2_lut_LC_6_27_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1272_2_lut_LC_6_27_0  (
            .in0(N__25524),
            .in1(N__25523),
            .in2(N__24416),
            .in3(N__24168),
            .lcout(\nx.n1909 ),
            .ltout(),
            .carryin(bfn_6_27_0_),
            .carryout(\nx.n10819 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_3_lut_LC_6_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_3_lut_LC_6_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_3_lut_LC_6_27_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_1272_3_lut_LC_6_27_1  (
            .in0(N__24602),
            .in1(N__24601),
            .in2(N__24417),
            .in3(N__24165),
            .lcout(\nx.n1908 ),
            .ltout(),
            .carryin(\nx.n10819 ),
            .carryout(\nx.n10820 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_4_lut_LC_6_27_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_4_lut_LC_6_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_4_lut_LC_6_27_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_4_lut_LC_6_27_2  (
            .in0(N__24626),
            .in1(N__24625),
            .in2(N__24511),
            .in3(N__24162),
            .lcout(\nx.n1907 ),
            .ltout(),
            .carryin(\nx.n10820 ),
            .carryout(\nx.n10821 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_5_lut_LC_6_27_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_5_lut_LC_6_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_5_lut_LC_6_27_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_5_lut_LC_6_27_3  (
            .in0(N__24159),
            .in1(N__24158),
            .in2(N__24514),
            .in3(N__24141),
            .lcout(\nx.n1906 ),
            .ltout(),
            .carryin(\nx.n10821 ),
            .carryout(\nx.n10822 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_6_lut_LC_6_27_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_6_lut_LC_6_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_6_lut_LC_6_27_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_6_lut_LC_6_27_4  (
            .in0(N__24134),
            .in1(N__24133),
            .in2(N__24512),
            .in3(N__24114),
            .lcout(\nx.n1905 ),
            .ltout(),
            .carryin(\nx.n10822 ),
            .carryout(\nx.n10823 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_7_lut_LC_6_27_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_7_lut_LC_6_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_7_lut_LC_6_27_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_7_lut_LC_6_27_5  (
            .in0(N__24674),
            .in1(N__24673),
            .in2(N__24515),
            .in3(N__24111),
            .lcout(\nx.n1904 ),
            .ltout(),
            .carryin(\nx.n10823 ),
            .carryout(\nx.n10824 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_8_lut_LC_6_27_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_8_lut_LC_6_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_8_lut_LC_6_27_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_8_lut_LC_6_27_6  (
            .in0(N__24371),
            .in1(N__24370),
            .in2(N__24513),
            .in3(N__24351),
            .lcout(\nx.n1903 ),
            .ltout(),
            .carryin(\nx.n10824 ),
            .carryout(\nx.n10825 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_9_lut_LC_6_27_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_9_lut_LC_6_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_9_lut_LC_6_27_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_9_lut_LC_6_27_7  (
            .in0(N__24581),
            .in1(N__24580),
            .in2(N__24516),
            .in3(N__24348),
            .lcout(\nx.n1902 ),
            .ltout(),
            .carryin(\nx.n10825 ),
            .carryout(\nx.n10826 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_10_lut_LC_6_28_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_10_lut_LC_6_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_10_lut_LC_6_28_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_10_lut_LC_6_28_0  (
            .in0(N__24344),
            .in1(N__24343),
            .in2(N__24504),
            .in3(N__24324),
            .lcout(\nx.n1901 ),
            .ltout(),
            .carryin(bfn_6_28_0_),
            .carryout(\nx.n10827 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_11_lut_LC_6_28_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_11_lut_LC_6_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_11_lut_LC_6_28_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_11_lut_LC_6_28_1  (
            .in0(N__24320),
            .in1(N__24319),
            .in2(N__24508),
            .in3(N__24300),
            .lcout(\nx.n1900 ),
            .ltout(),
            .carryin(\nx.n10827 ),
            .carryout(\nx.n10828 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_12_lut_LC_6_28_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_12_lut_LC_6_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_12_lut_LC_6_28_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_12_lut_LC_6_28_2  (
            .in0(N__24561),
            .in1(N__24560),
            .in2(N__24505),
            .in3(N__24297),
            .lcout(\nx.n1899 ),
            .ltout(),
            .carryin(\nx.n10828 ),
            .carryout(\nx.n10829 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_13_lut_LC_6_28_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_13_lut_LC_6_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_13_lut_LC_6_28_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_13_lut_LC_6_28_3  (
            .in0(N__24696),
            .in1(N__24695),
            .in2(N__24509),
            .in3(N__24294),
            .lcout(\nx.n1898 ),
            .ltout(),
            .carryin(\nx.n10829 ),
            .carryout(\nx.n10830 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_14_lut_LC_6_28_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_14_lut_LC_6_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_14_lut_LC_6_28_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_14_lut_LC_6_28_4  (
            .in0(N__24648),
            .in1(N__24647),
            .in2(N__24506),
            .in3(N__24291),
            .lcout(\nx.n1897 ),
            .ltout(),
            .carryin(\nx.n10830 ),
            .carryout(\nx.n10831 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_15_lut_LC_6_28_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1272_15_lut_LC_6_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_15_lut_LC_6_28_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_15_lut_LC_6_28_5  (
            .in0(N__24288),
            .in1(N__24287),
            .in2(N__24510),
            .in3(N__24270),
            .lcout(\nx.n1896 ),
            .ltout(),
            .carryin(\nx.n10831 ),
            .carryout(\nx.n10832 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1272_16_lut_LC_6_28_6 .C_ON=1'b0;
    defparam \nx.mod_5_add_1272_16_lut_LC_6_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1272_16_lut_LC_6_28_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_1272_16_lut_LC_6_28_6  (
            .in0(N__24539),
            .in1(N__24540),
            .in2(N__24507),
            .in3(N__24267),
            .lcout(\nx.n1895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_adj_133_LC_6_29_0 .C_ON=1'b0;
    defparam \nx.i20_4_lut_adj_133_LC_6_29_0 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_adj_133_LC_6_29_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i20_4_lut_adj_133_LC_6_29_0  (
            .in0(N__25941),
            .in1(N__25978),
            .in2(N__24765),
            .in3(N__39921),
            .lcout(\nx.n48_adj_778 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_69_LC_6_29_2 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_69_LC_6_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_69_LC_6_29_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_69_LC_6_29_2  (
            .in0(N__24702),
            .in1(N__24694),
            .in2(N__24678),
            .in3(N__24654),
            .lcout(),
            .ltout(\nx.n26_adj_719_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_70_LC_6_29_3 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_70_LC_6_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_70_LC_6_29_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_70_LC_6_29_3  (
            .in0(N__24640),
            .in1(N__24627),
            .in2(N__24606),
            .in3(N__24522),
            .lcout(\nx.n1829 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5924_2_lut_LC_6_29_4 .C_ON=1'b0;
    defparam \nx.i5924_2_lut_LC_6_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.i5924_2_lut_LC_6_29_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \nx.i5924_2_lut_LC_6_29_4  (
            .in0(N__25515),
            .in1(N__24603),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\nx.n9717_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8_4_lut_adj_68_LC_6_29_5 .C_ON=1'b0;
    defparam \nx.i8_4_lut_adj_68_LC_6_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.i8_4_lut_adj_68_LC_6_29_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i8_4_lut_adj_68_LC_6_29_5  (
            .in0(N__24582),
            .in1(N__24559),
            .in2(N__24543),
            .in3(N__24538),
            .lcout(\nx.n22_adj_718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9209_1_lut_LC_6_29_6 .C_ON=1'b0;
    defparam \nx.i9209_1_lut_LC_6_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9209_1_lut_LC_6_29_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.i9209_1_lut_LC_6_29_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24450),
            .lcout(\nx.n13605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7629_2_lut_3_lut_4_lut_4_lut_LC_7_16_0.C_ON=1'b0;
    defparam i7629_2_lut_3_lut_4_lut_4_lut_LC_7_16_0.SEQ_MODE=4'b0000;
    defparam i7629_2_lut_3_lut_4_lut_4_lut_LC_7_16_0.LUT_INIT=16'b1100110011001000;
    LogicCell40 i7629_2_lut_3_lut_4_lut_4_lut_LC_7_16_0 (
            .in0(N__44435),
            .in1(N__47519),
            .in2(N__45682),
            .in3(N__42627),
            .lcout(n11966),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i7_LC_7_16_1.C_ON=1'b0;
    defparam pin_output_enable__i7_LC_7_16_1.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i7_LC_7_16_1.LUT_INIT=16'b1011100010101010;
    LogicCell40 pin_output_enable__i7_LC_7_16_1 (
            .in0(N__24383),
            .in1(N__32424),
            .in2(N__47610),
            .in3(N__47153),
            .lcout(pin_oe_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46867),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.one_wire_108_LC_7_17_4 .C_ON=1'b0;
    defparam \nx.one_wire_108_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \nx.one_wire_108_LC_7_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.one_wire_108_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24955),
            .lcout(NEOPXL_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46857),
            .ce(N__24864),
            .sr(N__24855));
    defparam \nx.i8968_3_lut_LC_7_18_0 .C_ON=1'b0;
    defparam \nx.i8968_3_lut_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.i8968_3_lut_LC_7_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \nx.i8968_3_lut_LC_7_18_0  (
            .in0(N__26170),
            .in1(N__25025),
            .in2(_gnd_net_),
            .in3(N__26605),
            .lcout(\nx.n13363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_107_LC_7_18_1 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_107_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_107_LC_7_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \nx.i1_2_lut_adj_107_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(N__30811),
            .in2(_gnd_net_),
            .in3(N__26565),
            .lcout(\nx.n11156 ),
            .ltout(\nx.n11156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.bit_ctr_1__bdd_4_lut_LC_7_18_2 .C_ON=1'b0;
    defparam \nx.bit_ctr_1__bdd_4_lut_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.bit_ctr_1__bdd_4_lut_LC_7_18_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \nx.bit_ctr_1__bdd_4_lut_LC_7_18_2  (
            .in0(N__24846),
            .in1(N__24828),
            .in2(N__24822),
            .in3(N__24819),
            .lcout(),
            .ltout(\nx.n13619_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.n13619_bdd_4_lut_LC_7_18_3 .C_ON=1'b0;
    defparam \nx.n13619_bdd_4_lut_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.n13619_bdd_4_lut_LC_7_18_3 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \nx.n13619_bdd_4_lut_LC_7_18_3  (
            .in0(N__24771),
            .in1(N__26139),
            .in2(N__24813),
            .in3(N__24810),
            .lcout(\nx.n13622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i2_LC_7_18_4.C_ON=1'b0;
    defparam pin_output_enable__i2_LC_7_18_4.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i2_LC_7_18_4.LUT_INIT=16'b1101100011001100;
    LogicCell40 pin_output_enable__i2_LC_7_18_4 (
            .in0(N__24804),
            .in1(N__24782),
            .in2(N__47674),
            .in3(N__47157),
            .lcout(pin_oe_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46868),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8977_3_lut_LC_7_18_6 .C_ON=1'b0;
    defparam \nx.i8977_3_lut_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.i8977_3_lut_LC_7_18_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.i8977_3_lut_LC_7_18_6  (
            .in0(N__32221),
            .in1(_gnd_net_),
            .in2(N__26175),
            .in3(N__27289),
            .lcout(\nx.n13372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_84_LC_7_19_1 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_84_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_84_LC_7_19_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_84_LC_7_19_1  (
            .in0(N__33164),
            .in1(N__33131),
            .in2(N__32767),
            .in3(N__33092),
            .lcout(\nx.n44_adj_741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9204_1_lut_LC_7_19_3 .C_ON=1'b0;
    defparam \nx.i9204_1_lut_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9204_1_lut_LC_7_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \nx.i9204_1_lut_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29669),
            .lcout(\nx.n13600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.neo_pixel_transmitter_t0_i0_i28_LC_7_19_5 .C_ON=1'b0;
    defparam \nx.neo_pixel_transmitter_t0_i0_i28_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \nx.neo_pixel_transmitter_t0_i0_i28_LC_7_19_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.neo_pixel_transmitter_t0_i0_i28_LC_7_19_5  (
            .in0(N__25269),
            .in1(N__25067),
            .in2(_gnd_net_),
            .in3(N__25219),
            .lcout(neo_pixel_transmitter_t0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46872),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_7_20_0.C_ON=1'b0;
    defparam i1_4_lut_LC_7_20_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_7_20_0.LUT_INIT=16'b0110111111110110;
    LogicCell40 i1_4_lut_LC_7_20_0 (
            .in0(N__32222),
            .in1(N__24990),
            .in2(N__24983),
            .in3(N__25032),
            .lcout(n9_adj_847),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i13_LC_7_20_1.C_ON=1'b0;
    defparam neopxl_color_prev_i13_LC_7_20_1.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i13_LC_7_20_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 neopxl_color_prev_i13_LC_7_20_1 (
            .in0(N__25024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(neopxl_color_prev_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46873),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i13_LC_7_20_2.C_ON=1'b0;
    defparam neopxl_color_i13_LC_7_20_2.SEQ_MODE=4'b1000;
    defparam neopxl_color_i13_LC_7_20_2.LUT_INIT=16'b1111011100010000;
    LogicCell40 neopxl_color_i13_LC_7_20_2 (
            .in0(N__47516),
            .in1(N__43894),
            .in2(N__43692),
            .in3(N__25023),
            .lcout(neopxl_color_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46873),
            .ce(),
            .sr(_gnd_net_));
    defparam i9171_2_lut_3_lut_LC_7_20_3.C_ON=1'b0;
    defparam i9171_2_lut_3_lut_LC_7_20_3.SEQ_MODE=4'b0000;
    defparam i9171_2_lut_3_lut_LC_7_20_3.LUT_INIT=16'b0000000000010001;
    LogicCell40 i9171_2_lut_3_lut_LC_7_20_3 (
            .in0(N__43893),
            .in1(N__47515),
            .in2(_gnd_net_),
            .in3(N__43676),
            .lcout(current_pin_7__N_153),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i14_LC_7_20_4.C_ON=1'b0;
    defparam neopxl_color_prev_i14_LC_7_20_4.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i14_LC_7_20_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 neopxl_color_prev_i14_LC_7_20_4 (
            .in0(N__24979),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(neopxl_color_prev_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46873),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_7_20_5.C_ON=1'b0;
    defparam i3_4_lut_LC_7_20_5.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_7_20_5.LUT_INIT=16'b0110111111110110;
    LogicCell40 i3_4_lut_LC_7_20_5 (
            .in0(N__27027),
            .in1(N__27294),
            .in2(N__25026),
            .in3(N__25002),
            .lcout(n11_adj_845),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i4_LC_7_20_6.C_ON=1'b0;
    defparam neopxl_color_prev_i4_LC_7_20_6.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i4_LC_7_20_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 neopxl_color_prev_i4_LC_7_20_6 (
            .in0(N__32223),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(neopxl_color_prev_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46873),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i14_LC_7_20_7.C_ON=1'b0;
    defparam neopxl_color_i14_LC_7_20_7.SEQ_MODE=4'b1000;
    defparam neopxl_color_i14_LC_7_20_7.LUT_INIT=16'b1100110101001100;
    LogicCell40 neopxl_color_i14_LC_7_20_7 (
            .in0(N__43895),
            .in1(N__24978),
            .in2(N__47631),
            .in3(N__43680),
            .lcout(neopxl_color_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46873),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7605_3_lut_LC_7_21_0 .C_ON=1'b0;
    defparam \nx.i7605_3_lut_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.i7605_3_lut_LC_7_21_0 .LUT_INIT=16'b1111000011110011;
    LogicCell40 \nx.i7605_3_lut_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__25694),
            .in2(N__25368),
            .in3(N__25677),
            .lcout(\nx.n11941 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i675_3_lut_LC_7_21_1 .C_ON=1'b0;
    defparam \nx.mod_5_i675_3_lut_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i675_3_lut_LC_7_21_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i675_3_lut_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__25713),
            .in2(N__25731),
            .in3(N__25358),
            .lcout(\nx.n1008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9197_2_lut_LC_7_21_2 .C_ON=1'b0;
    defparam \nx.i9197_2_lut_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i9197_2_lut_LC_7_21_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \nx.i9197_2_lut_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25367),
            .in3(N__25676),
            .lcout(\nx.n1006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_25_LC_7_21_3 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_25_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_25_LC_7_21_3 .LUT_INIT=16'b1111110011111100;
    LogicCell40 \nx.i1_2_lut_adj_25_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__25580),
            .in2(N__25599),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\nx.n12837_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i604_4_lut_LC_7_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i604_4_lut_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i604_4_lut_LC_7_21_4 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \nx.mod_5_i604_4_lut_LC_7_21_4  (
            .in0(N__25563),
            .in1(_gnd_net_),
            .in2(N__25380),
            .in3(N__25807),
            .lcout(\nx.n905 ),
            .ltout(\nx.n905_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_44_LC_7_21_5 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_44_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_44_LC_7_21_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \nx.i1_4_lut_adj_44_LC_7_21_5  (
            .in0(N__25535),
            .in1(N__25657),
            .in2(N__25377),
            .in3(N__25374),
            .lcout(\nx.n11174 ),
            .ltout(\nx.n11174_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9198_1_lut_LC_7_21_6 .C_ON=1'b0;
    defparam \nx.i9198_1_lut_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9198_1_lut_LC_7_21_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \nx.i9198_1_lut_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25335),
            .in3(_gnd_net_),
            .lcout(\nx.n13594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i605_4_lut_LC_7_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_i605_4_lut_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i605_4_lut_LC_7_21_7 .LUT_INIT=16'b1010101010101001;
    LogicCell40 \nx.mod_5_i605_4_lut_LC_7_21_7  (
            .in0(N__25595),
            .in1(N__25579),
            .in2(N__25809),
            .in3(N__25562),
            .lcout(\nx.n906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_2_lut_LC_7_22_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_2_lut_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_2_lut_LC_7_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_2_lut_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__25327),
            .in2(_gnd_net_),
            .in3(N__25272),
            .lcout(\nx.n977 ),
            .ltout(),
            .carryin(bfn_7_22_0_),
            .carryout(\nx.n10738 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_3_lut_LC_7_22_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_3_lut_LC_7_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_3_lut_LC_7_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_3_lut_LC_7_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25730),
            .in3(N__25707),
            .lcout(\nx.n976 ),
            .ltout(),
            .carryin(\nx.n10738 ),
            .carryout(\nx.n10739 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_4_lut_LC_7_22_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_4_lut_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_4_lut_LC_7_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_4_lut_LC_7_22_2  (
            .in0(_gnd_net_),
            .in1(N__41616),
            .in2(N__25704),
            .in3(N__25680),
            .lcout(\nx.n975 ),
            .ltout(),
            .carryin(\nx.n10739 ),
            .carryout(\nx.n10740 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_5_lut_LC_7_22_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_5_lut_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_5_lut_LC_7_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_5_lut_LC_7_22_3  (
            .in0(_gnd_net_),
            .in1(N__41619),
            .in2(N__25539),
            .in3(N__25668),
            .lcout(\nx.n974 ),
            .ltout(),
            .carryin(\nx.n10740 ),
            .carryout(\nx.n10741 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_6_lut_LC_7_22_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_669_6_lut_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_6_lut_LC_7_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_669_6_lut_LC_7_22_4  (
            .in0(_gnd_net_),
            .in1(N__41617),
            .in2(N__25664),
            .in3(N__25635),
            .lcout(\nx.n973 ),
            .ltout(),
            .carryin(\nx.n10741 ),
            .carryout(\nx.n10742 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_669_7_lut_LC_7_22_5 .C_ON=1'b0;
    defparam \nx.mod_5_add_669_7_lut_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_669_7_lut_LC_7_22_5 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_669_7_lut_LC_7_22_5  (
            .in0(N__41618),
            .in1(N__25632),
            .in2(N__25626),
            .in3(N__25617),
            .lcout(\nx.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i538_3_lut_2_lut_LC_7_22_6 .C_ON=1'b0;
    defparam \nx.mod_5_i538_3_lut_2_lut_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i538_3_lut_2_lut_LC_7_22_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \nx.mod_5_i538_3_lut_2_lut_LC_7_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25855),
            .in3(N__25827),
            .lcout(\nx.n807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9153_3_lut_LC_7_22_7 .C_ON=1'b0;
    defparam \nx.i9153_3_lut_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.i9153_3_lut_LC_7_22_7 .LUT_INIT=16'b1111000011000011;
    LogicCell40 \nx.i9153_3_lut_LC_7_22_7  (
            .in0(_gnd_net_),
            .in1(N__25808),
            .in2(N__25581),
            .in3(N__25561),
            .lcout(\nx.n11868 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_137_LC_7_23_0 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_137_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_137_LC_7_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_137_LC_7_23_0  (
            .in0(N__35232),
            .in1(N__25522),
            .in2(N__25481),
            .in3(N__29328),
            .lcout(\nx.n44_adj_782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1665_3_lut_4_lut_LC_7_23_1 .C_ON=1'b0;
    defparam \nx.i1665_3_lut_4_lut_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1665_3_lut_4_lut_LC_7_23_1 .LUT_INIT=16'b1000001000001000;
    LogicCell40 \nx.i1665_3_lut_4_lut_LC_7_23_1  (
            .in0(N__25894),
            .in1(N__26073),
            .in2(N__26033),
            .in3(N__25985),
            .lcout(\nx.n11912 ),
            .ltout(\nx.n11912_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5757_2_lut_3_lut_4_lut_LC_7_23_2 .C_ON=1'b0;
    defparam \nx.i5757_2_lut_3_lut_4_lut_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.i5757_2_lut_3_lut_4_lut_LC_7_23_2 .LUT_INIT=16'b1101110111010111;
    LogicCell40 \nx.i5757_2_lut_3_lut_4_lut_LC_7_23_2  (
            .in0(N__25926),
            .in1(N__25895),
            .in2(N__26091),
            .in3(N__25828),
            .lcout(\nx.n58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6008_2_lut_4_lut_3_lut_LC_7_23_4 .C_ON=1'b0;
    defparam \nx.i6008_2_lut_4_lut_3_lut_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.i6008_2_lut_4_lut_3_lut_LC_7_23_4 .LUT_INIT=16'b0011100000111000;
    LogicCell40 \nx.i6008_2_lut_4_lut_3_lut_LC_7_23_4  (
            .in0(N__26074),
            .in1(N__26029),
            .in2(N__25989),
            .in3(_gnd_net_),
            .lcout(\nx.n9803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_adj_87_LC_7_23_5 .C_ON=1'b0;
    defparam \nx.i20_4_lut_adj_87_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_adj_87_LC_7_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i20_4_lut_adj_87_LC_7_23_5  (
            .in0(N__32975),
            .in1(N__33293),
            .in2(N__32847),
            .in3(N__32891),
            .lcout(\nx.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1940_2_lut_3_lut_4_lut_LC_7_23_6 .C_ON=1'b0;
    defparam \nx.i1940_2_lut_3_lut_4_lut_LC_7_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.i1940_2_lut_3_lut_4_lut_LC_7_23_6 .LUT_INIT=16'b0010001000101000;
    LogicCell40 \nx.i1940_2_lut_3_lut_4_lut_LC_7_23_6  (
            .in0(N__25927),
            .in1(N__25896),
            .in2(N__25857),
            .in3(N__25829),
            .lcout(\nx.n5703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_170_LC_7_24_0.C_ON=1'b0;
    defparam i2_4_lut_adj_170_LC_7_24_0.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_170_LC_7_24_0.LUT_INIT=16'b0110111111110110;
    LogicCell40 i2_4_lut_adj_170_LC_7_24_0 (
            .in0(N__25776),
            .in1(N__26127),
            .in2(N__25770),
            .in3(N__25737),
            .lcout(n10_adj_846),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i7_LC_7_24_1.C_ON=1'b0;
    defparam neopxl_color_prev_i7_LC_7_24_1.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i7_LC_7_24_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 neopxl_color_prev_i7_LC_7_24_1 (
            .in0(N__26129),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(neopxl_color_prev_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46879),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i15_LC_7_24_2.C_ON=1'b0;
    defparam neopxl_color_prev_i15_LC_7_24_2.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i15_LC_7_24_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 neopxl_color_prev_i15_LC_7_24_2 (
            .in0(N__25769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(neopxl_color_prev_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46879),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_7_24_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_7_24_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_7_24_3.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_2_lut_3_lut_LC_7_24_3 (
            .in0(N__26128),
            .in1(N__43897),
            .in2(_gnd_net_),
            .in3(N__47518),
            .lcout(n22_adj_793),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8978_3_lut_LC_7_24_5 .C_ON=1'b0;
    defparam \nx.i8978_3_lut_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.i8978_3_lut_LC_7_24_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.i8978_3_lut_LC_7_24_5  (
            .in0(N__26126),
            .in1(N__26208),
            .in2(_gnd_net_),
            .in3(N__26161),
            .lcout(\nx.n13373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_191_LC_7_24_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_191_LC_7_24_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_191_LC_7_24_6.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_2_lut_3_lut_adj_191_LC_7_24_6 (
            .in0(N__27293),
            .in1(N__43892),
            .in2(_gnd_net_),
            .in3(N__47514),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_194_LC_7_24_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_194_LC_7_24_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_194_LC_7_24_7.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_2_lut_3_lut_adj_194_LC_7_24_7 (
            .in0(N__32220),
            .in1(N__43896),
            .in2(_gnd_net_),
            .in3(N__47517),
            .lcout(n22_adj_787),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i7_LC_7_25_0.C_ON=1'b0;
    defparam neopxl_color_i7_LC_7_25_0.SEQ_MODE=4'b1001;
    defparam neopxl_color_i7_LC_7_25_0.LUT_INIT=16'b0000111100001000;
    LogicCell40 neopxl_color_i7_LC_7_25_0 (
            .in0(N__47539),
            .in1(N__43898),
            .in2(N__43715),
            .in3(N__26130),
            .lcout(neopxl_color_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46883),
            .ce(),
            .sr(N__26109));
    defparam \nx.i5_3_lut_LC_7_25_6 .C_ON=1'b0;
    defparam \nx.i5_3_lut_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.i5_3_lut_LC_7_25_6 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \nx.i5_3_lut_LC_7_25_6  (
            .in0(_gnd_net_),
            .in1(N__26348),
            .in2(N__26313),
            .in3(N__26653),
            .lcout(\nx.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1356_3_lut_LC_7_25_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1356_3_lut_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1356_3_lut_LC_7_25_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i1356_3_lut_LC_7_25_7  (
            .in0(N__26349),
            .in1(N__26325),
            .in2(_gnd_net_),
            .in3(N__27543),
            .lcout(\nx.n2009 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_27_LC_7_26_0 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_27_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_27_LC_7_26_0 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i1_2_lut_adj_27_LC_7_26_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26505),
            .in3(N__26543),
            .lcout(\nx.n16_adj_678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_26_LC_7_26_1 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_26_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_26_LC_7_26_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_26_LC_7_26_1  (
            .in0(N__27127),
            .in1(N__26248),
            .in2(N__27089),
            .in3(N__26275),
            .lcout(),
            .ltout(\nx.n26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_28_LC_7_26_2 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_28_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_28_LC_7_26_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_28_LC_7_26_2  (
            .in0(N__27601),
            .in1(N__27355),
            .in2(N__26100),
            .in3(N__26097),
            .lcout(),
            .ltout(\nx.n28_adj_679_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_29_LC_7_26_3 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_29_LC_7_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_29_LC_7_26_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_29_LC_7_26_3  (
            .in0(N__26416),
            .in1(N__26523),
            .in2(N__26367),
            .in3(N__26364),
            .lcout(\nx.n1928 ),
            .ltout(\nx.n1928_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1354_3_lut_LC_7_26_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1354_3_lut_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1354_3_lut_LC_7_26_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1354_3_lut_LC_7_26_4  (
            .in0(N__26276),
            .in1(_gnd_net_),
            .in2(N__26358),
            .in3(N__26259),
            .lcout(\nx.n2007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1352_3_lut_LC_7_26_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1352_3_lut_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1352_3_lut_LC_7_26_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1352_3_lut_LC_7_26_5  (
            .in0(N__26417),
            .in1(_gnd_net_),
            .in2(N__27545),
            .in3(N__26400),
            .lcout(\nx.n2005 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1353_3_lut_LC_7_26_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1353_3_lut_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1353_3_lut_LC_7_26_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1353_3_lut_LC_7_26_6  (
            .in0(N__26249),
            .in1(_gnd_net_),
            .in2(N__26232),
            .in3(N__27518),
            .lcout(\nx.n2006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1355_3_lut_LC_7_26_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1355_3_lut_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1355_3_lut_LC_7_26_7 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \nx.mod_5_i1355_3_lut_LC_7_26_7  (
            .in0(N__26308),
            .in1(N__26286),
            .in2(N__27544),
            .in3(_gnd_net_),
            .lcout(\nx.n2008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_2_lut_LC_7_27_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_2_lut_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_2_lut_LC_7_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_2_lut_LC_7_27_0  (
            .in0(_gnd_net_),
            .in1(N__26355),
            .in2(_gnd_net_),
            .in3(N__26316),
            .lcout(\nx.n1977 ),
            .ltout(),
            .carryin(bfn_7_27_0_),
            .carryout(\nx.n10833 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_3_lut_LC_7_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_3_lut_LC_7_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_3_lut_LC_7_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_3_lut_LC_7_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26309),
            .in3(N__26280),
            .lcout(\nx.n1976 ),
            .ltout(),
            .carryin(\nx.n10833 ),
            .carryout(\nx.n10834 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_4_lut_LC_7_27_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_4_lut_LC_7_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_4_lut_LC_7_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_4_lut_LC_7_27_2  (
            .in0(_gnd_net_),
            .in1(N__41627),
            .in2(N__26277),
            .in3(N__26253),
            .lcout(\nx.n1975 ),
            .ltout(),
            .carryin(\nx.n10834 ),
            .carryout(\nx.n10835 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_5_lut_LC_7_27_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_5_lut_LC_7_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_5_lut_LC_7_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_5_lut_LC_7_27_3  (
            .in0(_gnd_net_),
            .in1(N__41630),
            .in2(N__26250),
            .in3(N__26223),
            .lcout(\nx.n1974 ),
            .ltout(),
            .carryin(\nx.n10835 ),
            .carryout(\nx.n10836 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_6_lut_LC_7_27_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_6_lut_LC_7_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_6_lut_LC_7_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_6_lut_LC_7_27_4  (
            .in0(_gnd_net_),
            .in1(N__41628),
            .in2(N__26418),
            .in3(N__26394),
            .lcout(\nx.n1973 ),
            .ltout(),
            .carryin(\nx.n10836 ),
            .carryout(\nx.n10837 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_7_lut_LC_7_27_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_7_lut_LC_7_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_7_lut_LC_7_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_7_lut_LC_7_27_5  (
            .in0(_gnd_net_),
            .in1(N__41631),
            .in2(N__27088),
            .in3(N__26391),
            .lcout(\nx.n1972 ),
            .ltout(),
            .carryin(\nx.n10837 ),
            .carryout(\nx.n10838 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_8_lut_LC_7_27_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_8_lut_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_8_lut_LC_7_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_8_lut_LC_7_27_6  (
            .in0(_gnd_net_),
            .in1(N__41629),
            .in2(N__26654),
            .in3(N__26388),
            .lcout(\nx.n1971 ),
            .ltout(),
            .carryin(\nx.n10838 ),
            .carryout(\nx.n10839 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_9_lut_LC_7_27_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_9_lut_LC_7_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_9_lut_LC_7_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_9_lut_LC_7_27_7  (
            .in0(_gnd_net_),
            .in1(N__41632),
            .in2(N__27131),
            .in3(N__26385),
            .lcout(\nx.n1970 ),
            .ltout(),
            .carryin(\nx.n10839 ),
            .carryout(\nx.n10840 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_10_lut_LC_7_28_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_10_lut_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_10_lut_LC_7_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_10_lut_LC_7_28_0  (
            .in0(_gnd_net_),
            .in1(N__42201),
            .in2(N__27605),
            .in3(N__26382),
            .lcout(\nx.n1969 ),
            .ltout(),
            .carryin(bfn_7_28_0_),
            .carryout(\nx.n10841 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_11_lut_LC_7_28_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_11_lut_LC_7_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_11_lut_LC_7_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_11_lut_LC_7_28_1  (
            .in0(_gnd_net_),
            .in1(N__42205),
            .in2(N__27356),
            .in3(N__26379),
            .lcout(\nx.n1968 ),
            .ltout(),
            .carryin(\nx.n10841 ),
            .carryout(\nx.n10842 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_12_lut_LC_7_28_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_12_lut_LC_7_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_12_lut_LC_7_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_12_lut_LC_7_28_2  (
            .in0(_gnd_net_),
            .in1(N__42202),
            .in2(N__27170),
            .in3(N__26376),
            .lcout(\nx.n1967 ),
            .ltout(),
            .carryin(\nx.n10842 ),
            .carryout(\nx.n10843 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_13_lut_LC_7_28_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_13_lut_LC_7_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_13_lut_LC_7_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_13_lut_LC_7_28_3  (
            .in0(_gnd_net_),
            .in1(N__42206),
            .in2(N__27212),
            .in3(N__26373),
            .lcout(\nx.n1966 ),
            .ltout(),
            .carryin(\nx.n10843 ),
            .carryout(\nx.n10844 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_14_lut_LC_7_28_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_14_lut_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_14_lut_LC_7_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_14_lut_LC_7_28_4  (
            .in0(_gnd_net_),
            .in1(N__42203),
            .in2(N__26468),
            .in3(N__26370),
            .lcout(\nx.n1965 ),
            .ltout(),
            .carryin(\nx.n10844 ),
            .carryout(\nx.n10845 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_15_lut_LC_7_28_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_15_lut_LC_7_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_15_lut_LC_7_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_15_lut_LC_7_28_5  (
            .in0(_gnd_net_),
            .in1(N__42207),
            .in2(N__26436),
            .in3(N__26550),
            .lcout(\nx.n1964 ),
            .ltout(),
            .carryin(\nx.n10845 ),
            .carryout(\nx.n10846 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_16_lut_LC_7_28_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1339_16_lut_LC_7_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_16_lut_LC_7_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1339_16_lut_LC_7_28_6  (
            .in0(_gnd_net_),
            .in1(N__42204),
            .in2(N__26504),
            .in3(N__26547),
            .lcout(\nx.n1963 ),
            .ltout(),
            .carryin(\nx.n10846 ),
            .carryout(\nx.n10847 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1339_17_lut_LC_7_28_7 .C_ON=1'b0;
    defparam \nx.mod_5_add_1339_17_lut_LC_7_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1339_17_lut_LC_7_28_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \nx.mod_5_add_1339_17_lut_LC_7_28_7  (
            .in0(N__27552),
            .in1(N__42208),
            .in2(N__26544),
            .in3(N__26526),
            .lcout(\nx.n1994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_LC_7_29_1 .C_ON=1'b0;
    defparam \nx.i9_4_lut_LC_7_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_LC_7_29_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_LC_7_29_1  (
            .in0(N__27163),
            .in1(N__27205),
            .in2(N__26467),
            .in3(N__26431),
            .lcout(\nx.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1342_3_lut_LC_7_29_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1342_3_lut_LC_7_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1342_3_lut_LC_7_29_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \nx.mod_5_i1342_3_lut_LC_7_29_2  (
            .in0(_gnd_net_),
            .in1(N__27551),
            .in2(N__26514),
            .in3(N__26500),
            .lcout(\nx.n1995 ),
            .ltout(\nx.n1995_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9_4_lut_adj_33_LC_7_29_3 .C_ON=1'b0;
    defparam \nx.i9_4_lut_adj_33_LC_7_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.i9_4_lut_adj_33_LC_7_29_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i9_4_lut_adj_33_LC_7_29_3  (
            .in0(N__28964),
            .in1(N__29143),
            .in2(N__26478),
            .in3(N__27407),
            .lcout(\nx.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1344_3_lut_LC_7_29_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1344_3_lut_LC_7_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1344_3_lut_LC_7_29_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1344_3_lut_LC_7_29_4  (
            .in0(_gnd_net_),
            .in1(N__26475),
            .in2(N__26469),
            .in3(N__27546),
            .lcout(\nx.n1997 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1343_3_lut_LC_7_29_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1343_3_lut_LC_7_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1343_3_lut_LC_7_29_5 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \nx.mod_5_i1343_3_lut_LC_7_29_5  (
            .in0(N__26442),
            .in1(N__26432),
            .in2(N__27567),
            .in3(_gnd_net_),
            .lcout(\nx.n1996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1350_3_lut_LC_7_29_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1350_3_lut_LC_7_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1350_3_lut_LC_7_29_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1350_3_lut_LC_7_29_6  (
            .in0(_gnd_net_),
            .in1(N__26667),
            .in2(N__26658),
            .in3(N__27550),
            .lcout(\nx.n2003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8965_4_lut_LC_7_31_2.C_ON=1'b0;
    defparam i8965_4_lut_LC_7_31_2.SEQ_MODE=4'b0000;
    defparam i8965_4_lut_LC_7_31_2.LUT_INIT=16'b1011101000100010;
    LogicCell40 i8965_4_lut_LC_7_31_2 (
            .in0(N__27884),
            .in1(N__27815),
            .in2(N__27843),
            .in3(N__27863),
            .lcout(n13360),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8966_4_lut_LC_7_31_5.C_ON=1'b0;
    defparam i8966_4_lut_LC_7_31_5.SEQ_MODE=4'b0000;
    defparam i8966_4_lut_LC_7_31_5.LUT_INIT=16'b1111111011000100;
    LogicCell40 i8966_4_lut_LC_7_31_5 (
            .in0(N__27864),
            .in1(N__27842),
            .in2(N__27819),
            .in3(N__27885),
            .lcout(),
            .ltout(n13361_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8967_3_lut_LC_7_31_6.C_ON=1'b0;
    defparam i8967_3_lut_LC_7_31_6.SEQ_MODE=4'b0000;
    defparam i8967_3_lut_LC_7_31_6.LUT_INIT=16'b0000111101010101;
    LogicCell40 i8967_3_lut_LC_7_31_6 (
            .in0(N__26628),
            .in1(_gnd_net_),
            .in2(N__26622),
            .in3(N__27789),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_103_LC_9_17_1 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_103_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_103_LC_9_17_1 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \nx.i1_4_lut_adj_103_LC_9_17_1  (
            .in0(N__33483),
            .in1(N__33516),
            .in2(N__34024),
            .in3(N__27924),
            .lcout(\nx.n12817 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i12_LC_9_17_2.C_ON=1'b0;
    defparam neopxl_color_i12_LC_9_17_2.SEQ_MODE=4'b1000;
    defparam neopxl_color_i12_LC_9_17_2.LUT_INIT=16'b1111011100010000;
    LogicCell40 neopxl_color_i12_LC_9_17_2 (
            .in0(N__47598),
            .in1(N__43932),
            .in2(N__43691),
            .in3(N__26596),
            .lcout(neopxl_color_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46869),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2147_3_lut_LC_9_17_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2147_3_lut_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2147_3_lut_LC_9_17_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2147_3_lut_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__34131),
            .in2(N__34025),
            .in3(N__34098),
            .lcout(\nx.n59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9112_3_lut_LC_9_17_6 .C_ON=1'b0;
    defparam \nx.i9112_3_lut_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9112_3_lut_LC_9_17_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \nx.i9112_3_lut_LC_9_17_6  (
            .in0(N__30815),
            .in1(N__30747),
            .in2(_gnd_net_),
            .in3(N__26564),
            .lcout(\nx.color_bit_N_642_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2146_3_lut_LC_9_18_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2146_3_lut_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2146_3_lut_LC_9_18_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2146_3_lut_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__34047),
            .in2(N__34032),
            .in3(N__34080),
            .lcout(),
            .ltout(\nx.n61_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_106_LC_9_18_2 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_106_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_106_LC_9_18_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_106_LC_9_18_2  (
            .in0(N__26574),
            .in1(N__33861),
            .in2(N__26568),
            .in3(N__26676),
            .lcout(\nx.n11153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.state_i0_LC_9_18_5 .C_ON=1'b0;
    defparam \nx.state_i0_LC_9_18_5 .SEQ_MODE=4'b1001;
    defparam \nx.state_i0_LC_9_18_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \nx.state_i0_LC_9_18_5  (
            .in0(N__26880),
            .in1(N__26859),
            .in2(N__26823),
            .in3(N__26814),
            .lcout(state_0_adj_792),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46874),
            .ce(N__26715),
            .sr(N__26697));
    defparam \nx.i1_4_lut_adj_104_LC_9_18_6 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_104_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_104_LC_9_18_6 .LUT_INIT=16'b1111101111111000;
    LogicCell40 \nx.i1_4_lut_adj_104_LC_9_18_6  (
            .in0(N__33432),
            .in1(N__34027),
            .in2(N__26688),
            .in3(N__33468),
            .lcout(),
            .ltout(\nx.n12819_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_105_LC_9_18_7 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_105_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_105_LC_9_18_7 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \nx.i1_4_lut_adj_105_LC_9_18_7  (
            .in0(N__34028),
            .in1(N__33387),
            .in2(N__26679),
            .in3(N__33417),
            .lcout(\nx.n12821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2036_3_lut_LC_9_19_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2036_3_lut_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2036_3_lut_LC_9_19_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i2036_3_lut_LC_9_19_3  (
            .in0(N__35205),
            .in1(N__35259),
            .in2(_gnd_net_),
            .in3(N__37321),
            .lcout(\nx.n3009 ),
            .ltout(\nx.n3009_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_3_lut_LC_9_19_4 .C_ON=1'b0;
    defparam \nx.i13_3_lut_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.i13_3_lut_LC_9_19_4 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \nx.i13_3_lut_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__29338),
            .in2(N__26670),
            .in3(N__29227),
            .lcout(\nx.n39_adj_671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1967_3_lut_LC_9_19_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1967_3_lut_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1967_3_lut_LC_9_19_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1967_3_lut_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__28233),
            .in2(N__26910),
            .in3(N__37517),
            .lcout(\nx.n2908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1966_3_lut_LC_9_19_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1966_3_lut_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1966_3_lut_LC_9_19_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1966_3_lut_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__26895),
            .in2(N__37564),
            .in3(N__28082),
            .lcout(\nx.n2907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_66_LC_9_20_0 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_66_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_66_LC_9_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_66_LC_9_20_0  (
            .in0(N__37766),
            .in1(N__27046),
            .in2(N__27974),
            .in3(N__26981),
            .lcout(\nx.n38_adj_713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_117_LC_9_20_1 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_117_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_117_LC_9_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_117_LC_9_20_1  (
            .in0(N__37339),
            .in1(N__35449),
            .in2(N__35517),
            .in3(N__35401),
            .lcout(\nx.n42_adj_765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1899_3_lut_LC_9_20_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1899_3_lut_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1899_3_lut_LC_9_20_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1899_3_lut_LC_9_20_2  (
            .in0(N__28278),
            .in1(_gnd_net_),
            .in2(N__30009),
            .in3(N__31270),
            .lcout(\nx.n2808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1950_3_lut_LC_9_20_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1950_3_lut_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1950_3_lut_LC_9_20_3 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \nx.mod_5_i1950_3_lut_LC_9_20_3  (
            .in0(N__27047),
            .in1(N__27000),
            .in2(N__37595),
            .in3(_gnd_net_),
            .lcout(\nx.n2891 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1947_3_lut_LC_9_20_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1947_3_lut_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1947_3_lut_LC_9_20_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1947_3_lut_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__26955),
            .in2(N__28344),
            .in3(N__37556),
            .lcout(\nx.n2888 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1882_3_lut_LC_9_20_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1882_3_lut_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1882_3_lut_LC_9_20_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1882_3_lut_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__31574),
            .in2(N__31278),
            .in3(N__28458),
            .lcout(\nx.n2791 ),
            .ltout(\nx.n2791_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1949_3_lut_LC_9_20_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1949_3_lut_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1949_3_lut_LC_9_20_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1949_3_lut_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__26970),
            .in2(N__26916),
            .in3(N__37560),
            .lcout(\nx.n2890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_2_lut_LC_9_21_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_2_lut_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_2_lut_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_2_lut_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__28206),
            .in2(_gnd_net_),
            .in3(N__26913),
            .lcout(\nx.n2877 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\nx.n11004 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_3_lut_LC_9_21_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_3_lut_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_3_lut_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_3_lut_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__28229),
            .in2(_gnd_net_),
            .in3(N__26898),
            .lcout(\nx.n2876 ),
            .ltout(),
            .carryin(\nx.n11004 ),
            .carryout(\nx.n11005 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_4_lut_LC_9_21_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_4_lut_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_4_lut_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_4_lut_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__41742),
            .in2(N__28083),
            .in3(N__26886),
            .lcout(\nx.n2875 ),
            .ltout(),
            .carryin(\nx.n11005 ),
            .carryout(\nx.n11006 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_5_lut_LC_9_21_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_5_lut_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_5_lut_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_5_lut_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__41745),
            .in2(N__28031),
            .in3(N__26883),
            .lcout(\nx.n2874 ),
            .ltout(),
            .carryin(\nx.n11006 ),
            .carryout(\nx.n11007 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_6_lut_LC_9_21_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_6_lut_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_6_lut_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_6_lut_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__41743),
            .in2(N__34817),
            .in3(N__26943),
            .lcout(\nx.n2873 ),
            .ltout(),
            .carryin(\nx.n11007 ),
            .carryout(\nx.n11008 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_7_lut_LC_9_21_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_7_lut_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_7_lut_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_7_lut_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__41746),
            .in2(N__33844),
            .in3(N__26940),
            .lcout(\nx.n2872 ),
            .ltout(),
            .carryin(\nx.n11008 ),
            .carryout(\nx.n11009 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_8_lut_LC_9_21_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_8_lut_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_8_lut_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_8_lut_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__41744),
            .in2(N__36845),
            .in3(N__26937),
            .lcout(\nx.n2871 ),
            .ltout(),
            .carryin(\nx.n11009 ),
            .carryout(\nx.n11010 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_9_lut_LC_9_21_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_9_lut_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_9_lut_LC_9_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_9_lut_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__41747),
            .in2(N__34172),
            .in3(N__26934),
            .lcout(\nx.n2870 ),
            .ltout(),
            .carryin(\nx.n11010 ),
            .carryout(\nx.n11011 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_10_lut_LC_9_22_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_10_lut_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_10_lut_LC_9_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_10_lut_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__41935),
            .in2(N__28161),
            .in3(N__26931),
            .lcout(\nx.n2869 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\nx.n11012 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_11_lut_LC_9_22_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_11_lut_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_11_lut_LC_9_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_11_lut_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__41811),
            .in2(N__28108),
            .in3(N__26928),
            .lcout(\nx.n2868 ),
            .ltout(),
            .carryin(\nx.n11012 ),
            .carryout(\nx.n11013 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_12_lut_LC_9_22_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_12_lut_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_12_lut_LC_9_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_12_lut_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__41936),
            .in2(N__29774),
            .in3(N__26925),
            .lcout(\nx.n2867 ),
            .ltout(),
            .carryin(\nx.n11013 ),
            .carryout(\nx.n11014 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_13_lut_LC_9_22_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_13_lut_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_13_lut_LC_9_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_13_lut_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__41812),
            .in2(N__31440),
            .in3(N__26922),
            .lcout(\nx.n2866 ),
            .ltout(),
            .carryin(\nx.n11014 ),
            .carryout(\nx.n11015 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_14_lut_LC_9_22_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_14_lut_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_14_lut_LC_9_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_14_lut_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__41937),
            .in2(N__33804),
            .in3(N__26919),
            .lcout(\nx.n2865 ),
            .ltout(),
            .carryin(\nx.n11015 ),
            .carryout(\nx.n11016 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_15_lut_LC_9_22_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_15_lut_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_15_lut_LC_9_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_15_lut_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__41813),
            .in2(N__34882),
            .in3(N__27015),
            .lcout(\nx.n2864 ),
            .ltout(),
            .carryin(\nx.n11016 ),
            .carryout(\nx.n11017 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_16_lut_LC_9_22_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_16_lut_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_16_lut_LC_9_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_16_lut_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__41938),
            .in2(N__31143),
            .in3(N__27012),
            .lcout(\nx.n2863 ),
            .ltout(),
            .carryin(\nx.n11017 ),
            .carryout(\nx.n11018 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_17_lut_LC_9_22_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_17_lut_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_17_lut_LC_9_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_17_lut_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(N__41814),
            .in2(N__28136),
            .in3(N__27009),
            .lcout(\nx.n2862 ),
            .ltout(),
            .carryin(\nx.n11018 ),
            .carryout(\nx.n11019 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_18_lut_LC_9_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_18_lut_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_18_lut_LC_9_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_18_lut_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__41939),
            .in2(N__37654),
            .in3(N__27006),
            .lcout(\nx.n2861 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\nx.n11020 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_19_lut_LC_9_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_19_lut_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_19_lut_LC_9_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_19_lut_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__37762),
            .in2(N__42187),
            .in3(N__27003),
            .lcout(\nx.n2860 ),
            .ltout(),
            .carryin(\nx.n11020 ),
            .carryout(\nx.n11021 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_20_lut_LC_9_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_20_lut_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_20_lut_LC_9_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_20_lut_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__41943),
            .in2(N__27048),
            .in3(N__26991),
            .lcout(\nx.n2859 ),
            .ltout(),
            .carryin(\nx.n11021 ),
            .carryout(\nx.n11022 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_21_lut_LC_9_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_21_lut_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_21_lut_LC_9_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_21_lut_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__41805),
            .in2(N__26988),
            .in3(N__26961),
            .lcout(\nx.n2858 ),
            .ltout(),
            .carryin(\nx.n11022 ),
            .carryout(\nx.n11023 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_22_lut_LC_9_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_22_lut_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_22_lut_LC_9_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_22_lut_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__41944),
            .in2(N__27970),
            .in3(N__26958),
            .lcout(\nx.n2857 ),
            .ltout(),
            .carryin(\nx.n11023 ),
            .carryout(\nx.n11024 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_23_lut_LC_9_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_23_lut_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_23_lut_LC_9_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_23_lut_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__41806),
            .in2(N__28340),
            .in3(N__26946),
            .lcout(\nx.n2856 ),
            .ltout(),
            .carryin(\nx.n11024 ),
            .carryout(\nx.n11025 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_24_lut_LC_9_23_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_24_lut_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_24_lut_LC_9_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_24_lut_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__31331),
            .in2(N__42071),
            .in3(N__27057),
            .lcout(\nx.n2855 ),
            .ltout(),
            .carryin(\nx.n11025 ),
            .carryout(\nx.n11026 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_25_lut_LC_9_23_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1942_25_lut_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_25_lut_LC_9_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1942_25_lut_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__41810),
            .in2(N__29946),
            .in3(N__27054),
            .lcout(\nx.n2854 ),
            .ltout(),
            .carryin(\nx.n11026 ),
            .carryout(\nx.n11027 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1942_26_lut_LC_9_24_0 .C_ON=1'b0;
    defparam \nx.mod_5_add_1942_26_lut_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1942_26_lut_LC_9_24_0 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_1942_26_lut_LC_9_24_0  (
            .in0(N__42060),
            .in1(N__37596),
            .in2(N__28608),
            .in3(N__27051),
            .lcout(\nx.n2885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1885_3_lut_LC_9_24_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1885_3_lut_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1885_3_lut_LC_9_24_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1885_3_lut_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__31667),
            .in2(N__28488),
            .in3(N__31269),
            .lcout(\nx.n2794 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1892_3_lut_LC_9_24_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1892_3_lut_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1892_3_lut_LC_9_24_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1892_3_lut_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__28380),
            .in2(N__31277),
            .in3(N__34209),
            .lcout(\nx.n2801 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1880_3_lut_LC_9_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1880_3_lut_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1880_3_lut_LC_9_24_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1880_3_lut_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__31268),
            .in2(N__31611),
            .in3(N__28434),
            .lcout(\nx.n2789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1881_3_lut_LC_9_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1881_3_lut_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1881_3_lut_LC_9_24_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1881_3_lut_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(N__31637),
            .in2(N__31276),
            .in3(N__28443),
            .lcout(\nx.n2790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1883_3_lut_LC_9_24_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1883_3_lut_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1883_3_lut_LC_9_24_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1883_3_lut_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(N__31261),
            .in2(N__30087),
            .in3(N__28467),
            .lcout(\nx.n2792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_prev_i5_LC_9_24_6.C_ON=1'b0;
    defparam neopxl_color_prev_i5_LC_9_24_6.SEQ_MODE=4'b1000;
    defparam neopxl_color_prev_i5_LC_9_24_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 neopxl_color_prev_i5_LC_9_24_6 (
            .in0(N__27271),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(neopxl_color_prev_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46886),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1884_3_lut_LC_9_24_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1884_3_lut_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1884_3_lut_LC_9_24_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1884_3_lut_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(N__31260),
            .in2(N__30066),
            .in3(N__28476),
            .lcout(\nx.n2793 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i5_LC_9_25_0.C_ON=1'b0;
    defparam neopxl_color_i5_LC_9_25_0.SEQ_MODE=4'b1001;
    defparam neopxl_color_i5_LC_9_25_0.LUT_INIT=16'b0011001100100000;
    LogicCell40 neopxl_color_i5_LC_9_25_0 (
            .in0(N__43951),
            .in1(N__43716),
            .in2(N__47696),
            .in3(N__27270),
            .lcout(neopxl_color_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46891),
            .ce(),
            .sr(N__27243));
    defparam \nx.mod_5_i1345_3_lut_LC_9_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1345_3_lut_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1345_3_lut_LC_9_25_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1345_3_lut_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__27228),
            .in2(N__27582),
            .in3(N__27216),
            .lcout(\nx.n1998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1346_3_lut_LC_9_25_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1346_3_lut_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1346_3_lut_LC_9_25_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1346_3_lut_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__27189),
            .in2(N__27177),
            .in3(N__27576),
            .lcout(\nx.n1999 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1349_3_lut_LC_9_25_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1349_3_lut_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1349_3_lut_LC_9_25_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1349_3_lut_LC_9_25_3  (
            .in0(_gnd_net_),
            .in1(N__27147),
            .in2(N__27581),
            .in3(N__27135),
            .lcout(\nx.n2002 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1351_3_lut_LC_9_25_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1351_3_lut_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1351_3_lut_LC_9_25_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1351_3_lut_LC_9_25_4  (
            .in0(_gnd_net_),
            .in1(N__27108),
            .in2(N__27096),
            .in3(N__27572),
            .lcout(\nx.n2004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1547_3_lut_LC_9_25_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1547_3_lut_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1547_3_lut_LC_9_25_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1547_3_lut_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(N__30213),
            .in2(N__32304),
            .in3(N__32579),
            .lcout(\nx.n2296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_2_lut_LC_9_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_2_lut_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_2_lut_LC_9_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_2_lut_LC_9_26_0  (
            .in0(_gnd_net_),
            .in1(N__28929),
            .in2(_gnd_net_),
            .in3(N__27063),
            .lcout(\nx.n2077 ),
            .ltout(),
            .carryin(bfn_9_26_0_),
            .carryout(\nx.n10848 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_3_lut_LC_9_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_3_lut_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_3_lut_LC_9_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_3_lut_LC_9_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29204),
            .in3(N__27060),
            .lcout(\nx.n2076 ),
            .ltout(),
            .carryin(\nx.n10848 ),
            .carryout(\nx.n10849 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_4_lut_LC_9_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_4_lut_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_4_lut_LC_9_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_4_lut_LC_9_26_2  (
            .in0(_gnd_net_),
            .in1(N__42086),
            .in2(N__29020),
            .in3(N__27321),
            .lcout(\nx.n2075 ),
            .ltout(),
            .carryin(\nx.n10849 ),
            .carryout(\nx.n10850 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_5_lut_LC_9_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_5_lut_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_5_lut_LC_9_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_5_lut_LC_9_26_3  (
            .in0(_gnd_net_),
            .in1(N__42061),
            .in2(N__28869),
            .in3(N__27318),
            .lcout(\nx.n2074 ),
            .ltout(),
            .carryin(\nx.n10850 ),
            .carryout(\nx.n10851 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_6_lut_LC_9_26_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_6_lut_LC_9_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_6_lut_LC_9_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_6_lut_LC_9_26_4  (
            .in0(_gnd_net_),
            .in1(N__42087),
            .in2(N__28711),
            .in3(N__27315),
            .lcout(\nx.n2073 ),
            .ltout(),
            .carryin(\nx.n10851 ),
            .carryout(\nx.n10852 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_7_lut_LC_9_26_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_7_lut_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_7_lut_LC_9_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_7_lut_LC_9_26_5  (
            .in0(_gnd_net_),
            .in1(N__42062),
            .in2(N__28679),
            .in3(N__27312),
            .lcout(\nx.n2072 ),
            .ltout(),
            .carryin(\nx.n10852 ),
            .carryout(\nx.n10853 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_8_lut_LC_9_26_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_8_lut_LC_9_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_8_lut_LC_9_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_8_lut_LC_9_26_6  (
            .in0(_gnd_net_),
            .in1(N__42088),
            .in2(N__28790),
            .in3(N__27309),
            .lcout(\nx.n2071 ),
            .ltout(),
            .carryin(\nx.n10853 ),
            .carryout(\nx.n10854 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_9_lut_LC_9_26_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_9_lut_LC_9_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_9_lut_LC_9_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_9_lut_LC_9_26_7  (
            .in0(_gnd_net_),
            .in1(N__42063),
            .in2(N__28848),
            .in3(N__27306),
            .lcout(\nx.n2070 ),
            .ltout(),
            .carryin(\nx.n10854 ),
            .carryout(\nx.n10855 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_10_lut_LC_9_27_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_10_lut_LC_9_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_10_lut_LC_9_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_10_lut_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__42089),
            .in2(N__28644),
            .in3(N__27303),
            .lcout(\nx.n2069 ),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\nx.n10856 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_11_lut_LC_9_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_11_lut_LC_9_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_11_lut_LC_9_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_11_lut_LC_9_27_1  (
            .in0(_gnd_net_),
            .in1(N__42064),
            .in2(N__28554),
            .in3(N__27300),
            .lcout(\nx.n2068 ),
            .ltout(),
            .carryin(\nx.n10856 ),
            .carryout(\nx.n10857 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_12_lut_LC_9_27_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_12_lut_LC_9_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_12_lut_LC_9_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_12_lut_LC_9_27_2  (
            .in0(_gnd_net_),
            .in1(N__42090),
            .in2(N__28821),
            .in3(N__27297),
            .lcout(\nx.n2067 ),
            .ltout(),
            .carryin(\nx.n10857 ),
            .carryout(\nx.n10858 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_13_lut_LC_9_27_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_13_lut_LC_9_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_13_lut_LC_9_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_13_lut_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(N__42065),
            .in2(N__28530),
            .in3(N__27426),
            .lcout(\nx.n2066 ),
            .ltout(),
            .carryin(\nx.n10858 ),
            .carryout(\nx.n10859 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_14_lut_LC_9_27_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_14_lut_LC_9_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_14_lut_LC_9_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_14_lut_LC_9_27_4  (
            .in0(_gnd_net_),
            .in1(N__42091),
            .in2(N__28755),
            .in3(N__27423),
            .lcout(\nx.n2065 ),
            .ltout(),
            .carryin(\nx.n10859 ),
            .carryout(\nx.n10860 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_15_lut_LC_9_27_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_15_lut_LC_9_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_15_lut_LC_9_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_15_lut_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(N__42066),
            .in2(N__28982),
            .in3(N__27420),
            .lcout(\nx.n2064 ),
            .ltout(),
            .carryin(\nx.n10860 ),
            .carryout(\nx.n10861 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_16_lut_LC_9_27_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_16_lut_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_16_lut_LC_9_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_16_lut_LC_9_27_6  (
            .in0(_gnd_net_),
            .in1(N__42092),
            .in2(N__29157),
            .in3(N__27417),
            .lcout(\nx.n2063 ),
            .ltout(),
            .carryin(\nx.n10861 ),
            .carryout(\nx.n10862 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_17_lut_LC_9_27_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1406_17_lut_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_17_lut_LC_9_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1406_17_lut_LC_9_27_7  (
            .in0(_gnd_net_),
            .in1(N__42067),
            .in2(N__27392),
            .in3(N__27414),
            .lcout(\nx.n2062 ),
            .ltout(),
            .carryin(\nx.n10862 ),
            .carryout(\nx.n10863 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1406_18_lut_LC_9_28_0 .C_ON=1'b0;
    defparam \nx.mod_5_add_1406_18_lut_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1406_18_lut_LC_9_28_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1406_18_lut_LC_9_28_0  (
            .in0(N__42216),
            .in1(N__27411),
            .in2(N__29125),
            .in3(N__27396),
            .lcout(\nx.n2093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1409_3_lut_LC_9_28_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1409_3_lut_LC_9_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1409_3_lut_LC_9_28_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1409_3_lut_LC_9_28_1  (
            .in0(_gnd_net_),
            .in1(N__29112),
            .in2(N__27393),
            .in3(N__27366),
            .lcout(\nx.n2094 ),
            .ltout(\nx.n2094_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_35_LC_9_28_2 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_35_LC_9_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_35_LC_9_28_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i1_2_lut_adj_35_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27360),
            .in3(N__30854),
            .lcout(\nx.n18_adj_682 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1347_3_lut_LC_9_28_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1347_3_lut_LC_9_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1347_3_lut_LC_9_28_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1347_3_lut_LC_9_28_3  (
            .in0(_gnd_net_),
            .in1(N__27357),
            .in2(N__27580),
            .in3(N__27330),
            .lcout(\nx.n2000 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1348_3_lut_LC_9_28_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1348_3_lut_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1348_3_lut_LC_9_28_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1348_3_lut_LC_9_28_4  (
            .in0(_gnd_net_),
            .in1(N__27621),
            .in2(N__27612),
            .in3(N__27568),
            .lcout(\nx.n2001 ),
            .ltout(\nx.n2001_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1415_3_lut_LC_9_28_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1415_3_lut_LC_9_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1415_3_lut_LC_9_28_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1415_3_lut_LC_9_28_5  (
            .in0(_gnd_net_),
            .in1(N__27489),
            .in2(N__27483),
            .in3(N__29111),
            .lcout(\nx.n2100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1414_3_lut_LC_9_28_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1414_3_lut_LC_9_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1414_3_lut_LC_9_28_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1414_3_lut_LC_9_28_6  (
            .in0(_gnd_net_),
            .in1(N__28819),
            .in2(N__29126),
            .in3(N__27480),
            .lcout(\nx.n2099 ),
            .ltout(\nx.n2099_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_38_LC_9_28_7 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_38_LC_9_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_38_LC_9_28_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_38_LC_9_28_7  (
            .in0(N__30337),
            .in1(N__36580),
            .in2(N__27474),
            .in3(N__30712),
            .lcout(\nx.n28_adj_686 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i0_LC_9_29_0.C_ON=1'b1;
    defparam blink_counter_635__i0_LC_9_29_0.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i0_LC_9_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i0_LC_9_29_0 (
            .in0(_gnd_net_),
            .in1(N__27471),
            .in2(_gnd_net_),
            .in3(N__27465),
            .lcout(n26_adj_798),
            .ltout(),
            .carryin(bfn_9_29_0_),
            .carryout(n10644),
            .clk(N__46913),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i1_LC_9_29_1.C_ON=1'b1;
    defparam blink_counter_635__i1_LC_9_29_1.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i1_LC_9_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i1_LC_9_29_1 (
            .in0(_gnd_net_),
            .in1(N__27462),
            .in2(_gnd_net_),
            .in3(N__27456),
            .lcout(n25),
            .ltout(),
            .carryin(n10644),
            .carryout(n10645),
            .clk(N__46913),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i2_LC_9_29_2.C_ON=1'b1;
    defparam blink_counter_635__i2_LC_9_29_2.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i2_LC_9_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i2_LC_9_29_2 (
            .in0(_gnd_net_),
            .in1(N__27453),
            .in2(_gnd_net_),
            .in3(N__27447),
            .lcout(n24),
            .ltout(),
            .carryin(n10645),
            .carryout(n10646),
            .clk(N__46913),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i3_LC_9_29_3.C_ON=1'b1;
    defparam blink_counter_635__i3_LC_9_29_3.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i3_LC_9_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i3_LC_9_29_3 (
            .in0(_gnd_net_),
            .in1(N__27444),
            .in2(_gnd_net_),
            .in3(N__27438),
            .lcout(n23),
            .ltout(),
            .carryin(n10646),
            .carryout(n10647),
            .clk(N__46913),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i4_LC_9_29_4.C_ON=1'b1;
    defparam blink_counter_635__i4_LC_9_29_4.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i4_LC_9_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i4_LC_9_29_4 (
            .in0(_gnd_net_),
            .in1(N__27435),
            .in2(_gnd_net_),
            .in3(N__27429),
            .lcout(n22_adj_799),
            .ltout(),
            .carryin(n10647),
            .carryout(n10648),
            .clk(N__46913),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i5_LC_9_29_5.C_ON=1'b1;
    defparam blink_counter_635__i5_LC_9_29_5.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i5_LC_9_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i5_LC_9_29_5 (
            .in0(_gnd_net_),
            .in1(N__27693),
            .in2(_gnd_net_),
            .in3(N__27687),
            .lcout(n21),
            .ltout(),
            .carryin(n10648),
            .carryout(n10649),
            .clk(N__46913),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i6_LC_9_29_6.C_ON=1'b1;
    defparam blink_counter_635__i6_LC_9_29_6.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i6_LC_9_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i6_LC_9_29_6 (
            .in0(_gnd_net_),
            .in1(N__27684),
            .in2(_gnd_net_),
            .in3(N__27678),
            .lcout(n20),
            .ltout(),
            .carryin(n10649),
            .carryout(n10650),
            .clk(N__46913),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i7_LC_9_29_7.C_ON=1'b1;
    defparam blink_counter_635__i7_LC_9_29_7.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i7_LC_9_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i7_LC_9_29_7 (
            .in0(_gnd_net_),
            .in1(N__27675),
            .in2(_gnd_net_),
            .in3(N__27669),
            .lcout(n19_adj_800),
            .ltout(),
            .carryin(n10650),
            .carryout(n10651),
            .clk(N__46913),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i8_LC_9_30_0.C_ON=1'b1;
    defparam blink_counter_635__i8_LC_9_30_0.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i8_LC_9_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i8_LC_9_30_0 (
            .in0(_gnd_net_),
            .in1(N__27666),
            .in2(_gnd_net_),
            .in3(N__27660),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_9_30_0_),
            .carryout(n10652),
            .clk(N__46915),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i9_LC_9_30_1.C_ON=1'b1;
    defparam blink_counter_635__i9_LC_9_30_1.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i9_LC_9_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i9_LC_9_30_1 (
            .in0(_gnd_net_),
            .in1(N__27657),
            .in2(_gnd_net_),
            .in3(N__27651),
            .lcout(n17),
            .ltout(),
            .carryin(n10652),
            .carryout(n10653),
            .clk(N__46915),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i10_LC_9_30_2.C_ON=1'b1;
    defparam blink_counter_635__i10_LC_9_30_2.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i10_LC_9_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i10_LC_9_30_2 (
            .in0(_gnd_net_),
            .in1(N__27648),
            .in2(_gnd_net_),
            .in3(N__27642),
            .lcout(n16),
            .ltout(),
            .carryin(n10653),
            .carryout(n10654),
            .clk(N__46915),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i11_LC_9_30_3.C_ON=1'b1;
    defparam blink_counter_635__i11_LC_9_30_3.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i11_LC_9_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i11_LC_9_30_3 (
            .in0(_gnd_net_),
            .in1(N__27639),
            .in2(_gnd_net_),
            .in3(N__27633),
            .lcout(n15),
            .ltout(),
            .carryin(n10654),
            .carryout(n10655),
            .clk(N__46915),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i12_LC_9_30_4.C_ON=1'b1;
    defparam blink_counter_635__i12_LC_9_30_4.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i12_LC_9_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i12_LC_9_30_4 (
            .in0(_gnd_net_),
            .in1(N__27630),
            .in2(_gnd_net_),
            .in3(N__27624),
            .lcout(n14_adj_802),
            .ltout(),
            .carryin(n10655),
            .carryout(n10656),
            .clk(N__46915),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i13_LC_9_30_5.C_ON=1'b1;
    defparam blink_counter_635__i13_LC_9_30_5.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i13_LC_9_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i13_LC_9_30_5 (
            .in0(_gnd_net_),
            .in1(N__27765),
            .in2(_gnd_net_),
            .in3(N__27759),
            .lcout(n13),
            .ltout(),
            .carryin(n10656),
            .carryout(n10657),
            .clk(N__46915),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i14_LC_9_30_6.C_ON=1'b1;
    defparam blink_counter_635__i14_LC_9_30_6.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i14_LC_9_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i14_LC_9_30_6 (
            .in0(_gnd_net_),
            .in1(N__27756),
            .in2(_gnd_net_),
            .in3(N__27750),
            .lcout(n12),
            .ltout(),
            .carryin(n10657),
            .carryout(n10658),
            .clk(N__46915),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i15_LC_9_30_7.C_ON=1'b1;
    defparam blink_counter_635__i15_LC_9_30_7.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i15_LC_9_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i15_LC_9_30_7 (
            .in0(_gnd_net_),
            .in1(N__27747),
            .in2(_gnd_net_),
            .in3(N__27741),
            .lcout(n11),
            .ltout(),
            .carryin(n10658),
            .carryout(n10659),
            .clk(N__46915),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i16_LC_9_31_0.C_ON=1'b1;
    defparam blink_counter_635__i16_LC_9_31_0.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i16_LC_9_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i16_LC_9_31_0 (
            .in0(_gnd_net_),
            .in1(N__27738),
            .in2(_gnd_net_),
            .in3(N__27732),
            .lcout(n10_adj_806),
            .ltout(),
            .carryin(bfn_9_31_0_),
            .carryout(n10660),
            .clk(N__46921),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i17_LC_9_31_1.C_ON=1'b1;
    defparam blink_counter_635__i17_LC_9_31_1.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i17_LC_9_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i17_LC_9_31_1 (
            .in0(_gnd_net_),
            .in1(N__27729),
            .in2(_gnd_net_),
            .in3(N__27723),
            .lcout(n9_adj_807),
            .ltout(),
            .carryin(n10660),
            .carryout(n10661),
            .clk(N__46921),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i18_LC_9_31_2.C_ON=1'b1;
    defparam blink_counter_635__i18_LC_9_31_2.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i18_LC_9_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i18_LC_9_31_2 (
            .in0(_gnd_net_),
            .in1(N__27720),
            .in2(_gnd_net_),
            .in3(N__27714),
            .lcout(n8),
            .ltout(),
            .carryin(n10661),
            .carryout(n10662),
            .clk(N__46921),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i19_LC_9_31_3.C_ON=1'b1;
    defparam blink_counter_635__i19_LC_9_31_3.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i19_LC_9_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i19_LC_9_31_3 (
            .in0(_gnd_net_),
            .in1(N__27711),
            .in2(_gnd_net_),
            .in3(N__27705),
            .lcout(n7_adj_808),
            .ltout(),
            .carryin(n10662),
            .carryout(n10663),
            .clk(N__46921),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i20_LC_9_31_4.C_ON=1'b1;
    defparam blink_counter_635__i20_LC_9_31_4.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i20_LC_9_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i20_LC_9_31_4 (
            .in0(_gnd_net_),
            .in1(N__27702),
            .in2(_gnd_net_),
            .in3(N__27696),
            .lcout(n6_adj_809),
            .ltout(),
            .carryin(n10663),
            .carryout(n10664),
            .clk(N__46921),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i21_LC_9_31_5.C_ON=1'b1;
    defparam blink_counter_635__i21_LC_9_31_5.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i21_LC_9_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i21_LC_9_31_5 (
            .in0(_gnd_net_),
            .in1(N__27878),
            .in2(_gnd_net_),
            .in3(N__27867),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n10664),
            .carryout(n10665),
            .clk(N__46921),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i22_LC_9_31_6.C_ON=1'b1;
    defparam blink_counter_635__i22_LC_9_31_6.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i22_LC_9_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i22_LC_9_31_6 (
            .in0(_gnd_net_),
            .in1(N__27857),
            .in2(_gnd_net_),
            .in3(N__27846),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n10665),
            .carryout(n10666),
            .clk(N__46921),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i23_LC_9_31_7.C_ON=1'b1;
    defparam blink_counter_635__i23_LC_9_31_7.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i23_LC_9_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i23_LC_9_31_7 (
            .in0(_gnd_net_),
            .in1(N__27833),
            .in2(_gnd_net_),
            .in3(N__27822),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n10666),
            .carryout(n10667),
            .clk(N__46921),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i24_LC_9_32_0.C_ON=1'b1;
    defparam blink_counter_635__i24_LC_9_32_0.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i24_LC_9_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i24_LC_9_32_0 (
            .in0(_gnd_net_),
            .in1(N__27806),
            .in2(_gnd_net_),
            .in3(N__27795),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_9_32_0_),
            .carryout(n10668),
            .clk(N__46923),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_635__i25_LC_9_32_1.C_ON=1'b0;
    defparam blink_counter_635__i25_LC_9_32_1.SEQ_MODE=4'b1000;
    defparam blink_counter_635__i25_LC_9_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_635__i25_LC_9_32_1 (
            .in0(_gnd_net_),
            .in1(N__27782),
            .in2(_gnd_net_),
            .in3(N__27792),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46923),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_96_LC_10_17_0 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_96_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_96_LC_10_17_0 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \nx.i1_4_lut_adj_96_LC_10_17_0  (
            .in0(N__32943),
            .in1(N__32962),
            .in2(N__34006),
            .in3(N__30945),
            .lcout(\nx.n12775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2154_3_lut_LC_10_17_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2154_3_lut_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2154_3_lut_LC_10_17_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2154_3_lut_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__33663),
            .in2(N__33692),
            .in3(N__33984),
            .lcout(),
            .ltout(\nx.n45_adj_754_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_99_LC_10_17_2 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_99_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_99_LC_10_17_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_99_LC_10_17_2  (
            .in0(N__27918),
            .in1(N__30759),
            .in2(N__27771),
            .in3(N__27897),
            .lcout(),
            .ltout(\nx.n12809_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_100_LC_10_17_3 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_100_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_100_LC_10_17_3 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \nx.i1_4_lut_adj_100_LC_10_17_3  (
            .in0(N__33618),
            .in1(N__33648),
            .in2(N__27768),
            .in3(N__33985),
            .lcout(),
            .ltout(\nx.n12811_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_101_LC_10_17_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_101_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_101_LC_10_17_4 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \nx.i1_4_lut_adj_101_LC_10_17_4  (
            .in0(N__33986),
            .in1(N__33573),
            .in2(N__27930),
            .in3(N__33603),
            .lcout(),
            .ltout(\nx.n12813_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_102_LC_10_17_5 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_102_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_102_LC_10_17_5 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \nx.i1_4_lut_adj_102_LC_10_17_5  (
            .in0(N__33531),
            .in1(N__33554),
            .in2(N__27927),
            .in3(N__33987),
            .lcout(\nx.n12815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2155_3_lut_LC_10_17_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2155_3_lut_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2155_3_lut_LC_10_17_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2155_3_lut_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__33085),
            .in2(N__34007),
            .in3(N__33708),
            .lcout(\nx.n43_adj_753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_80_LC_10_18_0 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_80_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_80_LC_10_18_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_80_LC_10_18_0  (
            .in0(N__33238),
            .in1(N__33043),
            .in2(N__33205),
            .in3(N__32923),
            .lcout(),
            .ltout(\nx.n46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i23_4_lut_LC_10_18_1 .C_ON=1'b0;
    defparam \nx.i23_4_lut_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.i23_4_lut_LC_10_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i23_4_lut_LC_10_18_1  (
            .in0(N__32794),
            .in1(N__33361),
            .in2(N__27912),
            .in3(N__27891),
            .lcout(\nx.n50_adj_742 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2170_3_lut_LC_10_18_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2170_3_lut_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2170_3_lut_LC_10_18_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2170_3_lut_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__33027),
            .in2(N__33050),
            .in3(N__33988),
            .lcout(),
            .ltout(\nx.n13_adj_743_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_94_LC_10_18_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_94_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_94_LC_10_18_4 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \nx.i1_4_lut_adj_94_LC_10_18_4  (
            .in0(N__33989),
            .in1(N__33264),
            .in2(N__27909),
            .in3(N__33286),
            .lcout(),
            .ltout(\nx.n12787_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_98_LC_10_18_5 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_98_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_98_LC_10_18_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_98_LC_10_18_5  (
            .in0(N__30933),
            .in1(N__27906),
            .in2(N__27900),
            .in3(N__30960),
            .lcout(\nx.n12803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i8_3_lut_adj_81_LC_10_18_6 .C_ON=1'b0;
    defparam \nx.i8_3_lut_adj_81_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.i8_3_lut_adj_81_LC_10_18_6 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \nx.i8_3_lut_adj_81_LC_10_18_6  (
            .in0(N__32399),
            .in1(_gnd_net_),
            .in2(N__32353),
            .in3(N__33004),
            .lcout(\nx.n35_adj_738 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2035_3_lut_LC_10_19_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2035_3_lut_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2035_3_lut_LC_10_19_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2035_3_lut_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__35186),
            .in2(N__37322),
            .in3(N__35166),
            .lcout(\nx.n3008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2014_3_lut_LC_10_19_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2014_3_lut_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2014_3_lut_LC_10_19_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2014_3_lut_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__35611),
            .in2(N__35589),
            .in3(N__37311),
            .lcout(\nx.n2987 ),
            .ltout(\nx.n2987_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_LC_10_19_2 .C_ON=1'b0;
    defparam \nx.i15_4_lut_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_LC_10_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_LC_10_19_2  (
            .in0(N__29248),
            .in1(N__29476),
            .in2(N__28011),
            .in3(N__30919),
            .lcout(),
            .ltout(\nx.n41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i24_4_lut_LC_10_19_3 .C_ON=1'b0;
    defparam \nx.i24_4_lut_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.i24_4_lut_LC_10_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i24_4_lut_LC_10_19_3  (
            .in0(N__36933),
            .in1(N__34920),
            .in2(N__28008),
            .in3(N__31077),
            .lcout(),
            .ltout(\nx.n50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i25_4_lut_LC_10_19_4 .C_ON=1'b0;
    defparam \nx.i25_4_lut_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.i25_4_lut_LC_10_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i25_4_lut_LC_10_19_4  (
            .in0(N__28005),
            .in1(N__31383),
            .in2(N__27999),
            .in3(N__29514),
            .lcout(\nx.n3017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2034_3_lut_LC_10_19_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2034_3_lut_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2034_3_lut_LC_10_19_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i2034_3_lut_LC_10_19_5  (
            .in0(N__35118),
            .in1(_gnd_net_),
            .in2(N__35150),
            .in3(N__37307),
            .lcout(\nx.n3007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1968_3_lut_LC_10_19_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1968_3_lut_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1968_3_lut_LC_10_19_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1968_3_lut_LC_10_19_7  (
            .in0(N__27996),
            .in1(N__28215),
            .in2(_gnd_net_),
            .in3(N__37513),
            .lcout(\nx.n2909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1948_3_lut_LC_10_20_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1948_3_lut_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1948_3_lut_LC_10_20_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1948_3_lut_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__27987),
            .in2(N__37566),
            .in3(N__27975),
            .lcout(\nx.n2889 ),
            .ltout(\nx.n2889_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_3_lut_adj_112_LC_10_20_1 .C_ON=1'b0;
    defparam \nx.i5_3_lut_adj_112_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.i5_3_lut_adj_112_LC_10_20_1 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i5_3_lut_adj_112_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__35257),
            .in2(N__27942),
            .in3(N__35185),
            .lcout(\nx.n30_adj_759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1959_3_lut_LC_10_20_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1959_3_lut_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1959_3_lut_LC_10_20_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1959_3_lut_LC_10_20_2  (
            .in0(N__28110),
            .in1(_gnd_net_),
            .in2(N__37565),
            .in3(N__27939),
            .lcout(\nx.n2900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_61_LC_10_20_3 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_61_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_61_LC_10_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_61_LC_10_20_3  (
            .in0(N__28027),
            .in1(N__33845),
            .in2(N__34883),
            .in3(N__28109),
            .lcout(),
            .ltout(\nx.n40_adj_705_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_LC_10_20_4 .C_ON=1'b0;
    defparam \nx.i20_4_lut_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_LC_10_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i20_4_lut_LC_10_20_4  (
            .in0(N__37658),
            .in1(N__28081),
            .in2(N__28062),
            .in3(N__28167),
            .lcout(),
            .ltout(\nx.n44_adj_721_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i23_4_lut_adj_90_LC_10_20_5 .C_ON=1'b0;
    defparam \nx.i23_4_lut_adj_90_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.i23_4_lut_adj_90_LC_10_20_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i23_4_lut_adj_90_LC_10_20_5  (
            .in0(N__29484),
            .in1(N__28038),
            .in2(N__28059),
            .in3(N__28302),
            .lcout(\nx.n2819 ),
            .ltout(\nx.n2819_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1953_3_lut_LC_10_20_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1953_3_lut_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1953_3_lut_LC_10_20_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1953_3_lut_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__28056),
            .in2(N__28047),
            .in3(N__28137),
            .lcout(\nx.n2894 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1965_3_lut_LC_10_20_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1965_3_lut_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1965_3_lut_LC_10_20_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1965_3_lut_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(N__28044),
            .in2(N__28032),
            .in3(N__37521),
            .lcout(\nx.n2906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_74_LC_10_21_0 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_74_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_74_LC_10_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_74_LC_10_21_0  (
            .in0(N__28160),
            .in1(N__34804),
            .in2(N__29775),
            .in3(N__34168),
            .lcout(\nx.n42_adj_730 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1894_3_lut_LC_10_21_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1894_3_lut_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1894_3_lut_LC_10_21_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1894_3_lut_LC_10_21_1  (
            .in0(N__28407),
            .in1(_gnd_net_),
            .in2(N__31253),
            .in3(N__37817),
            .lcout(\nx.n2803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_3_lut_adj_114_LC_10_21_2 .C_ON=1'b0;
    defparam \nx.i13_3_lut_adj_114_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i13_3_lut_adj_114_LC_10_21_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \nx.i13_3_lut_adj_114_LC_10_21_2  (
            .in0(N__35528),
            .in1(_gnd_net_),
            .in2(N__35065),
            .in3(N__35861),
            .lcout(\nx.n38_adj_762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1898_3_lut_LC_10_21_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1898_3_lut_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1898_3_lut_LC_10_21_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1898_3_lut_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__28263),
            .in2(N__31252),
            .in3(N__35805),
            .lcout(\nx.n2807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1900_3_lut_LC_10_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1900_3_lut_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1900_3_lut_LC_10_21_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1900_3_lut_LC_10_21_4  (
            .in0(N__28293),
            .in1(N__30147),
            .in2(_gnd_net_),
            .in3(N__31205),
            .lcout(\nx.n2809 ),
            .ltout(\nx.n2809_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_3_lut_LC_10_21_5 .C_ON=1'b0;
    defparam \nx.i6_3_lut_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.i6_3_lut_LC_10_21_5 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \nx.i6_3_lut_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__28129),
            .in2(N__28218),
            .in3(N__28214),
            .lcout(\nx.n30_adj_704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1893_3_lut_LC_10_21_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1893_3_lut_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1893_3_lut_LC_10_21_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1893_3_lut_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__35771),
            .in2(N__28395),
            .in3(N__31212),
            .lcout(\nx.n2802 ),
            .ltout(\nx.n2802_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1960_3_lut_LC_10_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1960_3_lut_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1960_3_lut_LC_10_21_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1960_3_lut_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__28146),
            .in2(N__28140),
            .in3(N__37555),
            .lcout(\nx.n2901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1886_3_lut_LC_10_22_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1886_3_lut_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1886_3_lut_LC_10_22_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1886_3_lut_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__30035),
            .in2(N__31255),
            .in3(N__28500),
            .lcout(\nx.n2795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9135_3_lut_LC_10_22_1 .C_ON=1'b0;
    defparam \nx.i9135_3_lut_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.i9135_3_lut_LC_10_22_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.i9135_3_lut_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__28371),
            .in2(N__29898),
            .in3(N__31216),
            .lcout(\nx.n2800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1895_3_lut_LC_10_22_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1895_3_lut_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1895_3_lut_LC_10_22_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1895_3_lut_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__28239),
            .in2(N__31254),
            .in3(N__37856),
            .lcout(\nx.n2804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i22_4_lut_LC_10_22_3 .C_ON=1'b0;
    defparam \nx.i22_4_lut_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.i22_4_lut_LC_10_22_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i22_4_lut_LC_10_22_3  (
            .in0(N__29961),
            .in1(N__29832),
            .in2(N__29874),
            .in3(N__35745),
            .lcout(\nx.n2720 ),
            .ltout(\nx.n2720_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9137_3_lut_LC_10_22_4 .C_ON=1'b0;
    defparam \nx.i9137_3_lut_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.i9137_3_lut_LC_10_22_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.i9137_3_lut_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__28248),
            .in2(N__28113),
            .in3(N__29741),
            .lcout(\nx.n2805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1879_3_lut_LC_10_22_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1879_3_lut_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1879_3_lut_LC_10_22_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1879_3_lut_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__31220),
            .in2(N__31479),
            .in3(N__28425),
            .lcout(\nx.n2788 ),
            .ltout(\nx.n2788_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i2_2_lut_LC_10_22_6 .C_ON=1'b0;
    defparam \nx.i2_2_lut_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.i2_2_lut_LC_10_22_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i2_2_lut_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28347),
            .in3(N__28336),
            .lcout(),
            .ltout(\nx.n26_adj_706_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_78_LC_10_22_7 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_78_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_78_LC_10_22_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_78_LC_10_22_7  (
            .in0(N__28607),
            .in1(N__29938),
            .in2(N__28314),
            .in3(N__28311),
            .lcout(\nx.n43_adj_735 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_2_lut_LC_10_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_2_lut_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_2_lut_LC_10_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_2_lut_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__30142),
            .in2(_gnd_net_),
            .in3(N__28281),
            .lcout(\nx.n2777 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\nx.n10981 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_3_lut_LC_10_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_3_lut_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_3_lut_LC_10_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_3_lut_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29999),
            .in3(N__28266),
            .lcout(\nx.n2776 ),
            .ltout(),
            .carryin(\nx.n10981 ),
            .carryout(\nx.n10982 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_4_lut_LC_10_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_4_lut_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_4_lut_LC_10_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_4_lut_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__41748),
            .in2(N__35803),
            .in3(N__28254),
            .lcout(\nx.n2775 ),
            .ltout(),
            .carryin(\nx.n10982 ),
            .carryout(\nx.n10983 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_5_lut_LC_10_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_5_lut_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_5_lut_LC_10_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_5_lut_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(N__41751),
            .in2(N__31818),
            .in3(N__28251),
            .lcout(\nx.n2774 ),
            .ltout(),
            .carryin(\nx.n10983 ),
            .carryout(\nx.n10984 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_6_lut_LC_10_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_6_lut_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_6_lut_LC_10_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_6_lut_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__41749),
            .in2(N__29742),
            .in3(N__28242),
            .lcout(\nx.n2773 ),
            .ltout(),
            .carryin(\nx.n10984 ),
            .carryout(\nx.n10985 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_7_lut_LC_10_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_7_lut_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_7_lut_LC_10_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_7_lut_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(N__41752),
            .in2(N__37857),
            .in3(N__28410),
            .lcout(\nx.n2772 ),
            .ltout(),
            .carryin(\nx.n10985 ),
            .carryout(\nx.n10986 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_8_lut_LC_10_23_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_8_lut_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_8_lut_LC_10_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_8_lut_LC_10_23_6  (
            .in0(_gnd_net_),
            .in1(N__41750),
            .in2(N__37821),
            .in3(N__28398),
            .lcout(\nx.n2771 ),
            .ltout(),
            .carryin(\nx.n10986 ),
            .carryout(\nx.n10987 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_9_lut_LC_10_23_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_9_lut_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_9_lut_LC_10_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_9_lut_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(N__41753),
            .in2(N__35775),
            .in3(N__28383),
            .lcout(\nx.n2770 ),
            .ltout(),
            .carryin(\nx.n10987 ),
            .carryout(\nx.n10988 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_10_lut_LC_10_24_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_10_lut_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_10_lut_LC_10_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_10_lut_LC_10_24_0  (
            .in0(_gnd_net_),
            .in1(N__42047),
            .in2(N__34208),
            .in3(N__28374),
            .lcout(\nx.n2769 ),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\nx.n10989 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_11_lut_LC_10_24_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_11_lut_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_11_lut_LC_10_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_11_lut_LC_10_24_1  (
            .in0(_gnd_net_),
            .in1(N__42051),
            .in2(N__29894),
            .in3(N__28362),
            .lcout(\nx.n2768 ),
            .ltout(),
            .carryin(\nx.n10989 ),
            .carryout(\nx.n10990 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_12_lut_LC_10_24_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_12_lut_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_12_lut_LC_10_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_12_lut_LC_10_24_2  (
            .in0(_gnd_net_),
            .in1(N__42048),
            .in2(N__31536),
            .in3(N__28359),
            .lcout(\nx.n2767 ),
            .ltout(),
            .carryin(\nx.n10990 ),
            .carryout(\nx.n10991 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_13_lut_LC_10_24_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_13_lut_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_13_lut_LC_10_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_13_lut_LC_10_24_3  (
            .in0(_gnd_net_),
            .in1(N__42052),
            .in2(N__29922),
            .in3(N__28356),
            .lcout(\nx.n2766 ),
            .ltout(),
            .carryin(\nx.n10991 ),
            .carryout(\nx.n10992 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_14_lut_LC_10_24_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_14_lut_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_14_lut_LC_10_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_14_lut_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(N__42049),
            .in2(N__29858),
            .in3(N__28353),
            .lcout(\nx.n2765 ),
            .ltout(),
            .carryin(\nx.n10992 ),
            .carryout(\nx.n10993 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_15_lut_LC_10_24_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_15_lut_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_15_lut_LC_10_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_15_lut_LC_10_24_5  (
            .in0(_gnd_net_),
            .in1(N__42053),
            .in2(N__31301),
            .in3(N__28350),
            .lcout(\nx.n2764 ),
            .ltout(),
            .carryin(\nx.n10993 ),
            .carryout(\nx.n10994 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_16_lut_LC_10_24_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_16_lut_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_16_lut_LC_10_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_16_lut_LC_10_24_6  (
            .in0(_gnd_net_),
            .in1(N__42050),
            .in2(N__30036),
            .in3(N__28491),
            .lcout(\nx.n2763 ),
            .ltout(),
            .carryin(\nx.n10994 ),
            .carryout(\nx.n10995 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_17_lut_LC_10_24_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_17_lut_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_17_lut_LC_10_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_17_lut_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(N__42054),
            .in2(N__31668),
            .in3(N__28479),
            .lcout(\nx.n2762 ),
            .ltout(),
            .carryin(\nx.n10995 ),
            .carryout(\nx.n10996 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_18_lut_LC_10_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_18_lut_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_18_lut_LC_10_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_18_lut_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__42055),
            .in2(N__30062),
            .in3(N__28470),
            .lcout(\nx.n2761 ),
            .ltout(),
            .carryin(bfn_10_25_0_),
            .carryout(\nx.n10997 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_19_lut_LC_10_25_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_19_lut_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_19_lut_LC_10_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_19_lut_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(N__41966),
            .in2(N__30083),
            .in3(N__28461),
            .lcout(\nx.n2760 ),
            .ltout(),
            .carryin(\nx.n10997 ),
            .carryout(\nx.n10998 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_20_lut_LC_10_25_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_20_lut_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_20_lut_LC_10_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_20_lut_LC_10_25_2  (
            .in0(_gnd_net_),
            .in1(N__42056),
            .in2(N__31575),
            .in3(N__28446),
            .lcout(\nx.n2759 ),
            .ltout(),
            .carryin(\nx.n10998 ),
            .carryout(\nx.n10999 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_21_lut_LC_10_25_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_21_lut_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_21_lut_LC_10_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_21_lut_LC_10_25_3  (
            .in0(_gnd_net_),
            .in1(N__41967),
            .in2(N__31638),
            .in3(N__28437),
            .lcout(\nx.n2758 ),
            .ltout(),
            .carryin(\nx.n10999 ),
            .carryout(\nx.n11000 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_22_lut_LC_10_25_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_22_lut_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_22_lut_LC_10_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_22_lut_LC_10_25_4  (
            .in0(_gnd_net_),
            .in1(N__42057),
            .in2(N__31607),
            .in3(N__28428),
            .lcout(\nx.n2757 ),
            .ltout(),
            .carryin(\nx.n11000 ),
            .carryout(\nx.n11001 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_23_lut_LC_10_25_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_23_lut_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_23_lut_LC_10_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_23_lut_LC_10_25_5  (
            .in0(_gnd_net_),
            .in1(N__41968),
            .in2(N__31478),
            .in3(N__28416),
            .lcout(\nx.n2756 ),
            .ltout(),
            .carryin(\nx.n11001 ),
            .carryout(\nx.n11002 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_24_lut_LC_10_25_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1875_24_lut_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_24_lut_LC_10_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1875_24_lut_LC_10_25_6  (
            .in0(_gnd_net_),
            .in1(N__42058),
            .in2(N__31509),
            .in3(N__28413),
            .lcout(\nx.n2755 ),
            .ltout(),
            .carryin(\nx.n11002 ),
            .carryout(\nx.n11003 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1875_25_lut_LC_10_25_7 .C_ON=1'b0;
    defparam \nx.mod_5_add_1875_25_lut_LC_10_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1875_25_lut_LC_10_25_7 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1875_25_lut_LC_10_25_7  (
            .in0(N__42059),
            .in1(N__39983),
            .in2(N__31275),
            .in3(N__28611),
            .lcout(\nx.n2786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1417_3_lut_LC_10_26_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1417_3_lut_LC_10_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1417_3_lut_LC_10_26_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1417_3_lut_LC_10_26_0  (
            .in0(_gnd_net_),
            .in1(N__28843),
            .in2(N__28590),
            .in3(N__29120),
            .lcout(\nx.n2102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5916_2_lut_LC_10_26_1 .C_ON=1'b0;
    defparam \nx.i5916_2_lut_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.i5916_2_lut_LC_10_26_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \nx.i5916_2_lut_LC_10_26_1  (
            .in0(_gnd_net_),
            .in1(N__28937),
            .in2(_gnd_net_),
            .in3(N__29200),
            .lcout(),
            .ltout(\nx.n9709_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_31_LC_10_26_2 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_31_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_31_LC_10_26_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_31_LC_10_26_2  (
            .in0(N__28522),
            .in1(N__28744),
            .in2(N__28581),
            .in3(N__28636),
            .lcout(),
            .ltout(\nx.n26_adj_681_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_34_LC_10_26_3 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_34_LC_10_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_34_LC_10_26_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_34_LC_10_26_3  (
            .in0(N__28797),
            .in1(N__28578),
            .in2(N__28566),
            .in3(N__28536),
            .lcout(\nx.n2027 ),
            .ltout(\nx.n2027_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1421_3_lut_LC_10_26_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1421_3_lut_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1421_3_lut_LC_10_26_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1421_3_lut_LC_10_26_4  (
            .in0(N__28868),
            .in1(_gnd_net_),
            .in2(N__28563),
            .in3(N__28560),
            .lcout(\nx.n2106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_30_LC_10_26_5 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_30_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_30_LC_10_26_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_30_LC_10_26_5  (
            .in0(N__28672),
            .in1(N__28712),
            .in2(N__28789),
            .in3(N__28553),
            .lcout(\nx.n28_adj_680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1413_3_lut_LC_10_26_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1413_3_lut_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1413_3_lut_LC_10_26_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1413_3_lut_LC_10_26_6  (
            .in0(N__28523),
            .in1(_gnd_net_),
            .in2(N__28509),
            .in3(N__29121),
            .lcout(\nx.n2098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_32_LC_10_26_7 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_32_LC_10_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_32_LC_10_26_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_32_LC_10_26_7  (
            .in0(N__29021),
            .in1(N__28867),
            .in2(N__28847),
            .in3(N__28820),
            .lcout(\nx.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1418_3_lut_LC_10_27_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1418_3_lut_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1418_3_lut_LC_10_27_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1418_3_lut_LC_10_27_0  (
            .in0(N__28791),
            .in1(_gnd_net_),
            .in2(N__29122),
            .in3(N__28764),
            .lcout(\nx.n2103 ),
            .ltout(\nx.n2103_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_2_lut_LC_10_27_1 .C_ON=1'b0;
    defparam \nx.i7_2_lut_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.i7_2_lut_LC_10_27_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i7_2_lut_LC_10_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28758),
            .in3(N__30365),
            .lcout(\nx.n24_adj_684 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1412_3_lut_LC_10_27_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1412_3_lut_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1412_3_lut_LC_10_27_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1412_3_lut_LC_10_27_2  (
            .in0(_gnd_net_),
            .in1(N__28754),
            .in2(N__29124),
            .in3(N__28728),
            .lcout(\nx.n2097 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1420_3_lut_LC_10_27_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1420_3_lut_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1420_3_lut_LC_10_27_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1420_3_lut_LC_10_27_3  (
            .in0(_gnd_net_),
            .in1(N__28722),
            .in2(N__28716),
            .in3(N__29094),
            .lcout(\nx.n2105 ),
            .ltout(\nx.n2105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1487_3_lut_LC_10_27_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1487_3_lut_LC_10_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1487_3_lut_LC_10_27_4 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.mod_5_i1487_3_lut_LC_10_27_4  (
            .in0(N__36533),
            .in1(N__30354),
            .in2(N__28683),
            .in3(_gnd_net_),
            .lcout(\nx.n2204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1419_3_lut_LC_10_27_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1419_3_lut_LC_10_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1419_3_lut_LC_10_27_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1419_3_lut_LC_10_27_5  (
            .in0(_gnd_net_),
            .in1(N__28680),
            .in2(N__28653),
            .in3(N__29095),
            .lcout(\nx.n2104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1416_3_lut_LC_10_27_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1416_3_lut_LC_10_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1416_3_lut_LC_10_27_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1416_3_lut_LC_10_27_6  (
            .in0(_gnd_net_),
            .in1(N__28643),
            .in2(N__29123),
            .in3(N__28617),
            .lcout(\nx.n2101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1492_3_lut_LC_10_27_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1492_3_lut_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1492_3_lut_LC_10_27_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1492_3_lut_LC_10_27_7  (
            .in0(_gnd_net_),
            .in1(N__30528),
            .in2(N__30486),
            .in3(N__36532),
            .lcout(\nx.n2209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1422_3_lut_LC_10_28_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1422_3_lut_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1422_3_lut_LC_10_28_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1422_3_lut_LC_10_28_0  (
            .in0(_gnd_net_),
            .in1(N__29034),
            .in2(N__29025),
            .in3(N__29106),
            .lcout(\nx.n2107 ),
            .ltout(\nx.n2107_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_39_LC_10_28_1 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_39_LC_10_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_39_LC_10_28_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \nx.i12_4_lut_adj_39_LC_10_28_1  (
            .in0(N__30470),
            .in1(N__30533),
            .in2(N__28992),
            .in3(N__28989),
            .lcout(\nx.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1411_3_lut_LC_10_28_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1411_3_lut_LC_10_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1411_3_lut_LC_10_28_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1411_3_lut_LC_10_28_2  (
            .in0(_gnd_net_),
            .in1(N__28983),
            .in2(N__28953),
            .in3(N__29107),
            .lcout(\nx.n2096 ),
            .ltout(\nx.n2096_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_45_LC_10_28_3 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_45_LC_10_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_45_LC_10_28_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_45_LC_10_28_3  (
            .in0(N__30671),
            .in1(N__30628),
            .in2(N__28944),
            .in3(N__30562),
            .lcout(\nx.n27_adj_691 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1424_3_lut_LC_10_28_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1424_3_lut_LC_10_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1424_3_lut_LC_10_28_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i1424_3_lut_LC_10_28_4  (
            .in0(N__28941),
            .in1(N__28893),
            .in2(_gnd_net_),
            .in3(N__29105),
            .lcout(\nx.n2109 ),
            .ltout(\nx.n2109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1491_3_lut_LC_10_28_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1491_3_lut_LC_10_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1491_3_lut_LC_10_28_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1491_3_lut_LC_10_28_5  (
            .in0(N__30456),
            .in1(_gnd_net_),
            .in2(N__28881),
            .in3(N__36534),
            .lcout(\nx.n2208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1485_3_lut_LC_10_28_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1485_3_lut_LC_10_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1485_3_lut_LC_10_28_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1485_3_lut_LC_10_28_6  (
            .in0(_gnd_net_),
            .in1(N__30291),
            .in2(N__36559),
            .in3(N__30305),
            .lcout(\nx.n2202 ),
            .ltout(\nx.n2202_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i4_3_lut_LC_10_28_7 .C_ON=1'b0;
    defparam \nx.i4_3_lut_LC_10_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.i4_3_lut_LC_10_28_7 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \nx.i4_3_lut_LC_10_28_7  (
            .in0(N__31696),
            .in1(_gnd_net_),
            .in2(N__28878),
            .in3(N__31789),
            .lcout(\nx.n22_adj_693 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_37_LC_10_29_0 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_37_LC_10_29_0 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_37_LC_10_29_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_37_LC_10_29_0  (
            .in0(N__30446),
            .in1(N__30398),
            .in2(N__32707),
            .in3(N__28875),
            .lcout(\nx.n30_adj_685 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1478_3_lut_LC_10_29_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1478_3_lut_LC_10_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1478_3_lut_LC_10_29_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1478_3_lut_LC_10_29_1  (
            .in0(N__30596),
            .in1(_gnd_net_),
            .in2(N__30582),
            .in3(N__36525),
            .lcout(\nx.n2195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1476_3_lut_LC_10_29_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1476_3_lut_LC_10_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1476_3_lut_LC_10_29_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1476_3_lut_LC_10_29_2  (
            .in0(_gnd_net_),
            .in1(N__30887),
            .in2(N__36558),
            .in3(N__30873),
            .lcout(\nx.n2193 ),
            .ltout(\nx.n2193_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i10_4_lut_adj_47_LC_10_29_3 .C_ON=1'b0;
    defparam \nx.i10_4_lut_adj_47_LC_10_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.i10_4_lut_adj_47_LC_10_29_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i10_4_lut_adj_47_LC_10_29_3  (
            .in0(N__32596),
            .in1(N__32638),
            .in2(N__29208),
            .in3(N__30833),
            .lcout(\nx.n28_adj_692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1423_3_lut_LC_10_29_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1423_3_lut_LC_10_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1423_3_lut_LC_10_29_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1423_3_lut_LC_10_29_4  (
            .in0(_gnd_net_),
            .in1(N__29205),
            .in2(N__29175),
            .in3(N__29116),
            .lcout(\nx.n2108 ),
            .ltout(\nx.n2108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1490_3_lut_LC_10_29_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1490_3_lut_LC_10_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1490_3_lut_LC_10_29_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1490_3_lut_LC_10_29_5  (
            .in0(_gnd_net_),
            .in1(N__30432),
            .in2(N__29160),
            .in3(N__36524),
            .lcout(\nx.n2207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1488_3_lut_LC_10_29_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1488_3_lut_LC_10_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1488_3_lut_LC_10_29_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1488_3_lut_LC_10_29_6  (
            .in0(N__30381),
            .in1(_gnd_net_),
            .in2(N__36557),
            .in3(N__30399),
            .lcout(\nx.n2205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1410_3_lut_LC_10_29_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1410_3_lut_LC_10_29_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1410_3_lut_LC_10_29_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1410_3_lut_LC_10_29_7  (
            .in0(_gnd_net_),
            .in1(N__29153),
            .in2(N__29127),
            .in3(N__29043),
            .lcout(\nx.n2095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_15_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_15_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_15_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_82_LC_11_17_0 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_82_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_82_LC_11_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_82_LC_11_17_0  (
            .in0(N__33508),
            .in1(N__33412),
            .in2(N__33466),
            .in3(N__34126),
            .lcout(),
            .ltout(\nx.n42_adj_739_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i21_4_lut_adj_85_LC_11_17_1 .C_ON=1'b0;
    defparam \nx.i21_4_lut_adj_85_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.i21_4_lut_adj_85_LC_11_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i21_4_lut_adj_85_LC_11_17_1  (
            .in0(N__33328),
            .in1(N__34078),
            .in2(N__29397),
            .in3(N__33887),
            .lcout(\nx.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_2_lut_adj_83_LC_11_17_2 .C_ON=1'b0;
    defparam \nx.i5_2_lut_adj_83_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \nx.i5_2_lut_adj_83_LC_11_17_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \nx.i5_2_lut_adj_83_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__33685),
            .in2(_gnd_net_),
            .in3(N__33640),
            .lcout(),
            .ltout(\nx.n32_adj_740_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i22_4_lut_adj_86_LC_11_17_3 .C_ON=1'b0;
    defparam \nx.i22_4_lut_adj_86_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.i22_4_lut_adj_86_LC_11_17_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i22_4_lut_adj_86_LC_11_17_3  (
            .in0(N__33595),
            .in1(N__33553),
            .in2(N__29394),
            .in3(N__29391),
            .lcout(),
            .ltout(\nx.n49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i26_4_lut_LC_11_17_4 .C_ON=1'b0;
    defparam \nx.i26_4_lut_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \nx.i26_4_lut_LC_11_17_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i26_4_lut_LC_11_17_4  (
            .in0(N__29379),
            .in1(N__29373),
            .in2(N__29358),
            .in3(N__29355),
            .lcout(\nx.n3116 ),
            .ltout(\nx.n3116_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2167_3_lut_LC_11_17_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2167_3_lut_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2167_3_lut_LC_11_17_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2167_3_lut_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__32924),
            .in2(N__29349),
            .in3(N__32904),
            .lcout(\nx.n19_adj_745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_2_lut_LC_11_18_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_2_lut_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_2_lut_LC_11_18_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_2076_2_lut_LC_11_18_0  (
            .in0(N__29346),
            .in1(N__29345),
            .in2(N__29276),
            .in3(N__29301),
            .lcout(\nx.n3109 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\nx.n11053 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_3_lut_LC_11_18_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_3_lut_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_3_lut_LC_11_18_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \nx.mod_5_add_2076_3_lut_LC_11_18_1  (
            .in0(N__29298),
            .in1(N__29297),
            .in2(N__29277),
            .in3(N__29253),
            .lcout(\nx.n3108 ),
            .ltout(),
            .carryin(\nx.n11053 ),
            .carryout(\nx.n11054 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_4_lut_LC_11_18_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_4_lut_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_4_lut_LC_11_18_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_4_lut_LC_11_18_2  (
            .in0(N__29250),
            .in1(N__29249),
            .in2(N__29670),
            .in3(N__29232),
            .lcout(\nx.n3107 ),
            .ltout(),
            .carryin(\nx.n11054 ),
            .carryout(\nx.n11055 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_5_lut_LC_11_18_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_5_lut_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_5_lut_LC_11_18_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_5_lut_LC_11_18_3  (
            .in0(N__29229),
            .in1(N__29228),
            .in2(N__29673),
            .in3(N__29211),
            .lcout(\nx.n3106 ),
            .ltout(),
            .carryin(\nx.n11055 ),
            .carryout(\nx.n11056 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_6_lut_LC_11_18_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_6_lut_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_6_lut_LC_11_18_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_6_lut_LC_11_18_4  (
            .in0(N__34959),
            .in1(N__34958),
            .in2(N__29671),
            .in3(N__29424),
            .lcout(\nx.n3105 ),
            .ltout(),
            .carryin(\nx.n11056 ),
            .carryout(\nx.n11057 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_7_lut_LC_11_18_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_7_lut_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_7_lut_LC_11_18_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_7_lut_LC_11_18_5  (
            .in0(N__31050),
            .in1(N__31049),
            .in2(N__29674),
            .in3(N__29421),
            .lcout(\nx.n3104 ),
            .ltout(),
            .carryin(\nx.n11057 ),
            .carryout(\nx.n11058 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_8_lut_LC_11_18_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_8_lut_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_8_lut_LC_11_18_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_8_lut_LC_11_18_6  (
            .in0(N__34944),
            .in1(N__34943),
            .in2(N__29672),
            .in3(N__29418),
            .lcout(\nx.n3103 ),
            .ltout(),
            .carryin(\nx.n11058 ),
            .carryout(\nx.n11059 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_9_lut_LC_11_18_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_9_lut_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_9_lut_LC_11_18_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_9_lut_LC_11_18_7  (
            .in0(N__31068),
            .in1(N__31067),
            .in2(N__29675),
            .in3(N__29415),
            .lcout(\nx.n3102 ),
            .ltout(),
            .carryin(\nx.n11059 ),
            .carryout(\nx.n11060 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_10_lut_LC_11_19_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_10_lut_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_10_lut_LC_11_19_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_10_lut_LC_11_19_0  (
            .in0(N__36978),
            .in1(N__36977),
            .in2(N__29676),
            .in3(N__29412),
            .lcout(\nx.n3101 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\nx.n11061 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_11_lut_LC_11_19_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_11_lut_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_11_lut_LC_11_19_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_11_lut_LC_11_19_1  (
            .in0(N__31092),
            .in1(N__31091),
            .in2(N__29680),
            .in3(N__29409),
            .lcout(\nx.n3100 ),
            .ltout(),
            .carryin(\nx.n11061 ),
            .carryout(\nx.n11062 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_12_lut_LC_11_19_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_12_lut_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_12_lut_LC_11_19_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_12_lut_LC_11_19_2  (
            .in0(N__31112),
            .in1(N__31111),
            .in2(N__29677),
            .in3(N__29406),
            .lcout(\nx.n3099 ),
            .ltout(),
            .carryin(\nx.n11062 ),
            .carryout(\nx.n11063 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_13_lut_LC_11_19_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_13_lut_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_13_lut_LC_11_19_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_13_lut_LC_11_19_3  (
            .in0(N__34908),
            .in1(N__34907),
            .in2(N__29681),
            .in3(N__29403),
            .lcout(\nx.n3098 ),
            .ltout(),
            .carryin(\nx.n11063 ),
            .carryout(\nx.n11064 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_14_lut_LC_11_19_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_14_lut_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_14_lut_LC_11_19_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_14_lut_LC_11_19_4  (
            .in0(N__29478),
            .in1(N__29477),
            .in2(N__29678),
            .in3(N__29400),
            .lcout(\nx.n3097 ),
            .ltout(),
            .carryin(\nx.n11064 ),
            .carryout(\nx.n11065 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_15_lut_LC_11_19_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_15_lut_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_15_lut_LC_11_19_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_15_lut_LC_11_19_5  (
            .in0(N__31398),
            .in1(N__31397),
            .in2(N__29682),
            .in3(N__29451),
            .lcout(\nx.n3096 ),
            .ltout(),
            .carryin(\nx.n11065 ),
            .carryout(\nx.n11066 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_16_lut_LC_11_19_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_16_lut_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_16_lut_LC_11_19_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_16_lut_LC_11_19_6  (
            .in0(N__29505),
            .in1(N__29504),
            .in2(N__29679),
            .in3(N__29448),
            .lcout(\nx.n3095 ),
            .ltout(),
            .carryin(\nx.n11066 ),
            .carryout(\nx.n11067 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_17_lut_LC_11_19_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_17_lut_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_17_lut_LC_11_19_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_17_lut_LC_11_19_7  (
            .in0(N__36960),
            .in1(N__36959),
            .in2(N__29683),
            .in3(N__29445),
            .lcout(\nx.n3094 ),
            .ltout(),
            .carryin(\nx.n11067 ),
            .carryout(\nx.n11068 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_18_lut_LC_11_20_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_18_lut_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_18_lut_LC_11_20_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_18_lut_LC_11_20_0  (
            .in0(N__31013),
            .in1(N__31012),
            .in2(N__29684),
            .in3(N__29442),
            .lcout(\nx.n3093 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\nx.n11069 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_19_lut_LC_11_20_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_19_lut_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_19_lut_LC_11_20_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_19_lut_LC_11_20_1  (
            .in0(N__37167),
            .in1(N__37166),
            .in2(N__29688),
            .in3(N__29439),
            .lcout(\nx.n3092 ),
            .ltout(),
            .carryin(\nx.n11069 ),
            .carryout(\nx.n11070 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_20_lut_LC_11_20_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_20_lut_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_20_lut_LC_11_20_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_20_lut_LC_11_20_2  (
            .in0(N__37686),
            .in1(N__37685),
            .in2(N__29685),
            .in3(N__29436),
            .lcout(\nx.n3091 ),
            .ltout(),
            .carryin(\nx.n11070 ),
            .carryout(\nx.n11071 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_21_lut_LC_11_20_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_21_lut_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_21_lut_LC_11_20_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_21_lut_LC_11_20_3  (
            .in0(N__33732),
            .in1(N__33731),
            .in2(N__29689),
            .in3(N__29433),
            .lcout(\nx.n3090 ),
            .ltout(),
            .carryin(\nx.n11071 ),
            .carryout(\nx.n11072 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_22_lut_LC_11_20_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_22_lut_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_22_lut_LC_11_20_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_22_lut_LC_11_20_4  (
            .in0(N__36873),
            .in1(N__36872),
            .in2(N__29686),
            .in3(N__29430),
            .lcout(\nx.n3089 ),
            .ltout(),
            .carryin(\nx.n11072 ),
            .carryout(\nx.n11073 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_23_lut_LC_11_20_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_23_lut_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_23_lut_LC_11_20_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_23_lut_LC_11_20_5  (
            .in0(N__30924),
            .in1(N__30920),
            .in2(N__29690),
            .in3(N__29427),
            .lcout(\nx.n3088 ),
            .ltout(),
            .carryin(\nx.n11073 ),
            .carryout(\nx.n11074 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_24_lut_LC_11_20_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_24_lut_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_24_lut_LC_11_20_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_24_lut_LC_11_20_6  (
            .in0(N__31371),
            .in1(N__31370),
            .in2(N__29687),
            .in3(N__29727),
            .lcout(\nx.n3087 ),
            .ltout(),
            .carryin(\nx.n11074 ),
            .carryout(\nx.n11075 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_25_lut_LC_11_20_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_25_lut_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_25_lut_LC_11_20_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_25_lut_LC_11_20_7  (
            .in0(N__29724),
            .in1(N__29723),
            .in2(N__29691),
            .in3(N__29712),
            .lcout(\nx.n3086 ),
            .ltout(),
            .carryin(\nx.n11075 ),
            .carryout(\nx.n11076 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_26_lut_LC_11_21_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_26_lut_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_26_lut_LC_11_21_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_26_lut_LC_11_21_0  (
            .in0(N__33753),
            .in1(N__33752),
            .in2(N__29701),
            .in3(N__29709),
            .lcout(\nx.n3085 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\nx.n11077 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_27_lut_LC_11_21_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2076_27_lut_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_27_lut_LC_11_21_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_27_lut_LC_11_21_1  (
            .in0(N__29799),
            .in1(N__29798),
            .in2(N__29703),
            .in3(N__29706),
            .lcout(\nx.n3084 ),
            .ltout(),
            .carryin(\nx.n11077 ),
            .carryout(\nx.n11078 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2076_28_lut_LC_11_21_2 .C_ON=1'b0;
    defparam \nx.mod_5_add_2076_28_lut_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2076_28_lut_LC_11_21_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \nx.mod_5_add_2076_28_lut_LC_11_21_2  (
            .in0(N__35844),
            .in1(N__35843),
            .in2(N__29702),
            .in3(N__29517),
            .lcout(\nx.n3083 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_LC_11_21_3 .C_ON=1'b0;
    defparam \nx.i14_4_lut_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_LC_11_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_LC_11_21_3  (
            .in0(N__29497),
            .in1(N__31113),
            .in2(N__31014),
            .in3(N__29797),
            .lcout(\nx.n40_adj_670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2023_3_lut_LC_11_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2023_3_lut_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2023_3_lut_LC_11_21_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2023_3_lut_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__35307),
            .in2(N__37392),
            .in3(N__37313),
            .lcout(\nx.n2996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_79_LC_11_21_5 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_79_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_79_LC_11_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_79_LC_11_21_5  (
            .in0(N__31432),
            .in1(N__36841),
            .in2(N__31139),
            .in3(N__33796),
            .lcout(\nx.n41_adj_736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2025_3_lut_LC_11_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_i2025_3_lut_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2025_3_lut_LC_11_21_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2025_3_lut_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__35334),
            .in2(N__37323),
            .in3(N__35356),
            .lcout(\nx.n2998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1888_3_lut_LC_11_22_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1888_3_lut_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1888_3_lut_LC_11_22_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1888_3_lut_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__29841),
            .in2(N__29862),
            .in3(N__31230),
            .lcout(\nx.n2797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_41_LC_11_22_1 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_41_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_41_LC_11_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_41_LC_11_22_1  (
            .in0(N__31495),
            .in1(N__34201),
            .in2(N__39984),
            .in3(N__31542),
            .lcout(\nx.n41_adj_688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1890_3_lut_LC_11_22_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1890_3_lut_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1890_3_lut_LC_11_22_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \nx.mod_5_i1890_3_lut_LC_11_22_3  (
            .in0(N__29826),
            .in1(N__31529),
            .in2(N__31259),
            .in3(_gnd_net_),
            .lcout(\nx.n2799 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1945_3_lut_LC_11_22_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1945_3_lut_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1945_3_lut_LC_11_22_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1945_3_lut_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__29942),
            .in2(N__29817),
            .in3(N__37575),
            .lcout(\nx.n2886 ),
            .ltout(\nx.n2886_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2012_3_lut_LC_11_22_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2012_3_lut_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2012_3_lut_LC_11_22_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i2012_3_lut_LC_11_22_5  (
            .in0(N__37317),
            .in1(_gnd_net_),
            .in2(N__29802),
            .in3(N__35883),
            .lcout(\nx.n2985 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1897_3_lut_LC_11_22_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1897_3_lut_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1897_3_lut_LC_11_22_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1897_3_lut_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__31814),
            .in2(N__29784),
            .in3(N__31226),
            .lcout(\nx.n2806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1958_3_lut_LC_11_22_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1958_3_lut_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1958_3_lut_LC_11_22_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1958_3_lut_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__29773),
            .in2(N__37602),
            .in3(N__29751),
            .lcout(\nx.n2899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1813_3_lut_LC_11_23_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1813_3_lut_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1813_3_lut_LC_11_23_0 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.mod_5_i1813_3_lut_LC_11_23_0  (
            .in0(N__40098),
            .in1(N__39384),
            .in2(N__39410),
            .in3(_gnd_net_),
            .lcout(\nx.n2690 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1829_3_lut_LC_11_23_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1829_3_lut_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1829_3_lut_LC_11_23_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1829_3_lut_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__38784),
            .in2(N__38757),
            .in3(N__40097),
            .lcout(\nx.n2706 ),
            .ltout(\nx.n2706_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_40_LC_11_23_2 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_40_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_40_LC_11_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_40_LC_11_23_2  (
            .in0(N__29921),
            .in1(N__31813),
            .in2(N__29964),
            .in3(N__31528),
            .lcout(\nx.n40_adj_687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1819_3_lut_LC_11_23_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1819_3_lut_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1819_3_lut_LC_11_23_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1819_3_lut_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(N__39683),
            .in2(N__39669),
            .in3(N__40096),
            .lcout(\nx.n2696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1820_3_lut_LC_11_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1820_3_lut_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1820_3_lut_LC_11_23_4 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \nx.mod_5_i1820_3_lut_LC_11_23_4  (
            .in0(N__40099),
            .in1(N__39705),
            .in2(N__39735),
            .in3(_gnd_net_),
            .lcout(\nx.n2697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1878_3_lut_LC_11_23_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1878_3_lut_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1878_3_lut_LC_11_23_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1878_3_lut_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(N__31222),
            .in2(N__31505),
            .in3(N__29955),
            .lcout(\nx.n2787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1822_3_lut_LC_11_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1822_3_lut_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1822_3_lut_LC_11_23_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \nx.mod_5_i1822_3_lut_LC_11_23_6  (
            .in0(N__40100),
            .in1(_gnd_net_),
            .in2(N__39108),
            .in3(N__39138),
            .lcout(\nx.n2699 ),
            .ltout(\nx.n2699_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1889_3_lut_LC_11_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1889_3_lut_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1889_3_lut_LC_11_23_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1889_3_lut_LC_11_23_7  (
            .in0(N__29907),
            .in1(_gnd_net_),
            .in2(N__29901),
            .in3(N__31221),
            .lcout(\nx.n2798 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9134_3_lut_LC_11_24_0 .C_ON=1'b0;
    defparam \nx.i9134_3_lut_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.i9134_3_lut_LC_11_24_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.i9134_3_lut_LC_11_24_0  (
            .in0(N__39221),
            .in1(_gnd_net_),
            .in2(N__40094),
            .in3(N__39195),
            .lcout(\nx.n2701 ),
            .ltout(\nx.n2701_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_36_LC_11_24_1 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_36_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_36_LC_11_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_36_LC_11_24_1  (
            .in0(N__30093),
            .in1(N__31294),
            .in2(N__29877),
            .in3(N__30015),
            .lcout(\nx.n42_adj_683 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1821_3_lut_LC_11_24_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1821_3_lut_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1821_3_lut_LC_11_24_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1821_3_lut_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(N__39086),
            .in2(N__40093),
            .in3(N__39057),
            .lcout(\nx.n2698 ),
            .ltout(\nx.n2698_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i7_3_lut_LC_11_24_3 .C_ON=1'b0;
    defparam \nx.i7_3_lut_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.i7_3_lut_LC_11_24_3 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \nx.i7_3_lut_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__30132),
            .in2(N__30096),
            .in3(N__29995),
            .lcout(\nx.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1817_3_lut_LC_11_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1817_3_lut_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1817_3_lut_LC_11_24_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1817_3_lut_LC_11_24_4  (
            .in0(_gnd_net_),
            .in1(N__39567),
            .in2(N__40092),
            .in3(N__39600),
            .lcout(\nx.n2694 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1816_3_lut_LC_11_24_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1816_3_lut_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1816_3_lut_LC_11_24_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1816_3_lut_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__39549),
            .in2(N__39522),
            .in3(N__40058),
            .lcout(\nx.n2693 ),
            .ltout(\nx.n2693_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_23_LC_11_24_6 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_23_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_23_LC_11_24_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_23_LC_11_24_6  (
            .in0(N__30055),
            .in1(N__31657),
            .in2(N__30039),
            .in3(N__30031),
            .lcout(\nx.n37_adj_677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1832_3_lut_LC_11_24_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1832_3_lut_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1832_3_lut_LC_11_24_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i1832_3_lut_LC_11_24_7  (
            .in0(N__38920),
            .in1(N__38883),
            .in2(_gnd_net_),
            .in3(N__40051),
            .lcout(\nx.n2709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_2_lut_LC_11_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_2_lut_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_2_lut_LC_11_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_2_lut_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(N__31794),
            .in2(_gnd_net_),
            .in3(N__29976),
            .lcout(\nx.n2277 ),
            .ltout(),
            .carryin(bfn_11_25_0_),
            .carryout(\nx.n10881 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_3_lut_LC_11_25_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_3_lut_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_3_lut_LC_11_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_3_lut_LC_11_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31703),
            .in3(N__29973),
            .lcout(\nx.n2276 ),
            .ltout(),
            .carryin(\nx.n10881 ),
            .carryout(\nx.n10882 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_4_lut_LC_11_25_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_4_lut_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_4_lut_LC_11_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_4_lut_LC_11_25_2  (
            .in0(_gnd_net_),
            .in1(N__41559),
            .in2(N__32072),
            .in3(N__29970),
            .lcout(\nx.n2275 ),
            .ltout(),
            .carryin(\nx.n10882 ),
            .carryout(\nx.n10883 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_5_lut_LC_11_25_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_5_lut_LC_11_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_5_lut_LC_11_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_5_lut_LC_11_25_3  (
            .in0(_gnd_net_),
            .in1(N__41561),
            .in2(N__32106),
            .in3(N__29967),
            .lcout(\nx.n2274 ),
            .ltout(),
            .carryin(\nx.n10883 ),
            .carryout(\nx.n10884 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_6_lut_LC_11_25_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_6_lut_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_6_lut_LC_11_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_6_lut_LC_11_25_4  (
            .in0(_gnd_net_),
            .in1(N__31724),
            .in2(N__41963),
            .in3(N__30174),
            .lcout(\nx.n2273 ),
            .ltout(),
            .carryin(\nx.n10884 ),
            .carryout(\nx.n10885 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_7_lut_LC_11_25_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_7_lut_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_7_lut_LC_11_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_7_lut_LC_11_25_5  (
            .in0(_gnd_net_),
            .in1(N__41565),
            .in2(N__32025),
            .in3(N__30171),
            .lcout(\nx.n2272 ),
            .ltout(),
            .carryin(\nx.n10885 ),
            .carryout(\nx.n10886 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_8_lut_LC_11_25_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_8_lut_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_8_lut_LC_11_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_8_lut_LC_11_25_6  (
            .in0(_gnd_net_),
            .in1(N__41560),
            .in2(N__31955),
            .in3(N__30168),
            .lcout(\nx.n2271 ),
            .ltout(),
            .carryin(\nx.n10886 ),
            .carryout(\nx.n10887 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_9_lut_LC_11_25_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_9_lut_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_9_lut_LC_11_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_9_lut_LC_11_25_7  (
            .in0(_gnd_net_),
            .in1(N__41566),
            .in2(N__31883),
            .in3(N__30165),
            .lcout(\nx.n2270 ),
            .ltout(),
            .carryin(\nx.n10887 ),
            .carryout(\nx.n10888 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_10_lut_LC_11_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_10_lut_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_10_lut_LC_11_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_10_lut_LC_11_26_0  (
            .in0(_gnd_net_),
            .in1(N__41567),
            .in2(N__31904),
            .in3(N__30162),
            .lcout(\nx.n2269 ),
            .ltout(),
            .carryin(bfn_11_26_0_),
            .carryout(\nx.n10889 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_11_lut_LC_11_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_11_lut_LC_11_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_11_lut_LC_11_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_11_lut_LC_11_26_1  (
            .in0(_gnd_net_),
            .in1(N__41573),
            .in2(N__32673),
            .in3(N__30159),
            .lcout(\nx.n2268 ),
            .ltout(),
            .carryin(\nx.n10889 ),
            .carryout(\nx.n10890 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_12_lut_LC_11_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_12_lut_LC_11_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_12_lut_LC_11_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_12_lut_LC_11_26_2  (
            .in0(_gnd_net_),
            .in1(N__41568),
            .in2(N__36459),
            .in3(N__30156),
            .lcout(\nx.n2267 ),
            .ltout(),
            .carryin(\nx.n10890 ),
            .carryout(\nx.n10891 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_13_lut_LC_11_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_13_lut_LC_11_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_13_lut_LC_11_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_13_lut_LC_11_26_3  (
            .in0(_gnd_net_),
            .in1(N__31979),
            .in2(N__41964),
            .in3(N__30153),
            .lcout(\nx.n2266 ),
            .ltout(),
            .carryin(\nx.n10891 ),
            .carryout(\nx.n10892 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_14_lut_LC_11_26_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_14_lut_LC_11_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_14_lut_LC_11_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_14_lut_LC_11_26_4  (
            .in0(_gnd_net_),
            .in1(N__32133),
            .in2(N__41965),
            .in3(N__30150),
            .lcout(\nx.n2265 ),
            .ltout(),
            .carryin(\nx.n10892 ),
            .carryout(\nx.n10893 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_15_lut_LC_11_26_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_15_lut_LC_11_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_15_lut_LC_11_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_15_lut_LC_11_26_5  (
            .in0(_gnd_net_),
            .in1(N__41577),
            .in2(N__32297),
            .in3(N__30201),
            .lcout(\nx.n2264 ),
            .ltout(),
            .carryin(\nx.n10893 ),
            .carryout(\nx.n10894 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_16_lut_LC_11_26_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_16_lut_LC_11_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_16_lut_LC_11_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_16_lut_LC_11_26_6  (
            .in0(_gnd_net_),
            .in1(N__41572),
            .in2(N__32274),
            .in3(N__30198),
            .lcout(\nx.n2263 ),
            .ltout(),
            .carryin(\nx.n10894 ),
            .carryout(\nx.n10895 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_17_lut_LC_11_26_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_17_lut_LC_11_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_17_lut_LC_11_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_17_lut_LC_11_26_7  (
            .in0(_gnd_net_),
            .in1(N__41578),
            .in2(N__32609),
            .in3(N__30195),
            .lcout(\nx.n2262 ),
            .ltout(),
            .carryin(\nx.n10895 ),
            .carryout(\nx.n10896 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_18_lut_LC_11_27_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_18_lut_LC_11_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_18_lut_LC_11_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_18_lut_LC_11_27_0  (
            .in0(_gnd_net_),
            .in1(N__41589),
            .in2(N__32643),
            .in3(N__30192),
            .lcout(\nx.n2261 ),
            .ltout(),
            .carryin(bfn_11_27_0_),
            .carryout(\nx.n10897 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_19_lut_LC_11_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1540_19_lut_LC_11_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_19_lut_LC_11_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1540_19_lut_LC_11_27_1  (
            .in0(_gnd_net_),
            .in1(N__41590),
            .in2(N__30281),
            .in3(N__30189),
            .lcout(\nx.n2260 ),
            .ltout(),
            .carryin(\nx.n10897 ),
            .carryout(\nx.n10898 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1540_20_lut_LC_11_27_2 .C_ON=1'b0;
    defparam \nx.mod_5_add_1540_20_lut_LC_11_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1540_20_lut_LC_11_27_2 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_1540_20_lut_LC_11_27_2  (
            .in0(N__41591),
            .in1(N__32560),
            .in2(N__30840),
            .in3(N__30186),
            .lcout(\nx.n2291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1479_3_lut_LC_11_27_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1479_3_lut_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1479_3_lut_LC_11_27_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1479_3_lut_LC_11_27_3  (
            .in0(_gnd_net_),
            .in1(N__30612),
            .in2(N__30636),
            .in3(N__36538),
            .lcout(\nx.n2196 ),
            .ltout(\nx.n2196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1546_3_lut_LC_11_27_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1546_3_lut_LC_11_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1546_3_lut_LC_11_27_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1546_3_lut_LC_11_27_4  (
            .in0(_gnd_net_),
            .in1(N__30183),
            .in2(N__30177),
            .in3(N__32558),
            .lcout(\nx.n2295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_49_LC_11_27_5 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_49_LC_11_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_49_LC_11_27_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_49_LC_11_27_5  (
            .in0(N__32128),
            .in1(N__32062),
            .in2(N__31951),
            .in3(N__32665),
            .lcout(\nx.n30_adj_694 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1480_3_lut_LC_11_27_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1480_3_lut_LC_11_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1480_3_lut_LC_11_27_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1480_3_lut_LC_11_27_6  (
            .in0(N__30670),
            .in1(_gnd_net_),
            .in2(N__36560),
            .in3(N__30648),
            .lcout(\nx.n2197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1543_3_lut_LC_11_27_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1543_3_lut_LC_11_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1543_3_lut_LC_11_27_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i1543_3_lut_LC_11_27_7  (
            .in0(N__32559),
            .in1(_gnd_net_),
            .in2(N__30282),
            .in3(N__30264),
            .lcout(\nx.n2292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1477_3_lut_LC_11_28_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1477_3_lut_LC_11_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1477_3_lut_LC_11_28_0 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1477_3_lut_LC_11_28_0  (
            .in0(_gnd_net_),
            .in1(N__36548),
            .in2(N__30570),
            .in3(N__30546),
            .lcout(\nx.n2194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_46_LC_11_28_1 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_46_LC_11_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_46_LC_11_28_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_46_LC_11_28_1  (
            .in0(N__30258),
            .in1(N__30252),
            .in2(N__30243),
            .in3(N__30234),
            .lcout(\nx.n2126 ),
            .ltout(\nx.n2126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1489_3_lut_LC_11_28_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1489_3_lut_LC_11_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1489_3_lut_LC_11_28_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1489_3_lut_LC_11_28_2  (
            .in0(N__30408),
            .in1(_gnd_net_),
            .in2(N__30228),
            .in3(N__30422),
            .lcout(\nx.n2206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1482_3_lut_LC_11_28_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1482_3_lut_LC_11_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1482_3_lut_LC_11_28_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \nx.mod_5_i1482_3_lut_LC_11_28_3  (
            .in0(N__36552),
            .in1(_gnd_net_),
            .in2(N__30696),
            .in3(N__30722),
            .lcout(\nx.n2199 ),
            .ltout(\nx.n2199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_48_LC_11_28_4 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_48_LC_11_28_4 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_48_LC_11_28_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_48_LC_11_28_4  (
            .in0(N__31723),
            .in1(N__32092),
            .in2(N__30225),
            .in3(N__32011),
            .lcout(),
            .ltout(\nx.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_50_LC_11_28_5 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_50_LC_11_28_5 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_50_LC_11_28_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_50_LC_11_28_5  (
            .in0(N__36455),
            .in1(N__31873),
            .in2(N__30222),
            .in3(N__30219),
            .lcout(\nx.n34_adj_695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1486_3_lut_LC_11_28_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1486_3_lut_LC_11_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1486_3_lut_LC_11_28_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1486_3_lut_LC_11_28_7  (
            .in0(_gnd_net_),
            .in1(N__30318),
            .in2(N__36563),
            .in3(N__30338),
            .lcout(\nx.n2203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_2_lut_LC_11_29_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_2_lut_LC_11_29_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_2_lut_LC_11_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_2_lut_LC_11_29_0  (
            .in0(_gnd_net_),
            .in1(N__30532),
            .in2(_gnd_net_),
            .in3(N__30474),
            .lcout(\nx.n2177 ),
            .ltout(),
            .carryin(bfn_11_29_0_),
            .carryout(\nx.n10864 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_3_lut_LC_11_29_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_3_lut_LC_11_29_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_3_lut_LC_11_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_3_lut_LC_11_29_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30471),
            .in3(N__30450),
            .lcout(\nx.n2176 ),
            .ltout(),
            .carryin(\nx.n10864 ),
            .carryout(\nx.n10865 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_4_lut_LC_11_29_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_4_lut_LC_11_29_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_4_lut_LC_11_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_4_lut_LC_11_29_2  (
            .in0(_gnd_net_),
            .in1(N__42199),
            .in2(N__30447),
            .in3(N__30426),
            .lcout(\nx.n2175 ),
            .ltout(),
            .carryin(\nx.n10865 ),
            .carryout(\nx.n10866 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_5_lut_LC_11_29_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_5_lut_LC_11_29_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_5_lut_LC_11_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_5_lut_LC_11_29_3  (
            .in0(_gnd_net_),
            .in1(N__41592),
            .in2(N__30423),
            .in3(N__30402),
            .lcout(\nx.n2174 ),
            .ltout(),
            .carryin(\nx.n10866 ),
            .carryout(\nx.n10867 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_6_lut_LC_11_29_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_6_lut_LC_11_29_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_6_lut_LC_11_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_6_lut_LC_11_29_4  (
            .in0(_gnd_net_),
            .in1(N__30397),
            .in2(N__41974),
            .in3(N__30375),
            .lcout(\nx.n2173 ),
            .ltout(),
            .carryin(\nx.n10867 ),
            .carryout(\nx.n10868 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_7_lut_LC_11_29_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_7_lut_LC_11_29_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_7_lut_LC_11_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_7_lut_LC_11_29_5  (
            .in0(_gnd_net_),
            .in1(N__41596),
            .in2(N__30372),
            .in3(N__30345),
            .lcout(\nx.n2172 ),
            .ltout(),
            .carryin(\nx.n10868 ),
            .carryout(\nx.n10869 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_8_lut_LC_11_29_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_8_lut_LC_11_29_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_8_lut_LC_11_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_8_lut_LC_11_29_6  (
            .in0(_gnd_net_),
            .in1(N__42200),
            .in2(N__30342),
            .in3(N__30312),
            .lcout(\nx.n2171 ),
            .ltout(),
            .carryin(\nx.n10869 ),
            .carryout(\nx.n10870 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_9_lut_LC_11_29_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_9_lut_LC_11_29_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_9_lut_LC_11_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_9_lut_LC_11_29_7  (
            .in0(_gnd_net_),
            .in1(N__41597),
            .in2(N__30309),
            .in3(N__30285),
            .lcout(\nx.n2170 ),
            .ltout(),
            .carryin(\nx.n10870 ),
            .carryout(\nx.n10871 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_10_lut_LC_11_30_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_10_lut_LC_11_30_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_10_lut_LC_11_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_10_lut_LC_11_30_0  (
            .in0(_gnd_net_),
            .in1(N__41598),
            .in2(N__32708),
            .in3(N__30732),
            .lcout(\nx.n2169 ),
            .ltout(),
            .carryin(bfn_11_30_0_),
            .carryout(\nx.n10872 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_11_lut_LC_11_30_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_11_lut_LC_11_30_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_11_lut_LC_11_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_11_lut_LC_11_30_1  (
            .in0(_gnd_net_),
            .in1(N__41605),
            .in2(N__36593),
            .in3(N__30729),
            .lcout(\nx.n2168 ),
            .ltout(),
            .carryin(\nx.n10872 ),
            .carryout(\nx.n10873 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_12_lut_LC_11_30_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_12_lut_LC_11_30_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_12_lut_LC_11_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_12_lut_LC_11_30_2  (
            .in0(_gnd_net_),
            .in1(N__41599),
            .in2(N__30726),
            .in3(N__30684),
            .lcout(\nx.n2167 ),
            .ltout(),
            .carryin(\nx.n10873 ),
            .carryout(\nx.n10874 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_13_lut_LC_11_30_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_13_lut_LC_11_30_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_13_lut_LC_11_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_13_lut_LC_11_30_3  (
            .in0(_gnd_net_),
            .in1(N__41606),
            .in2(N__32166),
            .in3(N__30681),
            .lcout(\nx.n2166 ),
            .ltout(),
            .carryin(\nx.n10874 ),
            .carryout(\nx.n10875 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_14_lut_LC_11_30_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_14_lut_LC_11_30_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_14_lut_LC_11_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_14_lut_LC_11_30_4  (
            .in0(_gnd_net_),
            .in1(N__41600),
            .in2(N__30678),
            .in3(N__30639),
            .lcout(\nx.n2165 ),
            .ltout(),
            .carryin(\nx.n10875 ),
            .carryout(\nx.n10876 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_15_lut_LC_11_30_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_15_lut_LC_11_30_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_15_lut_LC_11_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_15_lut_LC_11_30_5  (
            .in0(_gnd_net_),
            .in1(N__30635),
            .in2(N__41975),
            .in3(N__30603),
            .lcout(\nx.n2164 ),
            .ltout(),
            .carryin(\nx.n10876 ),
            .carryout(\nx.n10877 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_16_lut_LC_11_30_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_16_lut_LC_11_30_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_16_lut_LC_11_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_16_lut_LC_11_30_6  (
            .in0(_gnd_net_),
            .in1(N__41604),
            .in2(N__30600),
            .in3(N__30573),
            .lcout(\nx.n2163 ),
            .ltout(),
            .carryin(\nx.n10877 ),
            .carryout(\nx.n10878 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_17_lut_LC_11_30_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_17_lut_LC_11_30_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_17_lut_LC_11_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_17_lut_LC_11_30_7  (
            .in0(_gnd_net_),
            .in1(N__41607),
            .in2(N__30569),
            .in3(N__30537),
            .lcout(\nx.n2162 ),
            .ltout(),
            .carryin(\nx.n10878 ),
            .carryout(\nx.n10879 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_18_lut_LC_11_31_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1473_18_lut_LC_11_31_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_18_lut_LC_11_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1473_18_lut_LC_11_31_0  (
            .in0(_gnd_net_),
            .in1(N__41608),
            .in2(N__30894),
            .in3(N__30864),
            .lcout(\nx.n2161 ),
            .ltout(),
            .carryin(bfn_11_31_0_),
            .carryout(\nx.n10880 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1473_19_lut_LC_11_31_1 .C_ON=1'b0;
    defparam \nx.mod_5_add_1473_19_lut_LC_11_31_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1473_19_lut_LC_11_31_1 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1473_19_lut_LC_11_31_1  (
            .in0(N__41609),
            .in1(N__30861),
            .in2(N__36561),
            .in3(N__30843),
            .lcout(\nx.n2192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2166_3_lut_LC_12_17_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2166_3_lut_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2166_3_lut_LC_12_17_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i2166_3_lut_LC_12_17_0  (
            .in0(N__32856),
            .in1(_gnd_net_),
            .in2(N__34005),
            .in3(N__32884),
            .lcout(),
            .ltout(\nx.n21_adj_750_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_93_LC_12_17_1 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_93_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_93_LC_12_17_1 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \nx.i1_4_lut_adj_93_LC_12_17_1  (
            .in0(N__33248),
            .in1(N__33222),
            .in2(N__30819),
            .in3(N__33977),
            .lcout(),
            .ltout(\nx.n12781_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_97_LC_12_17_2 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_97_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_97_LC_12_17_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \nx.i1_4_lut_adj_97_LC_12_17_2  (
            .in0(N__30816),
            .in1(N__30743),
            .in2(N__30762),
            .in3(N__30990),
            .lcout(\nx.n12801 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2163_3_lut_LC_12_17_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2163_3_lut_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2163_3_lut_LC_12_17_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2163_3_lut_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__32727),
            .in2(N__32769),
            .in3(N__33967),
            .lcout(),
            .ltout(\nx.n27_adj_744_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_89_LC_12_17_4 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_89_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_89_LC_12_17_4 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \nx.i1_4_lut_adj_89_LC_12_17_4  (
            .in0(N__33968),
            .in1(N__33306),
            .in2(N__30750),
            .in3(N__33329),
            .lcout(\nx.n12779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2172_3_lut_LC_12_17_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2172_3_lut_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2172_3_lut_LC_12_17_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i2172_3_lut_LC_12_17_5  (
            .in0(N__32370),
            .in1(N__32412),
            .in2(_gnd_net_),
            .in3(N__33972),
            .lcout(\nx.n3209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2164_3_lut_LC_12_17_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2164_3_lut_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2164_3_lut_LC_12_17_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2164_3_lut_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(N__32798),
            .in2(N__34004),
            .in3(N__32778),
            .lcout(),
            .ltout(\nx.n25_adj_748_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_92_LC_12_17_7 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_92_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_92_LC_12_17_7 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \nx.i1_4_lut_adj_92_LC_12_17_7  (
            .in0(N__33180),
            .in1(N__33209),
            .in2(N__30993),
            .in3(N__33973),
            .lcout(\nx.n12785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_88_LC_12_18_0 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_88_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_88_LC_12_18_0 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \nx.i1_4_lut_adj_88_LC_12_18_0  (
            .in0(N__32811),
            .in1(N__32833),
            .in2(N__34001),
            .in3(N__30984),
            .lcout(),
            .ltout(\nx.n12777_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_91_LC_12_18_1 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_91_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_91_LC_12_18_1 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \nx.i1_4_lut_adj_91_LC_12_18_1  (
            .in0(N__32985),
            .in1(N__33005),
            .in2(N__30978),
            .in3(N__33962),
            .lcout(\nx.n12789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2157_3_lut_LC_12_18_2 .C_ON=1'b0;
    defparam \nx.mod_5_i2157_3_lut_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2157_3_lut_LC_12_18_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2157_3_lut_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__33141),
            .in2(N__34003),
            .in3(N__33163),
            .lcout(),
            .ltout(\nx.n39_adj_747_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_4_lut_adj_95_LC_12_18_3 .C_ON=1'b0;
    defparam \nx.i1_4_lut_adj_95_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.i1_4_lut_adj_95_LC_12_18_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i1_4_lut_adj_95_LC_12_18_3  (
            .in0(N__30951),
            .in1(N__30975),
            .in2(N__30969),
            .in3(N__30966),
            .lcout(\nx.n12799 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2162_3_lut_LC_12_18_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2162_3_lut_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2162_3_lut_LC_12_18_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2162_3_lut_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__33345),
            .in2(N__34002),
            .in3(N__33365),
            .lcout(\nx.n29_adj_746 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2171_3_lut_LC_12_18_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2171_3_lut_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2171_3_lut_LC_12_18_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2171_3_lut_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__32325),
            .in2(N__32354),
            .in3(N__33955),
            .lcout(\nx.n11_adj_751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2156_3_lut_LC_12_18_7 .C_ON=1'b0;
    defparam \nx.mod_5_i2156_3_lut_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2156_3_lut_LC_12_18_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2156_3_lut_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__33124),
            .in2(N__33105),
            .in3(N__33966),
            .lcout(\nx.n41_adj_752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2016_3_lut_LC_12_19_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2016_3_lut_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2016_3_lut_LC_12_19_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2016_3_lut_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__35673),
            .in2(N__37103),
            .in3(N__37298),
            .lcout(\nx.n2989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2027_3_lut_LC_12_19_2 .C_ON=1'b0;
    defparam \nx.mod_5_i2027_3_lut_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2027_3_lut_LC_12_19_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2027_3_lut_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__35462),
            .in2(N__35430),
            .in3(N__37294),
            .lcout(\nx.n3000 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2028_3_lut_LC_12_19_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2028_3_lut_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2028_3_lut_LC_12_19_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2028_3_lut_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__35515),
            .in2(N__35481),
            .in3(N__37299),
            .lcout(\nx.n3001 ),
            .ltout(\nx.n3001_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_125_LC_12_19_5 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_125_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_125_LC_12_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_125_LC_12_19_5  (
            .in0(N__31066),
            .in1(N__31048),
            .in2(N__31080),
            .in3(N__35836),
            .lcout(\nx.n44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2030_3_lut_LC_12_19_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2030_3_lut_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2030_3_lut_LC_12_19_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2030_3_lut_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__37417),
            .in2(N__35001),
            .in3(N__37293),
            .lcout(\nx.n3003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2032_3_lut_LC_12_19_7 .C_ON=1'b0;
    defparam \nx.mod_5_i2032_3_lut_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2032_3_lut_LC_12_19_7 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \nx.mod_5_i2032_3_lut_LC_12_19_7  (
            .in0(N__35069),
            .in1(N__35040),
            .in2(N__37320),
            .in3(_gnd_net_),
            .lcout(\nx.n3005 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_113_LC_12_20_0 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_113_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_113_LC_12_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_113_LC_12_20_0  (
            .in0(N__35560),
            .in1(N__35612),
            .in2(N__36904),
            .in3(N__35282),
            .lcout(\nx.n39_adj_761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1954_3_lut_LC_12_20_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1954_3_lut_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1954_3_lut_LC_12_20_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1954_3_lut_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__31138),
            .in2(N__31032),
            .in3(N__37588),
            .lcout(\nx.n2895 ),
            .ltout(\nx.n2895_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2021_3_lut_LC_12_20_2 .C_ON=1'b0;
    defparam \nx.mod_5_i2021_3_lut_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2021_3_lut_LC_12_20_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2021_3_lut_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__35271),
            .in2(N__31017),
            .in3(N__37318),
            .lcout(\nx.n2994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_196_LC_12_20_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_196_LC_12_20_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_196_LC_12_20_3.LUT_INIT=16'b0001000100000000;
    LogicCell40 i1_2_lut_3_lut_adj_196_LC_12_20_3 (
            .in0(N__43925),
            .in1(N__47594),
            .in2(_gnd_net_),
            .in3(N__43681),
            .lcout(n7992),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1957_3_lut_LC_12_20_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1957_3_lut_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1957_3_lut_LC_12_20_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1957_3_lut_LC_12_20_4  (
            .in0(N__31439),
            .in1(_gnd_net_),
            .in2(N__37606),
            .in3(N__31413),
            .lcout(\nx.n2898 ),
            .ltout(\nx.n2898_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2024_3_lut_LC_12_20_5 .C_ON=1'b0;
    defparam \nx.mod_5_i2024_3_lut_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2024_3_lut_LC_12_20_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \nx.mod_5_i2024_3_lut_LC_12_20_5  (
            .in0(N__37319),
            .in1(_gnd_net_),
            .in2(N__31401),
            .in3(N__35319),
            .lcout(\nx.n2997 ),
            .ltout(\nx.n2997_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_LC_12_20_6 .C_ON=1'b0;
    defparam \nx.i19_4_lut_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_LC_12_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_LC_12_20_6  (
            .in0(N__33719),
            .in1(N__33745),
            .in2(N__31386),
            .in3(N__31369),
            .lcout(\nx.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2015_3_lut_LC_12_21_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2015_3_lut_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2015_3_lut_LC_12_21_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2015_3_lut_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__35657),
            .in2(N__35637),
            .in3(N__37312),
            .lcout(\nx.n2988 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1946_3_lut_LC_12_21_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1946_3_lut_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1946_3_lut_LC_12_21_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1946_3_lut_LC_12_21_2  (
            .in0(N__31353),
            .in1(_gnd_net_),
            .in2(N__31341),
            .in3(N__37607),
            .lcout(\nx.n2887 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1815_3_lut_LC_12_21_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1815_3_lut_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1815_3_lut_LC_12_21_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1815_3_lut_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(N__39471),
            .in2(N__39501),
            .in3(N__40106),
            .lcout(\nx.n2692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1887_3_lut_LC_12_21_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1887_3_lut_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1887_3_lut_LC_12_21_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1887_3_lut_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__31320),
            .in2(N__31308),
            .in3(N__31274),
            .lcout(\nx.n2796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_16_LC_12_21_7 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_16_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_16_LC_12_21_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_16_LC_12_21_7  (
            .in0(N__39251),
            .in1(N__39169),
            .in2(N__39306),
            .in3(N__39124),
            .lcout(\nx.n38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1757_rep_22_3_lut_LC_12_22_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1757_rep_22_3_lut_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1757_rep_22_3_lut_LC_12_22_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1757_rep_22_3_lut_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(N__40374),
            .in2(N__40347),
            .in3(N__40914),
            .lcout(\nx.n2602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1752_3_lut_LC_12_22_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1752_3_lut_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1752_3_lut_LC_12_22_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1752_3_lut_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__40729),
            .in2(N__40927),
            .in3(N__40707),
            .lcout(\nx.n2597 ),
            .ltout(\nx.n2597_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_17_LC_12_22_3 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_17_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_17_LC_12_22_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_17_LC_12_22_3  (
            .in0(N__39214),
            .in1(N__39727),
            .in2(N__31641),
            .in3(N__39079),
            .lcout(\nx.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1814_3_lut_LC_12_22_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1814_3_lut_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1814_3_lut_LC_12_22_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1814_3_lut_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(N__39453),
            .in2(N__39435),
            .in3(N__40079),
            .lcout(\nx.n2691 ),
            .ltout(\nx.n2691_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_24_LC_12_22_5 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_24_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_24_LC_12_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_24_LC_12_22_5  (
            .in0(N__31459),
            .in1(N__31594),
            .in2(N__31578),
            .in3(N__31558),
            .lcout(\nx.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9151_3_lut_LC_12_22_6 .C_ON=1'b0;
    defparam \nx.i9151_3_lut_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.i9151_3_lut_LC_12_22_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.i9151_3_lut_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(N__39173),
            .in2(N__39153),
            .in3(N__40078),
            .lcout(\nx.n2700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1811_3_lut_LC_12_23_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1811_3_lut_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1811_3_lut_LC_12_23_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1811_3_lut_LC_12_23_0  (
            .in0(N__39951),
            .in1(_gnd_net_),
            .in2(N__40091),
            .in3(N__40119),
            .lcout(\nx.n2688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1812_3_lut_LC_12_23_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1812_3_lut_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1812_3_lut_LC_12_23_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1812_3_lut_LC_12_23_1  (
            .in0(N__40159),
            .in1(_gnd_net_),
            .in2(N__40134),
            .in3(N__40047),
            .lcout(\nx.n2689 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_LC_12_23_3 .C_ON=1'b0;
    defparam \nx.i12_4_lut_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_LC_12_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_LC_12_23_3  (
            .in0(N__40802),
            .in1(N__39400),
            .in2(N__40163),
            .in3(N__39950),
            .lcout(),
            .ltout(\nx.n34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_3_lut_LC_12_23_4 .C_ON=1'b0;
    defparam \nx.i17_3_lut_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.i17_3_lut_LC_12_23_4 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \nx.i17_3_lut_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__39342),
            .in2(N__31443),
            .in3(N__39372),
            .lcout(),
            .ltout(\nx.n39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i21_4_lut_LC_12_23_5 .C_ON=1'b0;
    defparam \nx.i21_4_lut_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.i21_4_lut_LC_12_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i21_4_lut_LC_12_23_5  (
            .in0(N__31839),
            .in1(N__31830),
            .in2(N__31824),
            .in3(N__37146),
            .lcout(\nx.n2621 ),
            .ltout(\nx.n2621_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1831_rep_15_3_lut_LC_12_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1831_rep_15_3_lut_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1831_rep_15_3_lut_LC_12_23_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1831_rep_15_3_lut_LC_12_23_6  (
            .in0(N__38844),
            .in1(_gnd_net_),
            .in2(N__31821),
            .in3(N__38865),
            .lcout(\nx.n2708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1830_3_lut_LC_12_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1830_3_lut_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1830_3_lut_LC_12_23_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1830_3_lut_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(N__38829),
            .in2(N__38802),
            .in3(N__40046),
            .lcout(\nx.n2707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1560_3_lut_LC_12_24_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1560_3_lut_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1560_3_lut_LC_12_24_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i1560_3_lut_LC_12_24_0  (
            .in0(N__31790),
            .in1(N__31746),
            .in2(_gnd_net_),
            .in3(N__32561),
            .lcout(\nx.n2309 ),
            .ltout(\nx.n2309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5904_2_lut_LC_12_24_1 .C_ON=1'b0;
    defparam \nx.i5904_2_lut_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.i5904_2_lut_LC_12_24_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \nx.i5904_2_lut_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31740),
            .in3(N__34329),
            .lcout(),
            .ltout(\nx.n9697_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_54_LC_12_24_2 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_54_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_54_LC_12_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_54_LC_12_24_2  (
            .in0(N__34528),
            .in1(N__37898),
            .in2(N__31737),
            .in3(N__34249),
            .lcout(\nx.n32_adj_698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1556_3_lut_LC_12_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1556_3_lut_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1556_3_lut_LC_12_24_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1556_3_lut_LC_12_24_3  (
            .in0(_gnd_net_),
            .in1(N__31734),
            .in2(N__32578),
            .in3(N__31728),
            .lcout(\nx.n2305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1559_3_lut_LC_12_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1559_3_lut_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1559_3_lut_LC_12_24_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1559_3_lut_LC_12_24_4  (
            .in0(_gnd_net_),
            .in1(N__31704),
            .in2(N__31677),
            .in3(N__32562),
            .lcout(\nx.n2308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1818_3_lut_LC_12_24_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1818_3_lut_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1818_3_lut_LC_12_24_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1818_3_lut_LC_12_24_5  (
            .in0(_gnd_net_),
            .in1(N__39648),
            .in2(N__39618),
            .in3(N__40076),
            .lcout(\nx.n2695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1746_3_lut_LC_12_24_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1746_3_lut_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1746_3_lut_LC_12_24_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1746_3_lut_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(N__40527),
            .in2(N__40500),
            .in3(N__40928),
            .lcout(\nx.n2591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_55_LC_12_25_0 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_55_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_55_LC_12_25_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_55_LC_12_25_0  (
            .in0(N__36415),
            .in1(N__34469),
            .in2(N__34572),
            .in3(N__34442),
            .lcout(\nx.n33_adj_699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1554_3_lut_LC_12_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1554_3_lut_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1554_3_lut_LC_12_25_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1554_3_lut_LC_12_25_1  (
            .in0(_gnd_net_),
            .in1(N__31956),
            .in2(N__31923),
            .in3(N__32572),
            .lcout(\nx.n2303 ),
            .ltout(\nx.n2303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1621_3_lut_LC_12_25_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1621_3_lut_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1621_3_lut_LC_12_25_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1621_3_lut_LC_12_25_2  (
            .in0(N__34455),
            .in1(_gnd_net_),
            .in2(N__31914),
            .in3(N__37987),
            .lcout(\nx.n2402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1552_3_lut_LC_12_25_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1552_3_lut_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1552_3_lut_LC_12_25_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1552_3_lut_LC_12_25_4  (
            .in0(_gnd_net_),
            .in1(N__31911),
            .in2(N__32580),
            .in3(N__31905),
            .lcout(\nx.n2301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1553_3_lut_LC_12_25_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1553_3_lut_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1553_3_lut_LC_12_25_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1553_3_lut_LC_12_25_5  (
            .in0(_gnd_net_),
            .in1(N__31884),
            .in2(N__31854),
            .in3(N__32571),
            .lcout(\nx.n2302 ),
            .ltout(\nx.n2302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1620_3_lut_LC_12_25_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1620_3_lut_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1620_3_lut_LC_12_25_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1620_3_lut_LC_12_25_6  (
            .in0(N__34428),
            .in1(_gnd_net_),
            .in2(N__31845),
            .in3(N__37988),
            .lcout(\nx.n2401 ),
            .ltout(\nx.n2401_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i14_4_lut_adj_58_LC_12_25_7 .C_ON=1'b0;
    defparam \nx.i14_4_lut_adj_58_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.i14_4_lut_adj_58_LC_12_25_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i14_4_lut_adj_58_LC_12_25_7  (
            .in0(N__35936),
            .in1(N__36274),
            .in2(N__31842),
            .in3(N__36202),
            .lcout(\nx.n34_adj_701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1612_3_lut_LC_12_26_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1612_3_lut_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1612_3_lut_LC_12_26_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1612_3_lut_LC_12_26_0  (
            .in0(N__34678),
            .in1(_gnd_net_),
            .in2(N__38015),
            .in3(N__34656),
            .lcout(\nx.n2393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1557_3_lut_LC_12_26_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1557_3_lut_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1557_3_lut_LC_12_26_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1557_3_lut_LC_12_26_1  (
            .in0(N__32112),
            .in1(_gnd_net_),
            .in2(N__32569),
            .in3(N__32105),
            .lcout(\nx.n2306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1558_3_lut_LC_12_26_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1558_3_lut_LC_12_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1558_3_lut_LC_12_26_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1558_3_lut_LC_12_26_2  (
            .in0(N__32073),
            .in1(_gnd_net_),
            .in2(N__32043),
            .in3(N__32538),
            .lcout(\nx.n2307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1555_3_lut_LC_12_26_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1555_3_lut_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1555_3_lut_LC_12_26_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1555_3_lut_LC_12_26_3  (
            .in0(N__32031),
            .in1(_gnd_net_),
            .in2(N__32570),
            .in3(N__32024),
            .lcout(\nx.n2304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1610_3_lut_LC_12_26_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1610_3_lut_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1610_3_lut_LC_12_26_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1610_3_lut_LC_12_26_4  (
            .in0(_gnd_net_),
            .in1(N__34601),
            .in2(N__38016),
            .in3(N__34587),
            .lcout(\nx.n2391 ),
            .ltout(\nx.n2391_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_62_LC_12_26_5 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_62_LC_12_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_62_LC_12_26_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_62_LC_12_26_5  (
            .in0(N__36359),
            .in1(N__38573),
            .in2(N__31992),
            .in3(N__38518),
            .lcout(\nx.n31_adj_707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i11_4_lut_adj_52_LC_12_26_6 .C_ON=1'b0;
    defparam \nx.i11_4_lut_adj_52_LC_12_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.i11_4_lut_adj_52_LC_12_26_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i11_4_lut_adj_52_LC_12_26_6  (
            .in0(N__36307),
            .in1(N__34643),
            .in2(N__34680),
            .in3(N__34717),
            .lcout(),
            .ltout(\nx.n30_adj_696_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_53_LC_12_26_7 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_53_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_53_LC_12_26_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_53_LC_12_26_7  (
            .in0(N__34600),
            .in1(N__34498),
            .in2(N__31989),
            .in3(N__34973),
            .lcout(\nx.n34_adj_697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1549_3_lut_LC_12_27_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1549_3_lut_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1549_3_lut_LC_12_27_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1549_3_lut_LC_12_27_0  (
            .in0(_gnd_net_),
            .in1(N__31986),
            .in2(N__31980),
            .in3(N__32554),
            .lcout(\nx.n2298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1550_3_lut_LC_12_27_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1550_3_lut_LC_12_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1550_3_lut_LC_12_27_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1550_3_lut_LC_12_27_1  (
            .in0(_gnd_net_),
            .in1(N__31962),
            .in2(N__32577),
            .in3(N__36454),
            .lcout(\nx.n2299 ),
            .ltout(\nx.n2299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_56_LC_12_27_2 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_56_LC_12_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_56_LC_12_27_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_56_LC_12_27_2  (
            .in0(N__34405),
            .in1(N__36664),
            .in2(N__32316),
            .in3(N__36631),
            .lcout(\nx.n31_adj_700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1611_3_lut_LC_12_27_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1611_3_lut_LC_12_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1611_3_lut_LC_12_27_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1611_3_lut_LC_12_27_3  (
            .in0(N__34642),
            .in1(_gnd_net_),
            .in2(N__38021),
            .in3(N__34620),
            .lcout(\nx.n2392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1548_3_lut_LC_12_27_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1548_3_lut_LC_12_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1548_3_lut_LC_12_27_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1548_3_lut_LC_12_27_4  (
            .in0(_gnd_net_),
            .in1(N__32132),
            .in2(N__32313),
            .in3(N__32553),
            .lcout(\nx.n2297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i3_2_lut_LC_12_27_5 .C_ON=1'b0;
    defparam \nx.i3_2_lut_LC_12_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.i3_2_lut_LC_12_27_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \nx.i3_2_lut_LC_12_27_5  (
            .in0(_gnd_net_),
            .in1(N__32290),
            .in2(_gnd_net_),
            .in3(N__32270),
            .lcout(),
            .ltout(\nx.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_51_LC_12_27_6 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_51_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_51_LC_12_27_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_51_LC_12_27_6  (
            .in0(N__32259),
            .in1(N__32253),
            .in2(N__32241),
            .in3(N__32238),
            .lcout(\nx.n2225 ),
            .ltout(\nx.n2225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1551_3_lut_LC_12_27_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1551_3_lut_LC_12_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1551_3_lut_LC_12_27_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1551_3_lut_LC_12_27_7  (
            .in0(N__32232),
            .in1(_gnd_net_),
            .in2(N__32226),
            .in3(N__32669),
            .lcout(\nx.n2300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam neopxl_color_i4_LC_12_28_0.C_ON=1'b0;
    defparam neopxl_color_i4_LC_12_28_0.SEQ_MODE=4'b1001;
    defparam neopxl_color_i4_LC_12_28_0.LUT_INIT=16'b0000000011101010;
    LogicCell40 neopxl_color_i4_LC_12_28_0 (
            .in0(N__32203),
            .in1(N__47693),
            .in2(N__43956),
            .in3(N__43711),
            .lcout(neopxl_color_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46916),
            .ce(),
            .sr(N__32181));
    defparam \nx.mod_5_i1481_3_lut_LC_12_28_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1481_3_lut_LC_12_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1481_3_lut_LC_12_28_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1481_3_lut_LC_12_28_1  (
            .in0(_gnd_net_),
            .in1(N__32162),
            .in2(N__36564),
            .in3(N__32142),
            .lcout(\nx.n2198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1484_3_lut_LC_12_28_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1484_3_lut_LC_12_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1484_3_lut_LC_12_28_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1484_3_lut_LC_12_28_2  (
            .in0(_gnd_net_),
            .in1(N__32718),
            .in2(N__32709),
            .in3(N__36553),
            .lcout(\nx.n2201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1544_3_lut_LC_12_28_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1544_3_lut_LC_12_28_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1544_3_lut_LC_12_28_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1544_3_lut_LC_12_28_6  (
            .in0(_gnd_net_),
            .in1(N__32649),
            .in2(N__32576),
            .in3(N__32642),
            .lcout(\nx.n2293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1545_3_lut_LC_12_28_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1545_3_lut_LC_12_28_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1545_3_lut_LC_12_28_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1545_3_lut_LC_12_28_7  (
            .in0(_gnd_net_),
            .in1(N__32622),
            .in2(N__32613),
            .in3(N__32552),
            .lcout(\nx.n2294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i4_LC_13_15_0.C_ON=1'b0;
    defparam pin_output_enable__i4_LC_13_15_0.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i4_LC_13_15_0.LUT_INIT=16'b1101100011001100;
    LogicCell40 pin_output_enable__i4_LC_13_15_0 (
            .in0(N__37119),
            .in1(N__32462),
            .in2(N__47657),
            .in3(N__47072),
            .lcout(pin_oe_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46881),
            .ce(),
            .sr(_gnd_net_));
    defparam i7633_2_lut_3_lut_4_lut_4_lut_LC_13_16_2.C_ON=1'b0;
    defparam i7633_2_lut_3_lut_4_lut_4_lut_LC_13_16_2.SEQ_MODE=4'b0000;
    defparam i7633_2_lut_3_lut_4_lut_4_lut_LC_13_16_2.LUT_INIT=16'b1111111000000000;
    LogicCell40 i7633_2_lut_3_lut_4_lut_4_lut_LC_13_16_2 (
            .in0(N__42614),
            .in1(N__44106),
            .in2(N__45649),
            .in3(N__47549),
            .lcout(),
            .ltout(n11970_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i0_LC_13_16_3.C_ON=1'b0;
    defparam pin_output_enable__i0_LC_13_16_3.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i0_LC_13_16_3.LUT_INIT=16'b1010110010101010;
    LogicCell40 pin_output_enable__i0_LC_13_16_3 (
            .in0(N__32435),
            .in1(N__47581),
            .in2(N__32451),
            .in3(N__47146),
            .lcout(pin_oe_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46877),
            .ce(),
            .sr(_gnd_net_));
    defparam i7631_3_lut_4_lut_4_lut_LC_13_16_7.C_ON=1'b0;
    defparam i7631_3_lut_4_lut_4_lut_LC_13_16_7.SEQ_MODE=4'b0000;
    defparam i7631_3_lut_4_lut_4_lut_LC_13_16_7.LUT_INIT=16'b1111000001110000;
    LogicCell40 i7631_3_lut_4_lut_4_lut_LC_13_16_7 (
            .in0(N__43429),
            .in1(N__45592),
            .in2(N__47635),
            .in3(N__42613),
            .lcout(n11968),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_2_lut_LC_13_17_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_2_lut_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_2_lut_LC_13_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_2_lut_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__32411),
            .in2(_gnd_net_),
            .in3(N__32361),
            .lcout(\nx.n3177 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\nx.n11079 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_3_lut_LC_13_17_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_3_lut_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_3_lut_LC_13_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_3_lut_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32358),
            .in3(N__32319),
            .lcout(\nx.n3176 ),
            .ltout(),
            .carryin(\nx.n11079 ),
            .carryout(\nx.n11080 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_4_lut_LC_13_17_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_4_lut_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_4_lut_LC_13_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_4_lut_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__41308),
            .in2(N__33054),
            .in3(N__33015),
            .lcout(\nx.n3175 ),
            .ltout(),
            .carryin(\nx.n11080 ),
            .carryout(\nx.n11081 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_5_lut_LC_13_17_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_5_lut_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_5_lut_LC_13_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_5_lut_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__41314),
            .in2(N__33012),
            .in3(N__32979),
            .lcout(\nx.n3174 ),
            .ltout(),
            .carryin(\nx.n11081 ),
            .carryout(\nx.n11082 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_6_lut_LC_13_17_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_6_lut_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_6_lut_LC_13_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_6_lut_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__41309),
            .in2(N__32976),
            .in3(N__32934),
            .lcout(\nx.n3173 ),
            .ltout(),
            .carryin(\nx.n11082 ),
            .carryout(\nx.n11083 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_7_lut_LC_13_17_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_7_lut_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_7_lut_LC_13_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_7_lut_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__41315),
            .in2(N__32931),
            .in3(N__32895),
            .lcout(\nx.n3172 ),
            .ltout(),
            .carryin(\nx.n11083 ),
            .carryout(\nx.n11084 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_8_lut_LC_13_17_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_8_lut_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_8_lut_LC_13_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_8_lut_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__41310),
            .in2(N__32892),
            .in3(N__32850),
            .lcout(\nx.n3171 ),
            .ltout(),
            .carryin(\nx.n11084 ),
            .carryout(\nx.n11085 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_9_lut_LC_13_17_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_9_lut_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_9_lut_LC_13_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_9_lut_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__32843),
            .in2(N__41638),
            .in3(N__32805),
            .lcout(\nx.n3170 ),
            .ltout(),
            .carryin(\nx.n11085 ),
            .carryout(\nx.n11086 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_10_lut_LC_13_18_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_10_lut_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_10_lut_LC_13_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_10_lut_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__41472),
            .in2(N__32802),
            .in3(N__32772),
            .lcout(\nx.n3169 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\nx.n11087 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_11_lut_LC_13_18_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_11_lut_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_11_lut_LC_13_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_11_lut_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__41476),
            .in2(N__32768),
            .in3(N__32721),
            .lcout(\nx.n3168 ),
            .ltout(),
            .carryin(\nx.n11087 ),
            .carryout(\nx.n11088 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_12_lut_LC_13_18_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_12_lut_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_12_lut_LC_13_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_12_lut_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__41473),
            .in2(N__33372),
            .in3(N__33339),
            .lcout(\nx.n3167 ),
            .ltout(),
            .carryin(\nx.n11088 ),
            .carryout(\nx.n11089 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_13_lut_LC_13_18_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_13_lut_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_13_lut_LC_13_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_13_lut_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__41477),
            .in2(N__33336),
            .in3(N__33300),
            .lcout(\nx.n3166 ),
            .ltout(),
            .carryin(\nx.n11089 ),
            .carryout(\nx.n11090 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_14_lut_LC_13_18_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_14_lut_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_14_lut_LC_13_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_14_lut_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__41474),
            .in2(N__33297),
            .in3(N__33255),
            .lcout(\nx.n3165 ),
            .ltout(),
            .carryin(\nx.n11090 ),
            .carryout(\nx.n11091 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_15_lut_LC_13_18_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_15_lut_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_15_lut_LC_13_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_15_lut_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__41478),
            .in2(N__33252),
            .in3(N__33216),
            .lcout(\nx.n3164 ),
            .ltout(),
            .carryin(\nx.n11091 ),
            .carryout(\nx.n11092 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_16_lut_LC_13_18_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_16_lut_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_16_lut_LC_13_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_16_lut_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__41475),
            .in2(N__33213),
            .in3(N__33174),
            .lcout(\nx.n3163 ),
            .ltout(),
            .carryin(\nx.n11092 ),
            .carryout(\nx.n11093 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_17_lut_LC_13_18_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_17_lut_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_17_lut_LC_13_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_17_lut_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__41479),
            .in2(N__33171),
            .in3(N__33135),
            .lcout(\nx.n3162 ),
            .ltout(),
            .carryin(\nx.n11093 ),
            .carryout(\nx.n11094 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_18_lut_LC_13_19_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_18_lut_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_18_lut_LC_13_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_18_lut_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__33132),
            .in2(N__41862),
            .in3(N__33096),
            .lcout(\nx.n3161 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\nx.n11095 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_19_lut_LC_13_19_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_19_lut_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_19_lut_LC_13_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_19_lut_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__41483),
            .in2(N__33093),
            .in3(N__33696),
            .lcout(\nx.n3160 ),
            .ltout(),
            .carryin(\nx.n11095 ),
            .carryout(\nx.n11096 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_20_lut_LC_13_19_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_20_lut_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_20_lut_LC_13_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_20_lut_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__33693),
            .in2(N__41863),
            .in3(N__33651),
            .lcout(\nx.n3159 ),
            .ltout(),
            .carryin(\nx.n11096 ),
            .carryout(\nx.n11097 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_21_lut_LC_13_19_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_21_lut_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_21_lut_LC_13_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_21_lut_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__33647),
            .in2(N__41866),
            .in3(N__33606),
            .lcout(\nx.n3158 ),
            .ltout(),
            .carryin(\nx.n11097 ),
            .carryout(\nx.n11098 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_22_lut_LC_13_19_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_22_lut_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_22_lut_LC_13_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_22_lut_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__33602),
            .in2(N__41864),
            .in3(N__33561),
            .lcout(\nx.n3157 ),
            .ltout(),
            .carryin(\nx.n11098 ),
            .carryout(\nx.n11099 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_23_lut_LC_13_19_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_23_lut_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_23_lut_LC_13_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_23_lut_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__33558),
            .in2(N__41867),
            .in3(N__33519),
            .lcout(\nx.n3156 ),
            .ltout(),
            .carryin(\nx.n11099 ),
            .carryout(\nx.n11100 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_24_lut_LC_13_19_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_24_lut_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_24_lut_LC_13_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_24_lut_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__33515),
            .in2(N__41865),
            .in3(N__33471),
            .lcout(\nx.n3155 ),
            .ltout(),
            .carryin(\nx.n11100 ),
            .carryout(\nx.n11101 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_25_lut_LC_13_19_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_25_lut_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_25_lut_LC_13_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_25_lut_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__33467),
            .in2(N__41868),
            .in3(N__33420),
            .lcout(\nx.n3154 ),
            .ltout(),
            .carryin(\nx.n11101 ),
            .carryout(\nx.n11102 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_26_lut_LC_13_20_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_26_lut_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_26_lut_LC_13_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_26_lut_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__33413),
            .in2(N__42120),
            .in3(N__33375),
            .lcout(\nx.n3153 ),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(\nx.n11103 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_27_lut_LC_13_20_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_27_lut_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_27_lut_LC_13_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_27_lut_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__34127),
            .in2(N__42122),
            .in3(N__34083),
            .lcout(\nx.n3152 ),
            .ltout(),
            .carryin(\nx.n11103 ),
            .carryout(\nx.n11104 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_28_lut_LC_13_20_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2143_28_lut_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_28_lut_LC_13_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2143_28_lut_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__34079),
            .in2(N__42121),
            .in3(N__34035),
            .lcout(\nx.n3151 ),
            .ltout(),
            .carryin(\nx.n11104 ),
            .carryout(\nx.n11105 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2143_29_lut_LC_13_20_3 .C_ON=1'b0;
    defparam \nx.mod_5_add_2143_29_lut_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2143_29_lut_LC_13_20_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \nx.mod_5_add_2143_29_lut_LC_13_20_3  (
            .in0(N__34026),
            .in1(N__41875),
            .in2(N__33891),
            .in3(N__33864),
            .lcout(\nx.n13280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1963_3_lut_LC_13_20_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1963_3_lut_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1963_3_lut_LC_13_20_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1963_3_lut_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__33849),
            .in2(N__33819),
            .in3(N__37579),
            .lcout(\nx.n2904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1956_3_lut_LC_13_20_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1956_3_lut_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1956_3_lut_LC_13_20_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1956_3_lut_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__33803),
            .in2(N__33771),
            .in3(N__37580),
            .lcout(\nx.n2897 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2013_3_lut_LC_13_21_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2013_3_lut_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2013_3_lut_LC_13_21_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2013_3_lut_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__35570),
            .in2(N__35547),
            .in3(N__37306),
            .lcout(\nx.n2986 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1826_rep_14_3_lut_LC_13_21_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1826_rep_14_3_lut_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1826_rep_14_3_lut_LC_13_21_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1826_rep_14_3_lut_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__39304),
            .in2(N__39273),
            .in3(N__40105),
            .lcout(\nx.n2703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2018_3_lut_LC_13_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2018_3_lut_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2018_3_lut_LC_13_21_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2018_3_lut_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__35685),
            .in2(N__37725),
            .in3(N__37305),
            .lcout(\nx.n2991 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1755_3_lut_LC_13_22_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1755_3_lut_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1755_3_lut_LC_13_22_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1755_3_lut_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__40263),
            .in2(N__40283),
            .in3(N__40907),
            .lcout(\nx.n2600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1756_3_lut_LC_13_22_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1756_3_lut_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1756_3_lut_LC_13_22_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1756_3_lut_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__40302),
            .in2(N__40922),
            .in3(N__40322),
            .lcout(\nx.n2601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1758_3_lut_LC_13_22_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1758_3_lut_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1758_3_lut_LC_13_22_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1758_3_lut_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(N__40389),
            .in2(N__40415),
            .in3(N__40903),
            .lcout(\nx.n2603 ),
            .ltout(\nx.n2603_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1825_3_lut_LC_13_22_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1825_3_lut_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1825_3_lut_LC_13_22_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1825_3_lut_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(N__39237),
            .in2(N__34212),
            .in3(N__40077),
            .lcout(\nx.n2702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1961_3_lut_LC_13_22_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1961_3_lut_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1961_3_lut_LC_13_22_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1961_3_lut_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(N__34176),
            .in2(N__34149),
            .in3(N__37597),
            .lcout(\nx.n2902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1685_3_lut_LC_13_22_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1685_3_lut_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1685_3_lut_LC_13_22_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1685_3_lut_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(N__36099),
            .in2(N__36132),
            .in3(N__38478),
            .lcout(\nx.n2498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1687_3_lut_LC_13_23_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1687_3_lut_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1687_3_lut_LC_13_23_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1687_3_lut_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__36147),
            .in2(N__36174),
            .in3(N__38461),
            .lcout(\nx.n2500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1688_3_lut_LC_13_23_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1688_3_lut_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1688_3_lut_LC_13_23_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1688_3_lut_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__36186),
            .in2(N__38497),
            .in3(N__36212),
            .lcout(\nx.n2501 ),
            .ltout(\nx.n2501_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_3_lut_adj_110_LC_13_23_2 .C_ON=1'b0;
    defparam \nx.i6_3_lut_adj_110_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.i6_3_lut_adj_110_LC_13_23_2 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \nx.i6_3_lut_adj_110_LC_13_23_2  (
            .in0(N__39923),
            .in1(_gnd_net_),
            .in2(N__34134),
            .in3(N__39838),
            .lcout(\nx.n27_adj_757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1694_3_lut_LC_13_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1694_3_lut_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1694_3_lut_LC_13_23_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1694_3_lut_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__35979),
            .in2(N__36003),
            .in3(N__38456),
            .lcout(\nx.n2507 ),
            .ltout(\nx.n2507_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_109_LC_13_23_5 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_109_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_109_LC_13_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_109_LC_13_23_5  (
            .in0(N__40321),
            .in1(N__40237),
            .in2(N__34215),
            .in3(N__40408),
            .lcout(\nx.n36_adj_756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1689_rep_26_3_lut_LC_13_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1689_rep_26_3_lut_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1689_rep_26_3_lut_LC_13_23_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1689_rep_26_3_lut_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__36222),
            .in2(N__36249),
            .in3(N__38460),
            .lcout(\nx.n2502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1691_3_lut_LC_13_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1691_3_lut_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1691_3_lut_LC_13_23_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \nx.mod_5_i1691_3_lut_LC_13_23_7  (
            .in0(N__35889),
            .in1(_gnd_net_),
            .in2(N__38496),
            .in3(N__35913),
            .lcout(\nx.n2504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1690_3_lut_LC_13_24_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1690_3_lut_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1690_3_lut_LC_13_24_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1690_3_lut_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__36258),
            .in2(N__36282),
            .in3(N__38474),
            .lcout(\nx.n2503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1626_3_lut_LC_13_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1626_3_lut_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1626_3_lut_LC_13_24_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1626_3_lut_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__34250),
            .in2(N__34230),
            .in3(N__37999),
            .lcout(\nx.n2407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1614_3_lut_LC_13_24_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1614_3_lut_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1614_3_lut_LC_13_24_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1614_3_lut_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__34695),
            .in2(N__34731),
            .in3(N__38000),
            .lcout(\nx.n2395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1627_3_lut_LC_13_24_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1627_3_lut_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1627_3_lut_LC_13_24_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1627_3_lut_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__34266),
            .in2(N__38017),
            .in3(N__34280),
            .lcout(\nx.n2408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1628_3_lut_LC_13_24_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1628_3_lut_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1628_3_lut_LC_13_24_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \nx.mod_5_i1628_3_lut_LC_13_24_7  (
            .in0(N__34296),
            .in1(N__34333),
            .in2(_gnd_net_),
            .in3(N__37995),
            .lcout(\nx.n2409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1623_3_lut_LC_13_25_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1623_3_lut_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1623_3_lut_LC_13_25_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1623_3_lut_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__34509),
            .in2(N__34535),
            .in3(N__37967),
            .lcout(\nx.n2404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1618_3_lut_LC_13_25_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1618_3_lut_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1618_3_lut_LC_13_25_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1618_3_lut_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__34413),
            .in2(N__38008),
            .in3(N__34389),
            .lcout(\nx.n2399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1624_3_lut_LC_13_25_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1624_3_lut_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1624_3_lut_LC_13_25_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1624_3_lut_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(N__34570),
            .in2(N__34548),
            .in3(N__37968),
            .lcout(\nx.n2405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1617_3_lut_LC_13_25_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1617_3_lut_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1617_3_lut_LC_13_25_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1617_3_lut_LC_13_25_3  (
            .in0(N__34767),
            .in1(_gnd_net_),
            .in2(N__38010),
            .in3(N__34749),
            .lcout(\nx.n2398 ),
            .ltout(\nx.n2398_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i15_4_lut_adj_63_LC_13_25_4 .C_ON=1'b0;
    defparam \nx.i15_4_lut_adj_63_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.i15_4_lut_adj_63_LC_13_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i15_4_lut_adj_63_LC_13_25_4  (
            .in0(N__35905),
            .in1(N__35995),
            .in2(N__34377),
            .in3(N__36238),
            .lcout(\nx.n35_adj_708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1622_3_lut_LC_13_25_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1622_3_lut_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1622_3_lut_LC_13_25_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \nx.mod_5_i1622_3_lut_LC_13_25_5  (
            .in0(N__34499),
            .in1(N__34479),
            .in2(N__38009),
            .in3(_gnd_net_),
            .lcout(\nx.n2403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_57_LC_13_25_6 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_57_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_57_LC_13_25_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_57_LC_13_25_6  (
            .in0(N__34374),
            .in1(N__34365),
            .in2(N__34359),
            .in3(N__34350),
            .lcout(\nx.n2324 ),
            .ltout(\nx.n2324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1625_3_lut_LC_13_25_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1625_3_lut_LC_13_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1625_3_lut_LC_13_25_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1625_3_lut_LC_13_25_7  (
            .in0(_gnd_net_),
            .in1(N__36071),
            .in2(N__34344),
            .in3(N__37896),
            .lcout(\nx.n2406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_2_lut_LC_13_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_2_lut_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_2_lut_LC_13_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_2_lut_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__34341),
            .in2(_gnd_net_),
            .in3(N__34287),
            .lcout(\nx.n2377 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\nx.n10899 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_3_lut_LC_13_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_3_lut_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_3_lut_LC_13_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_3_lut_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34284),
            .in3(N__34257),
            .lcout(\nx.n2376 ),
            .ltout(),
            .carryin(\nx.n10899 ),
            .carryout(\nx.n10900 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_4_lut_LC_13_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_4_lut_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_4_lut_LC_13_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_4_lut_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(N__41998),
            .in2(N__34254),
            .in3(N__34218),
            .lcout(\nx.n2375 ),
            .ltout(),
            .carryin(\nx.n10900 ),
            .carryout(\nx.n10901 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_5_lut_LC_13_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_5_lut_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_5_lut_LC_13_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_5_lut_LC_13_26_3  (
            .in0(_gnd_net_),
            .in1(N__42015),
            .in2(N__37897),
            .in3(N__34575),
            .lcout(\nx.n2374 ),
            .ltout(),
            .carryin(\nx.n10901 ),
            .carryout(\nx.n10902 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_6_lut_LC_13_26_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_6_lut_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_6_lut_LC_13_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_6_lut_LC_13_26_4  (
            .in0(_gnd_net_),
            .in1(N__34571),
            .in2(N__42210),
            .in3(N__34539),
            .lcout(\nx.n2373 ),
            .ltout(),
            .carryin(\nx.n10902 ),
            .carryout(\nx.n10903 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_7_lut_LC_13_26_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_7_lut_LC_13_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_7_lut_LC_13_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_7_lut_LC_13_26_5  (
            .in0(_gnd_net_),
            .in1(N__42019),
            .in2(N__34536),
            .in3(N__34503),
            .lcout(\nx.n2372 ),
            .ltout(),
            .carryin(\nx.n10903 ),
            .carryout(\nx.n10904 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_8_lut_LC_13_26_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_8_lut_LC_13_26_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_8_lut_LC_13_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_8_lut_LC_13_26_6  (
            .in0(_gnd_net_),
            .in1(N__41999),
            .in2(N__34500),
            .in3(N__34473),
            .lcout(\nx.n2371 ),
            .ltout(),
            .carryin(\nx.n10904 ),
            .carryout(\nx.n10905 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_9_lut_LC_13_26_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_9_lut_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_9_lut_LC_13_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_9_lut_LC_13_26_7  (
            .in0(_gnd_net_),
            .in1(N__42020),
            .in2(N__34470),
            .in3(N__34449),
            .lcout(\nx.n2370 ),
            .ltout(),
            .carryin(\nx.n10905 ),
            .carryout(\nx.n10906 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_10_lut_LC_13_27_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_10_lut_LC_13_27_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_10_lut_LC_13_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_10_lut_LC_13_27_0  (
            .in0(_gnd_net_),
            .in1(N__42025),
            .in2(N__34446),
            .in3(N__34419),
            .lcout(\nx.n2369 ),
            .ltout(),
            .carryin(bfn_13_27_0_),
            .carryout(\nx.n10907 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_11_lut_LC_13_27_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_11_lut_LC_13_27_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_11_lut_LC_13_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_11_lut_LC_13_27_1  (
            .in0(_gnd_net_),
            .in1(N__41976),
            .in2(N__36422),
            .in3(N__34416),
            .lcout(\nx.n2368 ),
            .ltout(),
            .carryin(\nx.n10907 ),
            .carryout(\nx.n10908 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_12_lut_LC_13_27_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_12_lut_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_12_lut_LC_13_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_12_lut_LC_13_27_2  (
            .in0(_gnd_net_),
            .in1(N__42026),
            .in2(N__34412),
            .in3(N__34380),
            .lcout(\nx.n2367 ),
            .ltout(),
            .carryin(\nx.n10908 ),
            .carryout(\nx.n10909 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_13_lut_LC_13_27_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_13_lut_LC_13_27_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_13_lut_LC_13_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_13_lut_LC_13_27_3  (
            .in0(_gnd_net_),
            .in1(N__34760),
            .in2(N__42211),
            .in3(N__34740),
            .lcout(\nx.n2366 ),
            .ltout(),
            .carryin(\nx.n10909 ),
            .carryout(\nx.n10910 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_14_lut_LC_13_27_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_14_lut_LC_13_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_14_lut_LC_13_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_14_lut_LC_13_27_4  (
            .in0(_gnd_net_),
            .in1(N__42030),
            .in2(N__36638),
            .in3(N__34737),
            .lcout(\nx.n2365 ),
            .ltout(),
            .carryin(\nx.n10910 ),
            .carryout(\nx.n10911 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_15_lut_LC_13_27_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_15_lut_LC_13_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_15_lut_LC_13_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_15_lut_LC_13_27_5  (
            .in0(_gnd_net_),
            .in1(N__41977),
            .in2(N__36671),
            .in3(N__34734),
            .lcout(\nx.n2364 ),
            .ltout(),
            .carryin(\nx.n10911 ),
            .carryout(\nx.n10912 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_16_lut_LC_13_27_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_16_lut_LC_13_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_16_lut_LC_13_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_16_lut_LC_13_27_6  (
            .in0(_gnd_net_),
            .in1(N__42031),
            .in2(N__34730),
            .in3(N__34686),
            .lcout(\nx.n2363 ),
            .ltout(),
            .carryin(\nx.n10912 ),
            .carryout(\nx.n10913 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_17_lut_LC_13_27_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_17_lut_LC_13_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_17_lut_LC_13_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_17_lut_LC_13_27_7  (
            .in0(_gnd_net_),
            .in1(N__41978),
            .in2(N__36318),
            .in3(N__34683),
            .lcout(\nx.n2362 ),
            .ltout(),
            .carryin(\nx.n10913 ),
            .carryout(\nx.n10914 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_18_lut_LC_13_28_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_18_lut_LC_13_28_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_18_lut_LC_13_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_18_lut_LC_13_28_0  (
            .in0(_gnd_net_),
            .in1(N__42212),
            .in2(N__34679),
            .in3(N__34647),
            .lcout(\nx.n2361 ),
            .ltout(),
            .carryin(bfn_13_28_0_),
            .carryout(\nx.n10915 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_19_lut_LC_13_28_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_19_lut_LC_13_28_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_19_lut_LC_13_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_19_lut_LC_13_28_1  (
            .in0(_gnd_net_),
            .in1(N__42215),
            .in2(N__34644),
            .in3(N__34614),
            .lcout(\nx.n2360 ),
            .ltout(),
            .carryin(\nx.n10915 ),
            .carryout(\nx.n10916 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_20_lut_LC_13_28_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1607_20_lut_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_20_lut_LC_13_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1607_20_lut_LC_13_28_2  (
            .in0(_gnd_net_),
            .in1(N__42213),
            .in2(N__34611),
            .in3(N__34578),
            .lcout(\nx.n2359 ),
            .ltout(),
            .carryin(\nx.n10916 ),
            .carryout(\nx.n10917 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1607_21_lut_LC_13_28_3 .C_ON=1'b0;
    defparam \nx.mod_5_add_1607_21_lut_LC_13_28_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1607_21_lut_LC_13_28_3 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_1607_21_lut_LC_13_28_3  (
            .in0(N__42214),
            .in1(N__38004),
            .in2(N__34983),
            .in3(N__34962),
            .lcout(\nx.n2390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2031_3_lut_LC_14_18_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2031_3_lut_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2031_3_lut_LC_14_18_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2031_3_lut_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__35028),
            .in2(N__35013),
            .in3(N__37255),
            .lcout(\nx.n3004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2033_3_lut_LC_14_18_1 .C_ON=1'b0;
    defparam \nx.mod_5_i2033_3_lut_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2033_3_lut_LC_14_18_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i2033_3_lut_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__35079),
            .in2(N__37304),
            .in3(N__35106),
            .lcout(\nx.n3006 ),
            .ltout(\nx.n3006_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_LC_14_18_2 .C_ON=1'b0;
    defparam \nx.i17_4_lut_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_LC_14_18_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_LC_14_18_2  (
            .in0(N__34936),
            .in1(N__34895),
            .in2(N__34923),
            .in3(N__36871),
            .lcout(\nx.n43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2026_3_lut_LC_14_18_3 .C_ON=1'b0;
    defparam \nx.mod_5_i2026_3_lut_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2026_3_lut_LC_14_18_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2026_3_lut_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__35412),
            .in2(N__37303),
            .in3(N__35382),
            .lcout(\nx.n2999 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1955_3_lut_LC_14_18_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1955_3_lut_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1955_3_lut_LC_14_18_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1955_3_lut_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__34884),
            .in2(N__37608),
            .in3(N__34851),
            .lcout(\nx.n2896 ),
            .ltout(\nx.n2896_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_115_LC_14_18_5 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_115_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_115_LC_14_18_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_115_LC_14_18_5  (
            .in0(N__35151),
            .in1(N__35369),
            .in2(N__34836),
            .in3(N__35105),
            .lcout(),
            .ltout(\nx.n43_adj_763_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i22_4_lut_adj_123_LC_14_18_6 .C_ON=1'b0;
    defparam \nx.i22_4_lut_adj_123_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \nx.i22_4_lut_adj_123_LC_14_18_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i22_4_lut_adj_123_LC_14_18_6  (
            .in0(N__36803),
            .in1(N__35027),
            .in2(N__34833),
            .in3(N__34830),
            .lcout(\nx.n47_adj_770 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1964_3_lut_LC_14_18_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1964_3_lut_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1964_3_lut_LC_14_18_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1964_3_lut_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__34818),
            .in2(N__34785),
            .in3(N__37598),
            .lcout(\nx.n2905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_2_lut_LC_14_19_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_2_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_2_lut_LC_14_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_2_lut_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__35258),
            .in2(_gnd_net_),
            .in3(N__35193),
            .lcout(\nx.n2977 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\nx.n11028 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_3_lut_LC_14_19_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_3_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_3_lut_LC_14_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_3_lut_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35190),
            .in3(N__35154),
            .lcout(\nx.n2976 ),
            .ltout(),
            .carryin(\nx.n11028 ),
            .carryout(\nx.n11029 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_4_lut_LC_14_19_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_4_lut_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_4_lut_LC_14_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_4_lut_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__41316),
            .in2(N__35146),
            .in3(N__35109),
            .lcout(\nx.n2975 ),
            .ltout(),
            .carryin(\nx.n11029 ),
            .carryout(\nx.n11030 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_5_lut_LC_14_19_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_5_lut_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_5_lut_LC_14_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_5_lut_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__41322),
            .in2(N__35099),
            .in3(N__35073),
            .lcout(\nx.n2974 ),
            .ltout(),
            .carryin(\nx.n11030 ),
            .carryout(\nx.n11031 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_6_lut_LC_14_19_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_6_lut_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_6_lut_LC_14_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_6_lut_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__41317),
            .in2(N__35070),
            .in3(N__35031),
            .lcout(\nx.n2973 ),
            .ltout(),
            .carryin(\nx.n11031 ),
            .carryout(\nx.n11032 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_7_lut_LC_14_19_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_7_lut_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_7_lut_LC_14_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_7_lut_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__35026),
            .in2(N__41639),
            .in3(N__35004),
            .lcout(\nx.n2972 ),
            .ltout(),
            .carryin(\nx.n11032 ),
            .carryout(\nx.n11033 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_8_lut_LC_14_19_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_8_lut_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_8_lut_LC_14_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_8_lut_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__41321),
            .in2(N__37418),
            .in3(N__34989),
            .lcout(\nx.n2971 ),
            .ltout(),
            .carryin(\nx.n11033 ),
            .carryout(\nx.n11034 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_9_lut_LC_14_19_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_9_lut_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_9_lut_LC_14_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_9_lut_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__41323),
            .in2(N__36802),
            .in3(N__34986),
            .lcout(\nx.n2970 ),
            .ltout(),
            .carryin(\nx.n11034 ),
            .carryout(\nx.n11035 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_10_lut_LC_14_20_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_10_lut_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_10_lut_LC_14_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_10_lut_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__41640),
            .in2(N__35516),
            .in3(N__35466),
            .lcout(\nx.n2969 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\nx.n11036 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_11_lut_LC_14_20_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_11_lut_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_11_lut_LC_14_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_11_lut_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__41644),
            .in2(N__35463),
            .in3(N__35415),
            .lcout(\nx.n2968 ),
            .ltout(),
            .carryin(\nx.n11036 ),
            .carryout(\nx.n11037 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_12_lut_LC_14_20_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_12_lut_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_12_lut_LC_14_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_12_lut_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__41641),
            .in2(N__35411),
            .in3(N__35373),
            .lcout(\nx.n2967 ),
            .ltout(),
            .carryin(\nx.n11037 ),
            .carryout(\nx.n11038 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_13_lut_LC_14_20_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_13_lut_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_13_lut_LC_14_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_13_lut_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__41645),
            .in2(N__35370),
            .in3(N__35322),
            .lcout(\nx.n2966 ),
            .ltout(),
            .carryin(\nx.n11038 ),
            .carryout(\nx.n11039 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_14_lut_LC_14_20_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_14_lut_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_14_lut_LC_14_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_14_lut_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__41642),
            .in2(N__37437),
            .in3(N__35310),
            .lcout(\nx.n2965 ),
            .ltout(),
            .carryin(\nx.n11039 ),
            .carryout(\nx.n11040 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_15_lut_LC_14_20_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_15_lut_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_15_lut_LC_14_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_15_lut_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__41646),
            .in2(N__37381),
            .in3(N__35295),
            .lcout(\nx.n2964 ),
            .ltout(),
            .carryin(\nx.n11040 ),
            .carryout(\nx.n11041 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_16_lut_LC_14_20_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_16_lut_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_16_lut_LC_14_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_16_lut_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__41643),
            .in2(N__37011),
            .in3(N__35292),
            .lcout(\nx.n2963 ),
            .ltout(),
            .carryin(\nx.n11041 ),
            .carryout(\nx.n11042 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_17_lut_LC_14_20_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_17_lut_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_17_lut_LC_14_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_17_lut_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__41647),
            .in2(N__35289),
            .in3(N__35262),
            .lcout(\nx.n2962 ),
            .ltout(),
            .carryin(\nx.n11042 ),
            .carryout(\nx.n11043 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_18_lut_LC_14_21_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_18_lut_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_18_lut_LC_14_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_18_lut_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__41648),
            .in2(N__37353),
            .in3(N__35691),
            .lcout(\nx.n2961 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\nx.n11044 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_19_lut_LC_14_21_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_19_lut_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_19_lut_LC_14_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_19_lut_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__37448),
            .in2(N__41997),
            .in3(N__35688),
            .lcout(\nx.n2960 ),
            .ltout(),
            .carryin(\nx.n11044 ),
            .carryout(\nx.n11045 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_20_lut_LC_14_21_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_20_lut_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_20_lut_LC_14_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_20_lut_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__41652),
            .in2(N__37718),
            .in3(N__35679),
            .lcout(\nx.n2959 ),
            .ltout(),
            .carryin(\nx.n11045 ),
            .carryout(\nx.n11046 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_21_lut_LC_14_21_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_21_lut_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_21_lut_LC_14_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_21_lut_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__41655),
            .in2(N__36915),
            .in3(N__35676),
            .lcout(\nx.n2958 ),
            .ltout(),
            .carryin(\nx.n11046 ),
            .carryout(\nx.n11047 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_22_lut_LC_14_21_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_22_lut_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_22_lut_LC_14_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_22_lut_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__41653),
            .in2(N__37107),
            .in3(N__35661),
            .lcout(\nx.n2957 ),
            .ltout(),
            .carryin(\nx.n11047 ),
            .carryout(\nx.n11048 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_23_lut_LC_14_21_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_23_lut_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_23_lut_LC_14_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_23_lut_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__41656),
            .in2(N__35658),
            .in3(N__35625),
            .lcout(\nx.n2956 ),
            .ltout(),
            .carryin(\nx.n11048 ),
            .carryout(\nx.n11049 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_24_lut_LC_14_21_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_24_lut_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_24_lut_LC_14_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_24_lut_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__41654),
            .in2(N__35622),
            .in3(N__35574),
            .lcout(\nx.n2955 ),
            .ltout(),
            .carryin(\nx.n11049 ),
            .carryout(\nx.n11050 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_25_lut_LC_14_21_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_25_lut_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_25_lut_LC_14_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_25_lut_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__41657),
            .in2(N__35571),
            .in3(N__35538),
            .lcout(\nx.n2954 ),
            .ltout(),
            .carryin(\nx.n11050 ),
            .carryout(\nx.n11051 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_26_lut_LC_14_22_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_2009_26_lut_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_26_lut_LC_14_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_2009_26_lut_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(N__41679),
            .in2(N__35535),
            .in3(N__35874),
            .lcout(\nx.n2953 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\nx.n11052 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_2009_27_lut_LC_14_22_1 .C_ON=1'b0;
    defparam \nx.mod_5_add_2009_27_lut_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_2009_27_lut_LC_14_22_1 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_2009_27_lut_LC_14_22_1  (
            .in0(N__41680),
            .in1(N__37263),
            .in2(N__35871),
            .in3(N__35847),
            .lcout(\nx.n2984 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_adj_128_LC_14_22_4 .C_ON=1'b0;
    defparam \nx.i18_4_lut_adj_128_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_adj_128_LC_14_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_adj_128_LC_14_22_4  (
            .in0(N__35817),
            .in1(N__35811),
            .in2(N__40203),
            .in3(N__40373),
            .lcout(\nx.n39_adj_773 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_42_LC_14_22_5 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_42_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_42_LC_14_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_42_LC_14_22_5  (
            .in0(N__35804),
            .in1(N__35764),
            .in2(N__37846),
            .in3(N__37804),
            .lcout(\nx.n39_adj_689 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1754_rep_17_3_lut_LC_14_22_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1754_rep_17_3_lut_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1754_rep_17_3_lut_LC_14_22_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1754_rep_17_3_lut_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(N__40241),
            .in2(N__40221),
            .in3(N__40902),
            .lcout(\nx.n2599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_60_LC_14_23_0 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_60_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_60_LC_14_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_60_LC_14_23_0  (
            .in0(N__38104),
            .in1(N__38254),
            .in2(N__36131),
            .in3(N__38173),
            .lcout(\nx.n32_adj_703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i5_3_lut_adj_59_LC_14_23_1 .C_ON=1'b0;
    defparam \nx.i5_3_lut_adj_59_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.i5_3_lut_adj_59_LC_14_23_1 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \nx.i5_3_lut_adj_59_LC_14_23_1  (
            .in0(N__36058),
            .in1(_gnd_net_),
            .in2(N__35970),
            .in3(N__38317),
            .lcout(),
            .ltout(\nx.n25_adj_702_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i17_4_lut_adj_64_LC_14_23_2 .C_ON=1'b0;
    defparam \nx.i17_4_lut_adj_64_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.i17_4_lut_adj_64_LC_14_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i17_4_lut_adj_64_LC_14_23_2  (
            .in0(N__38290),
            .in1(N__38143),
            .in2(N__35736),
            .in3(N__35733),
            .lcout(),
            .ltout(\nx.n37_adj_709_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i19_4_lut_adj_65_LC_14_23_3 .C_ON=1'b0;
    defparam \nx.i19_4_lut_adj_65_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.i19_4_lut_adj_65_LC_14_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i19_4_lut_adj_65_LC_14_23_3  (
            .in0(N__35721),
            .in1(N__35712),
            .in2(N__35706),
            .in3(N__35703),
            .lcout(\nx.n2423 ),
            .ltout(\nx.n2423_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1696_3_lut_LC_14_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1696_3_lut_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1696_3_lut_LC_14_23_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1696_3_lut_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(N__36059),
            .in2(N__36078),
            .in3(N__36015),
            .lcout(\nx.n2509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1693_3_lut_LC_14_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1693_3_lut_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1693_3_lut_LC_14_23_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1693_3_lut_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(N__35949),
            .in2(N__38498),
            .in3(N__35968),
            .lcout(\nx.n2506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1625_rep_29_3_lut_LC_14_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1625_rep_29_3_lut_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1625_rep_29_3_lut_LC_14_23_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1625_rep_29_3_lut_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__36075),
            .in2(N__35925),
            .in3(N__38465),
            .lcout(\nx.n13321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_2_lut_LC_14_24_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_2_lut_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_2_lut_LC_14_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_2_lut_LC_14_24_0  (
            .in0(_gnd_net_),
            .in1(N__36057),
            .in2(_gnd_net_),
            .in3(N__36009),
            .lcout(\nx.n2477 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\nx.n10918 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_3_lut_LC_14_24_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_3_lut_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_3_lut_LC_14_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_3_lut_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38321),
            .in3(N__36006),
            .lcout(\nx.n2476 ),
            .ltout(),
            .carryin(\nx.n10918 ),
            .carryout(\nx.n10919 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_4_lut_LC_14_24_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_4_lut_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_4_lut_LC_14_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_4_lut_LC_14_24_2  (
            .in0(_gnd_net_),
            .in1(N__42009),
            .in2(N__36002),
            .in3(N__35973),
            .lcout(\nx.n2475 ),
            .ltout(),
            .carryin(\nx.n10919 ),
            .carryout(\nx.n10920 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_5_lut_LC_14_24_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_5_lut_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_5_lut_LC_14_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_5_lut_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(N__42012),
            .in2(N__35969),
            .in3(N__35943),
            .lcout(\nx.n2474 ),
            .ltout(),
            .carryin(\nx.n10920 ),
            .carryout(\nx.n10921 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_6_lut_LC_14_24_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_6_lut_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_6_lut_LC_14_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_6_lut_LC_14_24_4  (
            .in0(_gnd_net_),
            .in1(N__42010),
            .in2(N__35940),
            .in3(N__35916),
            .lcout(\nx.n2473 ),
            .ltout(),
            .carryin(\nx.n10921 ),
            .carryout(\nx.n10922 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_7_lut_LC_14_24_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_7_lut_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_7_lut_LC_14_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_7_lut_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(N__42013),
            .in2(N__35912),
            .in3(N__36285),
            .lcout(\nx.n2472 ),
            .ltout(),
            .carryin(\nx.n10922 ),
            .carryout(\nx.n10923 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_8_lut_LC_14_24_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_8_lut_LC_14_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_8_lut_LC_14_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_8_lut_LC_14_24_6  (
            .in0(_gnd_net_),
            .in1(N__42011),
            .in2(N__36281),
            .in3(N__36252),
            .lcout(\nx.n2471 ),
            .ltout(),
            .carryin(\nx.n10923 ),
            .carryout(\nx.n10924 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_9_lut_LC_14_24_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_9_lut_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_9_lut_LC_14_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_9_lut_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(N__42014),
            .in2(N__36245),
            .in3(N__36216),
            .lcout(\nx.n2470 ),
            .ltout(),
            .carryin(\nx.n10924 ),
            .carryout(\nx.n10925 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_10_lut_LC_14_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_10_lut_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_10_lut_LC_14_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_10_lut_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(N__42000),
            .in2(N__36213),
            .in3(N__36177),
            .lcout(\nx.n2469 ),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(\nx.n10926 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_11_lut_LC_14_25_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_11_lut_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_11_lut_LC_14_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_11_lut_LC_14_25_1  (
            .in0(_gnd_net_),
            .in1(N__42021),
            .in2(N__36170),
            .in3(N__36138),
            .lcout(\nx.n2468 ),
            .ltout(),
            .carryin(\nx.n10926 ),
            .carryout(\nx.n10927 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_12_lut_LC_14_25_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_12_lut_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_12_lut_LC_14_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_12_lut_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(N__42001),
            .in2(N__38297),
            .in3(N__36135),
            .lcout(\nx.n2467 ),
            .ltout(),
            .carryin(\nx.n10927 ),
            .carryout(\nx.n10928 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_13_lut_LC_14_25_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_13_lut_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_13_lut_LC_14_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_13_lut_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(N__42022),
            .in2(N__36127),
            .in3(N__36087),
            .lcout(\nx.n2466 ),
            .ltout(),
            .carryin(\nx.n10928 ),
            .carryout(\nx.n10929 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_14_lut_LC_14_25_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_14_lut_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_14_lut_LC_14_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_14_lut_LC_14_25_4  (
            .in0(_gnd_net_),
            .in1(N__42002),
            .in2(N__38204),
            .in3(N__36084),
            .lcout(\nx.n2465 ),
            .ltout(),
            .carryin(\nx.n10929 ),
            .carryout(\nx.n10930 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_15_lut_LC_14_25_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_15_lut_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_15_lut_LC_14_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_15_lut_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__42023),
            .in2(N__38148),
            .in3(N__36081),
            .lcout(\nx.n2464 ),
            .ltout(),
            .carryin(\nx.n10930 ),
            .carryout(\nx.n10931 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_16_lut_LC_14_25_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_16_lut_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_16_lut_LC_14_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_16_lut_LC_14_25_6  (
            .in0(_gnd_net_),
            .in1(N__42003),
            .in2(N__38259),
            .in3(N__36381),
            .lcout(\nx.n2463 ),
            .ltout(),
            .carryin(\nx.n10931 ),
            .carryout(\nx.n10932 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_17_lut_LC_14_25_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_17_lut_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_17_lut_LC_14_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_17_lut_LC_14_25_7  (
            .in0(_gnd_net_),
            .in1(N__42024),
            .in2(N__38180),
            .in3(N__36378),
            .lcout(\nx.n2462 ),
            .ltout(),
            .carryin(\nx.n10932 ),
            .carryout(\nx.n10933 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_18_lut_LC_14_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_18_lut_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_18_lut_LC_14_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_18_lut_LC_14_26_0  (
            .in0(_gnd_net_),
            .in1(N__42004),
            .in2(N__38105),
            .in3(N__36375),
            .lcout(\nx.n2461 ),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(\nx.n10934 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_19_lut_LC_14_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_19_lut_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_19_lut_LC_14_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_19_lut_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(N__42032),
            .in2(N__38531),
            .in3(N__36372),
            .lcout(\nx.n2460 ),
            .ltout(),
            .carryin(\nx.n10934 ),
            .carryout(\nx.n10935 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_20_lut_LC_14_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_20_lut_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_20_lut_LC_14_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_20_lut_LC_14_26_2  (
            .in0(_gnd_net_),
            .in1(N__42005),
            .in2(N__38591),
            .in3(N__36369),
            .lcout(\nx.n2459 ),
            .ltout(),
            .carryin(\nx.n10935 ),
            .carryout(\nx.n10936 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_21_lut_LC_14_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1674_21_lut_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_21_lut_LC_14_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1674_21_lut_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(N__38054),
            .in2(N__42209),
            .in3(N__36366),
            .lcout(\nx.n2458 ),
            .ltout(),
            .carryin(\nx.n10936 ),
            .carryout(\nx.n10937 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1674_22_lut_LC_14_26_4 .C_ON=1'b0;
    defparam \nx.mod_5_add_1674_22_lut_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1674_22_lut_LC_14_26_4 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_1674_22_lut_LC_14_26_4  (
            .in0(N__42033),
            .in1(N__38500),
            .in2(N__36363),
            .in3(N__36342),
            .lcout(\nx.n2489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i18_LC_14_26_6.C_ON=1'b0;
    defparam pin_output_enable__i18_LC_14_26_6.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i18_LC_14_26_6.LUT_INIT=16'b1101100011001100;
    LogicCell40 pin_output_enable__i18_LC_14_26_6 (
            .in0(N__38964),
            .in1(N__36329),
            .in2(N__47694),
            .in3(N__47154),
            .lcout(pin_oe_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46917),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1613_3_lut_LC_14_27_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1613_3_lut_LC_14_27_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1613_3_lut_LC_14_27_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1613_3_lut_LC_14_27_2  (
            .in0(_gnd_net_),
            .in1(N__36317),
            .in2(N__36294),
            .in3(N__38011),
            .lcout(\nx.n2394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1615_3_lut_LC_14_27_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1615_3_lut_LC_14_27_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1615_3_lut_LC_14_27_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1615_3_lut_LC_14_27_4  (
            .in0(_gnd_net_),
            .in1(N__36672),
            .in2(N__36648),
            .in3(N__38012),
            .lcout(\nx.n2396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1616_3_lut_LC_14_27_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1616_3_lut_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1616_3_lut_LC_14_27_5 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \nx.mod_5_i1616_3_lut_LC_14_27_5  (
            .in0(N__38014),
            .in1(N__36639),
            .in2(N__36615),
            .in3(_gnd_net_),
            .lcout(\nx.n2397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1483_3_lut_LC_14_27_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1483_3_lut_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1483_3_lut_LC_14_27_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1483_3_lut_LC_14_27_6  (
            .in0(_gnd_net_),
            .in1(N__36606),
            .in2(N__36594),
            .in3(N__36562),
            .lcout(\nx.n2200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1619_3_lut_LC_14_27_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1619_3_lut_LC_14_27_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1619_3_lut_LC_14_27_7 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \nx.mod_5_i1619_3_lut_LC_14_27_7  (
            .in0(N__38013),
            .in1(N__36423),
            .in2(N__36396),
            .in3(_gnd_net_),
            .lcout(\nx.n2400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam state__i0_LC_15_14_4.C_ON=1'b0;
    defparam state__i0_LC_15_14_4.SEQ_MODE=4'b1000;
    defparam state__i0_LC_15_14_4.LUT_INIT=16'b0011000000110011;
    LogicCell40 state__i0_LC_15_14_4 (
            .in0(_gnd_net_),
            .in1(N__47325),
            .in2(N__43191),
            .in3(N__43822),
            .lcout(state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46893),
            .ce(N__42399),
            .sr(N__38390));
    defparam state__i2_LC_15_14_5.C_ON=1'b0;
    defparam state__i2_LC_15_14_5.SEQ_MODE=4'b1000;
    defparam state__i2_LC_15_14_5.LUT_INIT=16'b0001000100000000;
    LogicCell40 state__i2_LC_15_14_5 (
            .in0(N__47324),
            .in1(N__43186),
            .in2(_gnd_net_),
            .in3(N__43823),
            .lcout(state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46893),
            .ce(N__42399),
            .sr(N__38390));
    defparam i1_2_lut_LC_15_15_0.C_ON=1'b0;
    defparam i1_2_lut_LC_15_15_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_15_15_0.LUT_INIT=16'b1111111101010101;
    LogicCell40 i1_2_lut_LC_15_15_0 (
            .in0(N__43817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43584),
            .lcout(n7602),
            .ltout(n7602_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_195_LC_15_15_1.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_195_LC_15_15_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_195_LC_15_15_1.LUT_INIT=16'b1100110011000100;
    LogicCell40 i1_3_lut_4_lut_adj_195_LC_15_15_1 (
            .in0(N__36729),
            .in1(N__45902),
            .in2(N__36387),
            .in3(N__47299),
            .lcout(n7730),
            .ltout(n7730_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i9_LC_15_15_2.C_ON=1'b0;
    defparam pin_output_enable__i9_LC_15_15_2.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i9_LC_15_15_2.LUT_INIT=16'b1100110010101100;
    LogicCell40 pin_output_enable__i9_LC_15_15_2 (
            .in0(N__47301),
            .in1(N__36767),
            .in2(N__36384),
            .in3(N__42381),
            .lcout(pin_oe_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46888),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i10_LC_15_15_4.C_ON=1'b0;
    defparam pin_output_enable__i10_LC_15_15_4.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i10_LC_15_15_4.LUT_INIT=16'b1011100010101010;
    LogicCell40 pin_output_enable__i10_LC_15_15_4 (
            .in0(N__36746),
            .in1(N__36735),
            .in2(N__47431),
            .in3(N__47039),
            .lcout(pin_oe_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46888),
            .ce(),
            .sr(_gnd_net_));
    defparam i7623_2_lut_3_lut_4_lut_4_lut_LC_15_15_5.C_ON=1'b0;
    defparam i7623_2_lut_3_lut_4_lut_4_lut_LC_15_15_5.SEQ_MODE=4'b0000;
    defparam i7623_2_lut_3_lut_4_lut_4_lut_LC_15_15_5.LUT_INIT=16'b1100110011001000;
    LogicCell40 i7623_2_lut_3_lut_4_lut_4_lut_LC_15_15_5 (
            .in0(N__44430),
            .in1(N__47300),
            .in2(N__45681),
            .in3(N__44532),
            .lcout(n11960),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i308_2_lut_LC_15_16_2.C_ON=1'b0;
    defparam i308_2_lut_LC_15_16_2.SEQ_MODE=4'b0000;
    defparam i308_2_lut_LC_15_16_2.LUT_INIT=16'b1100110011111111;
    LogicCell40 i308_2_lut_LC_15_16_2 (
            .in0(_gnd_net_),
            .in1(N__38627),
            .in2(_gnd_net_),
            .in3(N__43184),
            .lcout(n2618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i3_LC_15_16_4.C_ON=1'b0;
    defparam pin_output_enable__i3_LC_15_16_4.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i3_LC_15_16_4.LUT_INIT=16'b1010001011100010;
    LogicCell40 pin_output_enable__i3_LC_15_16_4 (
            .in0(N__36713),
            .in1(N__47038),
            .in2(N__47577),
            .in3(N__38646),
            .lcout(pin_oe_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46885),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_164_LC_15_17_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_164_LC_15_17_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_164_LC_15_17_2.LUT_INIT=16'b1100110011001101;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_164_LC_15_17_2 (
            .in0(N__44968),
            .in1(N__44831),
            .in2(N__45664),
            .in3(N__44503),
            .lcout(),
            .ltout(n8_adj_825_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i9_LC_15_17_3.C_ON=1'b0;
    defparam pin_output_i0_i9_LC_15_17_3.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i9_LC_15_17_3.LUT_INIT=16'b0111111100100000;
    LogicCell40 pin_output_i0_i9_LC_15_17_3 (
            .in0(N__45898),
            .in1(N__46147),
            .in2(N__36702),
            .in3(N__36689),
            .lcout(pin_out_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46880),
            .ce(),
            .sr(_gnd_net_));
    defparam i9176_2_lut_3_lut_4_lut_3_lut_LC_15_17_4.C_ON=1'b0;
    defparam i9176_2_lut_3_lut_4_lut_3_lut_LC_15_17_4.SEQ_MODE=4'b0000;
    defparam i9176_2_lut_3_lut_4_lut_3_lut_LC_15_17_4.LUT_INIT=16'b0000000001100110;
    LogicCell40 i9176_2_lut_3_lut_4_lut_3_lut_LC_15_17_4 (
            .in0(N__43836),
            .in1(N__47367),
            .in2(_gnd_net_),
            .in3(N__43596),
            .lcout(n11789),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8974_3_lut_LC_15_18_1.C_ON=1'b0;
    defparam i8974_3_lut_LC_15_18_1.SEQ_MODE=4'b0000;
    defparam i8974_3_lut_LC_15_18_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i8974_3_lut_LC_15_18_1 (
            .in0(N__46385),
            .in1(N__36688),
            .in2(_gnd_net_),
            .in3(N__43340),
            .lcout(n13369),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_240_i6_2_lut_LC_15_18_4.C_ON=1'b0;
    defparam equal_240_i6_2_lut_LC_15_18_4.SEQ_MODE=4'b0000;
    defparam equal_240_i6_2_lut_LC_15_18_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 equal_240_i6_2_lut_LC_15_18_4 (
            .in0(_gnd_net_),
            .in1(N__46564),
            .in2(_gnd_net_),
            .in3(N__46386),
            .lcout(n6_adj_813),
            .ltout(n6_adj_813_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7637_2_lut_3_lut_4_lut_4_lut_LC_15_18_5.C_ON=1'b0;
    defparam i7637_2_lut_3_lut_4_lut_4_lut_LC_15_18_5.SEQ_MODE=4'b0000;
    defparam i7637_2_lut_3_lut_4_lut_4_lut_LC_15_18_5.LUT_INIT=16'b1100100011001100;
    LogicCell40 i7637_2_lut_3_lut_4_lut_4_lut_LC_15_18_5 (
            .in0(N__42578),
            .in1(N__47590),
            .in2(N__37122),
            .in3(N__45627),
            .lcout(n11974),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_adj_122_LC_15_19_2 .C_ON=1'b0;
    defparam \nx.i20_4_lut_adj_122_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_adj_122_LC_15_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i20_4_lut_adj_122_LC_15_19_2  (
            .in0(N__37714),
            .in1(N__37102),
            .in2(N__37065),
            .in3(N__37047),
            .lcout(),
            .ltout(\nx.n45_adj_769_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i24_4_lut_adj_124_LC_15_19_3 .C_ON=1'b0;
    defparam \nx.i24_4_lut_adj_124_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \nx.i24_4_lut_adj_124_LC_15_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i24_4_lut_adj_124_LC_15_19_3  (
            .in0(N__37359),
            .in1(N__37035),
            .in2(N__37020),
            .in3(N__37017),
            .lcout(\nx.n2918 ),
            .ltout(\nx.n2918_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2022_3_lut_LC_15_19_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2022_3_lut_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2022_3_lut_LC_15_19_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2022_3_lut_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__37007),
            .in2(N__36993),
            .in3(N__36990),
            .lcout(\nx.n2995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2029_3_lut_LC_15_19_6 .C_ON=1'b0;
    defparam \nx.mod_5_i2029_3_lut_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2029_3_lut_LC_15_19_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2029_3_lut_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__36984),
            .in2(N__36804),
            .in3(N__37262),
            .lcout(\nx.n3002 ),
            .ltout(\nx.n3002_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_LC_15_19_7 .C_ON=1'b0;
    defparam \nx.i16_4_lut_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_LC_15_19_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_LC_15_19_7  (
            .in0(N__36947),
            .in1(N__37159),
            .in2(N__36936),
            .in3(N__37673),
            .lcout(\nx.n42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2017_3_lut_LC_15_20_0 .C_ON=1'b0;
    defparam \nx.mod_5_i2017_3_lut_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2017_3_lut_LC_15_20_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i2017_3_lut_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__36921),
            .in2(N__36911),
            .in3(N__37227),
            .lcout(\nx.n2990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1962_3_lut_LC_15_20_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1962_3_lut_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1962_3_lut_LC_15_20_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1962_3_lut_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__36849),
            .in2(N__36822),
            .in3(N__37603),
            .lcout(\nx.n2903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1951_3_lut_LC_15_20_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1951_3_lut_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1951_3_lut_LC_15_20_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1951_3_lut_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__37773),
            .in2(N__37743),
            .in3(N__37605),
            .lcout(\nx.n2892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2019_3_lut_LC_15_20_4 .C_ON=1'b0;
    defparam \nx.mod_5_i2019_3_lut_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2019_3_lut_LC_15_20_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i2019_3_lut_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__37449),
            .in2(N__37695),
            .in3(N__37231),
            .lcout(\nx.n2992 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1952_3_lut_LC_15_20_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1952_3_lut_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1952_3_lut_LC_15_20_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1952_3_lut_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(N__37662),
            .in2(N__37626),
            .in3(N__37604),
            .lcout(\nx.n2893 ),
            .ltout(\nx.n2893_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_121_LC_15_20_6 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_121_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_121_LC_15_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_121_LC_15_20_6  (
            .in0(N__37436),
            .in1(N__37419),
            .in2(N__37395),
            .in3(N__37382),
            .lcout(\nx.n41_adj_768 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i2020_3_lut_LC_15_20_7 .C_ON=1'b0;
    defparam \nx.mod_5_i2020_3_lut_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i2020_3_lut_LC_15_20_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i2020_3_lut_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(N__37349),
            .in2(N__37276),
            .in3(N__37173),
            .lcout(\nx.n2993 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i18_4_lut_LC_15_21_0 .C_ON=1'b0;
    defparam \nx.i18_4_lut_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.i18_4_lut_LC_15_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i18_4_lut_LC_15_21_0  (
            .in0(N__38821),
            .in1(N__39592),
            .in2(N__37131),
            .in3(N__38067),
            .lcout(\nx.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1764_3_lut_LC_15_21_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1764_3_lut_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1764_3_lut_LC_15_21_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \nx.mod_5_i1764_3_lut_LC_15_21_1  (
            .in0(N__39927),
            .in1(N__39864),
            .in2(_gnd_net_),
            .in3(N__40894),
            .lcout(\nx.n2609 ),
            .ltout(\nx.n2609_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i6_3_lut_adj_155_LC_15_21_2 .C_ON=1'b0;
    defparam \nx.i6_3_lut_adj_155_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.i6_3_lut_adj_155_LC_15_21_2 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \nx.i6_3_lut_adj_155_LC_15_21_2  (
            .in0(N__38927),
            .in1(_gnd_net_),
            .in2(N__37134),
            .in3(N__39643),
            .lcout(\nx.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1761_3_lut_LC_15_21_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1761_3_lut_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1761_3_lut_LC_15_21_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1761_3_lut_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__39747),
            .in2(N__39774),
            .in3(N__40898),
            .lcout(\nx.n2606 ),
            .ltout(\nx.n2606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1828_3_lut_LC_15_21_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1828_3_lut_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1828_3_lut_LC_15_21_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1828_3_lut_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__39351),
            .in2(N__37860),
            .in3(N__40101),
            .lcout(\nx.n2705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1763_3_lut_LC_15_21_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1763_3_lut_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1763_3_lut_LC_15_21_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1763_3_lut_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__39819),
            .in2(N__40921),
            .in3(N__39848),
            .lcout(\nx.n2608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1827_3_lut_LC_15_21_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1827_3_lut_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1827_3_lut_LC_15_21_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1827_3_lut_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__39337),
            .in2(N__40107),
            .in3(N__39315),
            .lcout(\nx.n2704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1762_3_lut_LC_15_22_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1762_3_lut_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1762_3_lut_LC_15_22_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1762_3_lut_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__39806),
            .in2(N__39789),
            .in3(N__40863),
            .lcout(\nx.n2607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i16_4_lut_adj_126_LC_15_22_1 .C_ON=1'b0;
    defparam \nx.i16_4_lut_adj_126_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.i16_4_lut_adj_126_LC_15_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i16_4_lut_adj_126_LC_15_22_1  (
            .in0(N__39805),
            .in1(N__40474),
            .in2(N__40446),
            .in3(N__38028),
            .lcout(),
            .ltout(\nx.n37_adj_772_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i20_4_lut_adj_141_LC_15_22_2 .C_ON=1'b0;
    defparam \nx.i20_4_lut_adj_141_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.i20_4_lut_adj_141_LC_15_22_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i20_4_lut_adj_141_LC_15_22_2  (
            .in0(N__38217),
            .in1(N__38550),
            .in2(N__37785),
            .in3(N__37782),
            .lcout(\nx.n2522 ),
            .ltout(\nx.n2522_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1760_3_lut_LC_15_22_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1760_3_lut_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1760_3_lut_LC_15_22_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \nx.mod_5_i1760_3_lut_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__40458),
            .in2(N__37776),
            .in3(N__40475),
            .lcout(\nx.n2605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1753_3_lut_LC_15_22_5 .C_ON=1'b0;
    defparam \nx.mod_5_i1753_3_lut_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1753_3_lut_LC_15_22_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1753_3_lut_LC_15_22_5  (
            .in0(N__40201),
            .in1(_gnd_net_),
            .in2(N__40900),
            .in3(N__40176),
            .lcout(\nx.n2598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1747_3_lut_LC_15_22_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1747_3_lut_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1747_3_lut_LC_15_22_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1747_3_lut_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__40864),
            .in2(N__40569),
            .in3(N__40542),
            .lcout(\nx.n2592 ),
            .ltout(\nx.n2592_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_LC_15_22_7 .C_ON=1'b0;
    defparam \nx.i13_4_lut_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_LC_15_22_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_LC_15_22_7  (
            .in0(N__38773),
            .in1(N__39538),
            .in2(N__38070),
            .in3(N__39487),
            .lcout(\nx.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1677_3_lut_LC_15_23_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1677_3_lut_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1677_3_lut_LC_15_23_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1677_3_lut_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__38061),
            .in2(N__38499),
            .in3(N__38040),
            .lcout(\nx.n2490 ),
            .ltout(\nx.n2490_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i1_2_lut_adj_108_LC_15_23_1 .C_ON=1'b0;
    defparam \nx.i1_2_lut_adj_108_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.i1_2_lut_adj_108_LC_15_23_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \nx.i1_2_lut_adj_108_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38031),
            .in3(N__40946),
            .lcout(\nx.n22_adj_755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1749_3_lut_LC_15_23_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1749_3_lut_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1749_3_lut_LC_15_23_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1749_3_lut_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__40637),
            .in2(N__40623),
            .in3(N__40861),
            .lcout(\nx.n2594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1748_3_lut_LC_15_23_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1748_3_lut_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1748_3_lut_LC_15_23_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \nx.mod_5_i1748_3_lut_LC_15_23_3  (
            .in0(N__40860),
            .in1(_gnd_net_),
            .in2(N__40584),
            .in3(N__40604),
            .lcout(\nx.n2593 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1751_3_lut_LC_15_23_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1751_3_lut_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1751_3_lut_LC_15_23_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1751_3_lut_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(N__40692),
            .in2(N__40674),
            .in3(N__40859),
            .lcout(\nx.n2596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i9121_3_lut_4_lut_LC_15_23_5 .C_ON=1'b0;
    defparam \nx.i9121_3_lut_4_lut_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.i9121_3_lut_4_lut_LC_15_23_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \nx.i9121_3_lut_4_lut_LC_15_23_5  (
            .in0(N__38022),
            .in1(N__38470),
            .in2(N__37905),
            .in3(N__37869),
            .lcout(\nx.n2505 ),
            .ltout(\nx.n2505_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1759_3_lut_LC_15_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1759_3_lut_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1759_3_lut_LC_15_23_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1759_3_lut_LC_15_23_6  (
            .in0(N__40428),
            .in1(_gnd_net_),
            .in2(N__37863),
            .in3(N__40862),
            .lcout(\nx.n2604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1695_3_lut_LC_15_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1695_3_lut_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1695_3_lut_LC_15_23_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1695_3_lut_LC_15_23_7  (
            .in0(N__38334),
            .in1(_gnd_net_),
            .in2(N__38328),
            .in3(N__38469),
            .lcout(\nx.n2508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1686_3_lut_LC_15_24_0 .C_ON=1'b0;
    defparam \nx.mod_5_i1686_3_lut_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1686_3_lut_LC_15_24_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1686_3_lut_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__38298),
            .in2(N__38268),
            .in3(N__38492),
            .lcout(\nx.n2499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1682_3_lut_LC_15_24_1 .C_ON=1'b0;
    defparam \nx.mod_5_i1682_3_lut_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1682_3_lut_LC_15_24_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \nx.mod_5_i1682_3_lut_LC_15_24_1  (
            .in0(N__38258),
            .in1(_gnd_net_),
            .in2(N__38505),
            .in3(N__38229),
            .lcout(\nx.n2495 ),
            .ltout(\nx.n2495_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i13_4_lut_adj_111_LC_15_24_2 .C_ON=1'b0;
    defparam \nx.i13_4_lut_adj_111_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.i13_4_lut_adj_111_LC_15_24_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i13_4_lut_adj_111_LC_15_24_2  (
            .in0(N__40658),
            .in1(N__40690),
            .in2(N__38220),
            .in3(N__40736),
            .lcout(\nx.n34_adj_758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1684_3_lut_LC_15_24_3 .C_ON=1'b0;
    defparam \nx.mod_5_i1684_3_lut_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1684_3_lut_LC_15_24_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \nx.mod_5_i1684_3_lut_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__38208),
            .in2(N__38504),
            .in3(N__38187),
            .lcout(\nx.n2497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1681_3_lut_LC_15_24_4 .C_ON=1'b0;
    defparam \nx.mod_5_i1681_3_lut_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1681_3_lut_LC_15_24_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1681_3_lut_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__38181),
            .in2(N__38157),
            .in3(N__38487),
            .lcout(\nx.n2494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1683_3_lut_LC_15_24_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1683_3_lut_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1683_3_lut_LC_15_24_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \nx.mod_5_i1683_3_lut_LC_15_24_6  (
            .in0(N__38147),
            .in1(_gnd_net_),
            .in2(N__38118),
            .in3(N__38488),
            .lcout(\nx.n2496 ),
            .ltout(\nx.n2496_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1750_3_lut_LC_15_24_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1750_3_lut_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1750_3_lut_LC_15_24_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \nx.mod_5_i1750_3_lut_LC_15_24_7  (
            .in0(N__40647),
            .in1(_gnd_net_),
            .in2(N__38109),
            .in3(N__40901),
            .lcout(\nx.n2595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1680_3_lut_LC_15_25_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1680_3_lut_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1680_3_lut_LC_15_25_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1680_3_lut_LC_15_25_2  (
            .in0(_gnd_net_),
            .in1(N__38106),
            .in2(N__38079),
            .in3(N__38502),
            .lcout(\nx.n2493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i22_LC_15_25_3.C_ON=1'b0;
    defparam pin_output_enable__i22_LC_15_25_3.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i22_LC_15_25_3.LUT_INIT=16'b1101000011001100;
    LogicCell40 pin_output_enable__i22_LC_15_25_3 (
            .in0(N__42663),
            .in1(N__38603),
            .in2(N__47695),
            .in3(N__47155),
            .lcout(pin_oe_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46918),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1678_3_lut_LC_15_25_6 .C_ON=1'b0;
    defparam \nx.mod_5_i1678_3_lut_LC_15_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1678_3_lut_LC_15_25_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \nx.mod_5_i1678_3_lut_LC_15_25_6  (
            .in0(_gnd_net_),
            .in1(N__38592),
            .in2(N__38562),
            .in3(N__38503),
            .lcout(\nx.n2491 ),
            .ltout(\nx.n2491_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.i12_4_lut_adj_120_LC_15_25_7 .C_ON=1'b0;
    defparam \nx.i12_4_lut_adj_120_LC_15_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.i12_4_lut_adj_120_LC_15_25_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \nx.i12_4_lut_adj_120_LC_15_25_7  (
            .in0(N__40516),
            .in1(N__40600),
            .in2(N__38553),
            .in3(N__40558),
            .lcout(\nx.n33_adj_767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1679_3_lut_LC_15_26_2 .C_ON=1'b0;
    defparam \nx.mod_5_i1679_3_lut_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1679_3_lut_LC_15_26_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \nx.mod_5_i1679_3_lut_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(N__38541),
            .in2(N__38535),
            .in3(N__38501),
            .lcout(\nx.n2492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1745_3_lut_LC_15_26_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1745_3_lut_LC_15_26_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1745_3_lut_LC_15_26_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1745_3_lut_LC_15_26_7  (
            .in0(_gnd_net_),
            .in1(N__40926),
            .in2(N__42363),
            .in3(N__42345),
            .lcout(\nx.n2590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam state__i1_LC_16_14_5.C_ON=1'b0;
    defparam state__i1_LC_16_14_5.SEQ_MODE=4'b1000;
    defparam state__i1_LC_16_14_5.LUT_INIT=16'b0100101000001010;
    LogicCell40 state__i1_LC_16_14_5 (
            .in0(N__47323),
            .in1(N__38631),
            .in2(N__43875),
            .in3(N__43190),
            .lcout(state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46897),
            .ce(N__42398),
            .sr(N__38391));
    defparam counter_633__i0_LC_16_15_5.C_ON=1'b0;
    defparam counter_633__i0_LC_16_15_5.SEQ_MODE=4'b1000;
    defparam counter_633__i0_LC_16_15_5.LUT_INIT=16'b1111111000000100;
    LogicCell40 counter_633__i0_LC_16_15_5 (
            .in0(N__38370),
            .in1(N__40758),
            .in2(N__47459),
            .in3(N__42888),
            .lcout(counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46894),
            .ce(N__45961),
            .sr(_gnd_net_));
    defparam pin_output_enable__i11_LC_16_16_0.C_ON=1'b0;
    defparam pin_output_enable__i11_LC_16_16_0.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i11_LC_16_16_0.LUT_INIT=16'b1100010011100100;
    LogicCell40 pin_output_enable__i11_LC_16_16_0 (
            .in0(N__47037),
            .in1(N__38345),
            .in2(N__47489),
            .in3(N__44219),
            .lcout(pin_oe_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46889),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_243_i6_2_lut_LC_16_16_4.C_ON=1'b0;
    defparam equal_243_i6_2_lut_LC_16_16_4.SEQ_MODE=4'b0000;
    defparam equal_243_i6_2_lut_LC_16_16_4.LUT_INIT=16'b1100110011111111;
    LogicCell40 equal_243_i6_2_lut_LC_16_16_4 (
            .in0(_gnd_net_),
            .in1(N__46509),
            .in2(_gnd_net_),
            .in3(N__46321),
            .lcout(n6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_197_LC_16_16_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_197_LC_16_16_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_197_LC_16_16_5.LUT_INIT=16'b0000000011101111;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_197_LC_16_16_5 (
            .in0(N__43600),
            .in1(N__47368),
            .in2(N__43890),
            .in3(N__42887),
            .lcout(n6_adj_819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_244_i7_2_lut_LC_16_17_0.C_ON=1'b0;
    defparam equal_244_i7_2_lut_LC_16_17_0.SEQ_MODE=4'b0000;
    defparam equal_244_i7_2_lut_LC_16_17_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 equal_244_i7_2_lut_LC_16_17_0 (
            .in0(_gnd_net_),
            .in1(N__43240),
            .in2(_gnd_net_),
            .in3(N__45263),
            .lcout(n7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_241_i9_2_lut_3_lut_4_lut_LC_16_17_1.C_ON=1'b0;
    defparam equal_241_i9_2_lut_3_lut_4_lut_LC_16_17_1.SEQ_MODE=4'b0000;
    defparam equal_241_i9_2_lut_3_lut_4_lut_LC_16_17_1.LUT_INIT=16'b1111111111111011;
    LogicCell40 equal_241_i9_2_lut_3_lut_4_lut_LC_16_17_1 (
            .in0(N__43241),
            .in1(N__43398),
            .in2(N__45270),
            .in3(N__45481),
            .lcout(n9),
            .ltout(n9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_193_LC_16_17_2.C_ON=1'b0;
    defparam i1_2_lut_adj_193_LC_16_17_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_193_LC_16_17_2.LUT_INIT=16'b1111111100001111;
    LogicCell40 i1_2_lut_adj_193_LC_16_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38640),
            .in3(N__44830),
            .lcout(),
            .ltout(n8_adj_820_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i3_LC_16_17_3.C_ON=1'b0;
    defparam pin_output_i0_i3_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i3_LC_16_17_3.LUT_INIT=16'b0111111100100000;
    LogicCell40 pin_output_i0_i3_LC_16_17_3 (
            .in0(N__45899),
            .in1(N__46145),
            .in2(N__38637),
            .in3(N__38707),
            .lcout(pin_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46884),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_180_LC_16_17_5.C_ON=1'b0;
    defparam i2_2_lut_adj_180_LC_16_17_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_180_LC_16_17_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i2_2_lut_adj_180_LC_16_17_5 (
            .in0(_gnd_net_),
            .in1(N__42494),
            .in2(_gnd_net_),
            .in3(N__42509),
            .lcout(),
            .ltout(n6_adj_805_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_181_LC_16_17_6.C_ON=1'b0;
    defparam i3_4_lut_adj_181_LC_16_17_6.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_181_LC_16_17_6.LUT_INIT=16'b1111111011111010;
    LogicCell40 i3_4_lut_adj_181_LC_16_17_6 (
            .in0(N__42476),
            .in1(N__43239),
            .in2(N__38634),
            .in3(N__45262),
            .lcout(n1788),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i4_LC_16_17_7.C_ON=1'b0;
    defparam pin_output_i0_i4_LC_16_17_7.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i4_LC_16_17_7.LUT_INIT=16'b0111111100100000;
    LogicCell40 pin_output_i0_i4_LC_16_17_7 (
            .in0(N__45900),
            .in1(N__46146),
            .in2(N__38730),
            .in3(N__42694),
            .lcout(pin_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46884),
            .ce(),
            .sr(_gnd_net_));
    defparam i5698_2_lut_LC_16_18_1.C_ON=1'b0;
    defparam i5698_2_lut_LC_16_18_1.SEQ_MODE=4'b0000;
    defparam i5698_2_lut_LC_16_18_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i5698_2_lut_LC_16_18_1 (
            .in0(_gnd_net_),
            .in1(N__46322),
            .in2(_gnd_net_),
            .in3(N__46508),
            .lcout(n9488),
            .ltout(n9488_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_233_i9_2_lut_3_lut_4_lut_LC_16_18_2.C_ON=1'b0;
    defparam equal_233_i9_2_lut_3_lut_4_lut_LC_16_18_2.SEQ_MODE=4'b0000;
    defparam equal_233_i9_2_lut_3_lut_4_lut_LC_16_18_2.LUT_INIT=16'b1111111111011111;
    LogicCell40 equal_233_i9_2_lut_3_lut_4_lut_LC_16_18_2 (
            .in0(N__45254),
            .in1(N__43242),
            .in2(N__38736),
            .in3(N__45454),
            .lcout(n9_adj_812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_234_i7_2_lut_LC_16_18_3.C_ON=1'b0;
    defparam equal_234_i7_2_lut_LC_16_18_3.SEQ_MODE=4'b0000;
    defparam equal_234_i7_2_lut_LC_16_18_3.LUT_INIT=16'b1010101011111111;
    LogicCell40 equal_234_i7_2_lut_LC_16_18_3 (
            .in0(N__43243),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45253),
            .lcout(n7_adj_811),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_172_LC_16_18_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_172_LC_16_18_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_172_LC_16_18_5.LUT_INIT=16'b1111111100000001;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_172_LC_16_18_5 (
            .in0(N__42583),
            .in1(N__44389),
            .in2(N__45568),
            .in3(N__44873),
            .lcout(),
            .ltout(n7_adj_818_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i2_LC_16_18_6.C_ON=1'b0;
    defparam pin_output_i0_i2_LC_16_18_6.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i2_LC_16_18_6.LUT_INIT=16'b0111111100100000;
    LogicCell40 pin_output_i0_i2_LC_16_18_6 (
            .in0(N__45901),
            .in1(N__46142),
            .in2(N__38733),
            .in3(N__38672),
            .lcout(pin_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46890),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_166_LC_16_18_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_166_LC_16_18_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_166_LC_16_18_7.LUT_INIT=16'b1111111100010000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_166_LC_16_18_7 (
            .in0(N__42582),
            .in1(N__44063),
            .in2(N__45567),
            .in3(N__44872),
            .lcout(n7_adj_821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_173_LC_16_19_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_173_LC_16_19_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_173_LC_16_19_2.LUT_INIT=16'b1111111100000001;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_173_LC_16_19_2 (
            .in0(N__42603),
            .in1(N__44990),
            .in2(N__45588),
            .in3(N__44874),
            .lcout(n8_adj_817),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8960_3_lut_LC_16_19_5.C_ON=1'b0;
    defparam i8960_3_lut_LC_16_19_5.SEQ_MODE=4'b0000;
    defparam i8960_3_lut_LC_16_19_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 i8960_3_lut_LC_16_19_5 (
            .in0(N__38711),
            .in1(N__38671),
            .in2(_gnd_net_),
            .in3(N__46384),
            .lcout(),
            .ltout(n13355_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13625_bdd_4_lut_LC_16_19_6.C_ON=1'b0;
    defparam n13625_bdd_4_lut_LC_16_19_6.SEQ_MODE=4'b0000;
    defparam n13625_bdd_4_lut_LC_16_19_6.LUT_INIT=16'b1111101001000100;
    LogicCell40 n13625_bdd_4_lut_LC_16_19_6 (
            .in0(N__45493),
            .in1(N__38652),
            .in2(N__38655),
            .in3(N__42672),
            .lcout(n13628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8959_3_lut_LC_16_20_0.C_ON=1'b0;
    defparam i8959_3_lut_LC_16_20_0.SEQ_MODE=4'b0000;
    defparam i8959_3_lut_LC_16_20_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i8959_3_lut_LC_16_20_0 (
            .in0(N__38977),
            .in1(N__39019),
            .in2(_gnd_net_),
            .in3(N__46383),
            .lcout(n13354),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_174_LC_16_20_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_174_LC_16_20_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_174_LC_16_20_1.LUT_INIT=16'b1111000011110001;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_174_LC_16_20_1 (
            .in0(N__44091),
            .in1(N__45498),
            .in2(N__44913),
            .in3(N__42604),
            .lcout(),
            .ltout(n7_adj_840_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i0_LC_16_20_2.C_ON=1'b0;
    defparam pin_output_i0_i0_LC_16_20_2.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i0_LC_16_20_2.LUT_INIT=16'b0011101010101010;
    LogicCell40 pin_output_i0_i0_LC_16_20_2 (
            .in0(N__39020),
            .in1(N__46143),
            .in2(N__39039),
            .in3(N__45973),
            .lcout(pin_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46898),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i1_LC_16_20_4.C_ON=1'b0;
    defparam pin_output_i0_i1_LC_16_20_4.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i1_LC_16_20_4.LUT_INIT=16'b0010111010101010;
    LogicCell40 pin_output_i0_i1_LC_16_20_4 (
            .in0(N__38978),
            .in1(N__39003),
            .in2(N__46152),
            .in3(N__45972),
            .lcout(pin_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46898),
            .ce(),
            .sr(_gnd_net_));
    defparam i7615_2_lut_3_lut_4_lut_4_lut_LC_16_20_6.C_ON=1'b0;
    defparam i7615_2_lut_3_lut_4_lut_4_lut_LC_16_20_6.SEQ_MODE=4'b0000;
    defparam i7615_2_lut_3_lut_4_lut_4_lut_LC_16_20_6.LUT_INIT=16'b1111000011100000;
    LogicCell40 i7615_2_lut_3_lut_4_lut_4_lut_LC_16_20_6 (
            .in0(N__45497),
            .in1(N__44387),
            .in2(N__47599),
            .in3(N__45107),
            .lcout(n11952),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i8_LC_16_20_7.C_ON=1'b0;
    defparam pin_output_enable__i8_LC_16_20_7.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i8_LC_16_20_7.LUT_INIT=16'b1010110010101010;
    LogicCell40 pin_output_enable__i8_LC_16_20_7 (
            .in0(N__38942),
            .in1(N__47502),
            .in2(N__42648),
            .in3(N__47156),
            .lcout(pin_oe_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46898),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_2_lut_LC_16_21_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_2_lut_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_2_lut_LC_16_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_2_lut_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__38931),
            .in2(_gnd_net_),
            .in3(N__38868),
            .lcout(\nx.n2677 ),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(\nx.n10959 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_3_lut_LC_16_21_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_3_lut_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_3_lut_LC_16_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_3_lut_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38861),
            .in3(N__38832),
            .lcout(\nx.n2676 ),
            .ltout(),
            .carryin(\nx.n10959 ),
            .carryout(\nx.n10960 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_4_lut_LC_16_21_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_4_lut_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_4_lut_LC_16_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_4_lut_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__42123),
            .in2(N__38825),
            .in3(N__38787),
            .lcout(\nx.n2675 ),
            .ltout(),
            .carryin(\nx.n10960 ),
            .carryout(\nx.n10961 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_5_lut_LC_16_21_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_5_lut_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_5_lut_LC_16_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_5_lut_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__42126),
            .in2(N__38780),
            .in3(N__38739),
            .lcout(\nx.n2674 ),
            .ltout(),
            .carryin(\nx.n10961 ),
            .carryout(\nx.n10962 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_6_lut_LC_16_21_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_6_lut_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_6_lut_LC_16_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_6_lut_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__42124),
            .in2(N__39368),
            .in3(N__39345),
            .lcout(\nx.n2673 ),
            .ltout(),
            .carryin(\nx.n10962 ),
            .carryout(\nx.n10963 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_7_lut_LC_16_21_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_7_lut_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_7_lut_LC_16_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_7_lut_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(N__42127),
            .in2(N__39338),
            .in3(N__39309),
            .lcout(\nx.n2672 ),
            .ltout(),
            .carryin(\nx.n10963 ),
            .carryout(\nx.n10964 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_8_lut_LC_16_21_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_8_lut_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_8_lut_LC_16_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_8_lut_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(N__42125),
            .in2(N__39305),
            .in3(N__39261),
            .lcout(\nx.n2671 ),
            .ltout(),
            .carryin(\nx.n10964 ),
            .carryout(\nx.n10965 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_9_lut_LC_16_21_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_9_lut_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_9_lut_LC_16_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_9_lut_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(N__42128),
            .in2(N__39258),
            .in3(N__39225),
            .lcout(\nx.n2670 ),
            .ltout(),
            .carryin(\nx.n10965 ),
            .carryout(\nx.n10966 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_10_lut_LC_16_22_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_10_lut_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_10_lut_LC_16_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_10_lut_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__42138),
            .in2(N__39222),
            .in3(N__39180),
            .lcout(\nx.n2669 ),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(\nx.n10967 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_11_lut_LC_16_22_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_11_lut_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_11_lut_LC_16_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_11_lut_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(N__42168),
            .in2(N__39177),
            .in3(N__39141),
            .lcout(\nx.n2668 ),
            .ltout(),
            .carryin(\nx.n10967 ),
            .carryout(\nx.n10968 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_12_lut_LC_16_22_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_12_lut_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_12_lut_LC_16_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_12_lut_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(N__42139),
            .in2(N__39137),
            .in3(N__39090),
            .lcout(\nx.n2667 ),
            .ltout(),
            .carryin(\nx.n10968 ),
            .carryout(\nx.n10969 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_13_lut_LC_16_22_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_13_lut_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_13_lut_LC_16_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_13_lut_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__42169),
            .in2(N__39087),
            .in3(N__39042),
            .lcout(\nx.n2666 ),
            .ltout(),
            .carryin(\nx.n10969 ),
            .carryout(\nx.n10970 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_14_lut_LC_16_22_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_14_lut_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_14_lut_LC_16_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_14_lut_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(N__42140),
            .in2(N__39731),
            .in3(N__39690),
            .lcout(\nx.n2665 ),
            .ltout(),
            .carryin(\nx.n10970 ),
            .carryout(\nx.n10971 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_15_lut_LC_16_22_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_15_lut_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_15_lut_LC_16_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_15_lut_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(N__42170),
            .in2(N__39687),
            .in3(N__39651),
            .lcout(\nx.n2664 ),
            .ltout(),
            .carryin(\nx.n10971 ),
            .carryout(\nx.n10972 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_16_lut_LC_16_22_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_16_lut_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_16_lut_LC_16_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_16_lut_LC_16_22_6  (
            .in0(_gnd_net_),
            .in1(N__42141),
            .in2(N__39644),
            .in3(N__39603),
            .lcout(\nx.n2663 ),
            .ltout(),
            .carryin(\nx.n10972 ),
            .carryout(\nx.n10973 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_17_lut_LC_16_22_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_17_lut_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_17_lut_LC_16_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_17_lut_LC_16_22_7  (
            .in0(_gnd_net_),
            .in1(N__42171),
            .in2(N__39599),
            .in3(N__39552),
            .lcout(\nx.n2662 ),
            .ltout(),
            .carryin(\nx.n10973 ),
            .carryout(\nx.n10974 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_18_lut_LC_16_23_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_18_lut_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_18_lut_LC_16_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_18_lut_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(N__42041),
            .in2(N__39545),
            .in3(N__39504),
            .lcout(\nx.n2661 ),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(\nx.n10975 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_19_lut_LC_16_23_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_19_lut_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_19_lut_LC_16_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_19_lut_LC_16_23_1  (
            .in0(_gnd_net_),
            .in1(N__42172),
            .in2(N__39494),
            .in3(N__39456),
            .lcout(\nx.n2660 ),
            .ltout(),
            .carryin(\nx.n10975 ),
            .carryout(\nx.n10976 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_20_lut_LC_16_23_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_20_lut_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_20_lut_LC_16_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_20_lut_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(N__42042),
            .in2(N__39452),
            .in3(N__39417),
            .lcout(\nx.n2659 ),
            .ltout(),
            .carryin(\nx.n10976 ),
            .carryout(\nx.n10977 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_21_lut_LC_16_23_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_21_lut_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_21_lut_LC_16_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_21_lut_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(N__42173),
            .in2(N__39414),
            .in3(N__39375),
            .lcout(\nx.n2658 ),
            .ltout(),
            .carryin(\nx.n10977 ),
            .carryout(\nx.n10978 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_22_lut_LC_16_23_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_22_lut_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_22_lut_LC_16_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_22_lut_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(N__42043),
            .in2(N__40164),
            .in3(N__40122),
            .lcout(\nx.n2657 ),
            .ltout(),
            .carryin(\nx.n10978 ),
            .carryout(\nx.n10979 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_23_lut_LC_16_23_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1808_23_lut_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_23_lut_LC_16_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1808_23_lut_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(N__42174),
            .in2(N__39949),
            .in3(N__40110),
            .lcout(\nx.n2656 ),
            .ltout(),
            .carryin(\nx.n10979 ),
            .carryout(\nx.n10980 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1808_24_lut_LC_16_23_6 .C_ON=1'b0;
    defparam \nx.mod_5_add_1808_24_lut_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1808_24_lut_LC_16_23_6 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \nx.mod_5_add_1808_24_lut_LC_16_23_6  (
            .in0(N__42175),
            .in1(N__40095),
            .in2(N__40803),
            .in3(N__39987),
            .lcout(\nx.n2687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_i1744_3_lut_LC_16_23_7 .C_ON=1'b0;
    defparam \nx.mod_5_i1744_3_lut_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_i1744_3_lut_LC_16_23_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \nx.mod_5_i1744_3_lut_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(N__40899),
            .in2(N__42332),
            .in3(N__42312),
            .lcout(\nx.n2589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_2_lut_LC_16_24_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_2_lut_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_2_lut_LC_16_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_2_lut_LC_16_24_0  (
            .in0(_gnd_net_),
            .in1(N__39922),
            .in2(_gnd_net_),
            .in3(N__39852),
            .lcout(\nx.n2577 ),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(\nx.n10938 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_3_lut_LC_16_24_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_3_lut_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_3_lut_LC_16_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_3_lut_LC_16_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39849),
            .in3(N__39810),
            .lcout(\nx.n2576 ),
            .ltout(),
            .carryin(\nx.n10938 ),
            .carryout(\nx.n10939 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_4_lut_LC_16_24_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_4_lut_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_4_lut_LC_16_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_4_lut_LC_16_24_2  (
            .in0(_gnd_net_),
            .in1(N__42270),
            .in2(N__39807),
            .in3(N__39777),
            .lcout(\nx.n2575 ),
            .ltout(),
            .carryin(\nx.n10939 ),
            .carryout(\nx.n10940 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_5_lut_LC_16_24_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_5_lut_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_5_lut_LC_16_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_5_lut_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(N__39770),
            .in2(N__42297),
            .in3(N__39738),
            .lcout(\nx.n2574 ),
            .ltout(),
            .carryin(\nx.n10940 ),
            .carryout(\nx.n10941 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_6_lut_LC_16_24_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_6_lut_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_6_lut_LC_16_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_6_lut_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(N__42274),
            .in2(N__40482),
            .in3(N__40449),
            .lcout(\nx.n2573 ),
            .ltout(),
            .carryin(\nx.n10941 ),
            .carryout(\nx.n10942 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_7_lut_LC_16_24_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_7_lut_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_7_lut_LC_16_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_7_lut_LC_16_24_5  (
            .in0(_gnd_net_),
            .in1(N__42255),
            .in2(N__40445),
            .in3(N__40422),
            .lcout(\nx.n2572 ),
            .ltout(),
            .carryin(\nx.n10942 ),
            .carryout(\nx.n10943 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_8_lut_LC_16_24_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_8_lut_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_8_lut_LC_16_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_8_lut_LC_16_24_6  (
            .in0(_gnd_net_),
            .in1(N__42275),
            .in2(N__40419),
            .in3(N__40377),
            .lcout(\nx.n2571 ),
            .ltout(),
            .carryin(\nx.n10943 ),
            .carryout(\nx.n10944 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_9_lut_LC_16_24_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_9_lut_LC_16_24_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_9_lut_LC_16_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_9_lut_LC_16_24_7  (
            .in0(_gnd_net_),
            .in1(N__40372),
            .in2(N__42298),
            .in3(N__40332),
            .lcout(\nx.n2570 ),
            .ltout(),
            .carryin(\nx.n10944 ),
            .carryout(\nx.n10945 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_10_lut_LC_16_25_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_10_lut_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_10_lut_LC_16_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_10_lut_LC_16_25_0  (
            .in0(_gnd_net_),
            .in1(N__42256),
            .in2(N__40329),
            .in3(N__40290),
            .lcout(\nx.n2569 ),
            .ltout(),
            .carryin(bfn_16_25_0_),
            .carryout(\nx.n10946 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_11_lut_LC_16_25_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_11_lut_LC_16_25_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_11_lut_LC_16_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_11_lut_LC_16_25_1  (
            .in0(_gnd_net_),
            .in1(N__42262),
            .in2(N__40287),
            .in3(N__40251),
            .lcout(\nx.n2568 ),
            .ltout(),
            .carryin(\nx.n10946 ),
            .carryout(\nx.n10947 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_12_lut_LC_16_25_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_12_lut_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_12_lut_LC_16_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_12_lut_LC_16_25_2  (
            .in0(_gnd_net_),
            .in1(N__42257),
            .in2(N__40248),
            .in3(N__40206),
            .lcout(\nx.n2567 ),
            .ltout(),
            .carryin(\nx.n10947 ),
            .carryout(\nx.n10948 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_13_lut_LC_16_25_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_13_lut_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_13_lut_LC_16_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_13_lut_LC_16_25_3  (
            .in0(_gnd_net_),
            .in1(N__42263),
            .in2(N__40202),
            .in3(N__40167),
            .lcout(\nx.n2566 ),
            .ltout(),
            .carryin(\nx.n10948 ),
            .carryout(\nx.n10949 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_14_lut_LC_16_25_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_14_lut_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_14_lut_LC_16_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_14_lut_LC_16_25_4  (
            .in0(_gnd_net_),
            .in1(N__42258),
            .in2(N__40740),
            .in3(N__40695),
            .lcout(\nx.n2565 ),
            .ltout(),
            .carryin(\nx.n10949 ),
            .carryout(\nx.n10950 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_15_lut_LC_16_25_5 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_15_lut_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_15_lut_LC_16_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_15_lut_LC_16_25_5  (
            .in0(_gnd_net_),
            .in1(N__40691),
            .in2(N__42295),
            .in3(N__40662),
            .lcout(\nx.n2564 ),
            .ltout(),
            .carryin(\nx.n10950 ),
            .carryout(\nx.n10951 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_16_lut_LC_16_25_6 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_16_lut_LC_16_25_6 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_16_lut_LC_16_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_16_lut_LC_16_25_6  (
            .in0(_gnd_net_),
            .in1(N__40659),
            .in2(N__42296),
            .in3(N__40641),
            .lcout(\nx.n2563 ),
            .ltout(),
            .carryin(\nx.n10951 ),
            .carryout(\nx.n10952 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_17_lut_LC_16_25_7 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_17_lut_LC_16_25_7 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_17_lut_LC_16_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_17_lut_LC_16_25_7  (
            .in0(_gnd_net_),
            .in1(N__42267),
            .in2(N__40638),
            .in3(N__40611),
            .lcout(\nx.n2562 ),
            .ltout(),
            .carryin(\nx.n10952 ),
            .carryout(\nx.n10953 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_18_lut_LC_16_26_0 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_18_lut_LC_16_26_0 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_18_lut_LC_16_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_18_lut_LC_16_26_0  (
            .in0(_gnd_net_),
            .in1(N__42251),
            .in2(N__40608),
            .in3(N__40572),
            .lcout(\nx.n2561 ),
            .ltout(),
            .carryin(bfn_16_26_0_),
            .carryout(\nx.n10954 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_19_lut_LC_16_26_1 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_19_lut_LC_16_26_1 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_19_lut_LC_16_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_19_lut_LC_16_26_1  (
            .in0(_gnd_net_),
            .in1(N__42268),
            .in2(N__40565),
            .in3(N__40530),
            .lcout(\nx.n2560 ),
            .ltout(),
            .carryin(\nx.n10954 ),
            .carryout(\nx.n10955 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_20_lut_LC_16_26_2 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_20_lut_LC_16_26_2 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_20_lut_LC_16_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_20_lut_LC_16_26_2  (
            .in0(_gnd_net_),
            .in1(N__42252),
            .in2(N__40523),
            .in3(N__40485),
            .lcout(\nx.n2559 ),
            .ltout(),
            .carryin(\nx.n10955 ),
            .carryout(\nx.n10956 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_21_lut_LC_16_26_3 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_21_lut_LC_16_26_3 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_21_lut_LC_16_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_21_lut_LC_16_26_3  (
            .in0(_gnd_net_),
            .in1(N__42269),
            .in2(N__42362),
            .in3(N__42339),
            .lcout(\nx.n2558 ),
            .ltout(),
            .carryin(\nx.n10956 ),
            .carryout(\nx.n10957 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_22_lut_LC_16_26_4 .C_ON=1'b1;
    defparam \nx.mod_5_add_1741_22_lut_LC_16_26_4 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_22_lut_LC_16_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \nx.mod_5_add_1741_22_lut_LC_16_26_4  (
            .in0(_gnd_net_),
            .in1(N__42253),
            .in2(N__42336),
            .in3(N__42303),
            .lcout(\nx.n2557 ),
            .ltout(),
            .carryin(\nx.n10957 ),
            .carryout(\nx.n10958 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \nx.mod_5_add_1741_23_lut_LC_16_26_5 .C_ON=1'b0;
    defparam \nx.mod_5_add_1741_23_lut_LC_16_26_5 .SEQ_MODE=4'b0000;
    defparam \nx.mod_5_add_1741_23_lut_LC_16_26_5 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \nx.mod_5_add_1741_23_lut_LC_16_26_5  (
            .in0(N__42254),
            .in1(N__40947),
            .in2(N__40929),
            .in3(N__40806),
            .lcout(\nx.n2588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9207_1_lut_2_lut_3_lut_LC_17_14_3.C_ON=1'b0;
    defparam i9207_1_lut_2_lut_3_lut_LC_17_14_3.SEQ_MODE=4'b0000;
    defparam i9207_1_lut_2_lut_3_lut_LC_17_14_3.LUT_INIT=16'b0000000000100010;
    LogicCell40 i9207_1_lut_2_lut_3_lut_LC_17_14_3 (
            .in0(N__43818),
            .in1(N__47363),
            .in2(_gnd_net_),
            .in3(N__43592),
            .lcout(n13603),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i12_LC_17_14_4.C_ON=1'b0;
    defparam pin_output_enable__i12_LC_17_14_4.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i12_LC_17_14_4.LUT_INIT=16'b1011100010101010;
    LogicCell40 pin_output_enable__i12_LC_17_14_4 (
            .in0(N__40769),
            .in1(N__42807),
            .in2(N__47488),
            .in3(N__47120),
            .lcout(pin_oe_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46902),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_633_add_4_2_lut_LC_17_15_0.C_ON=1'b1;
    defparam counter_633_add_4_2_lut_LC_17_15_0.SEQ_MODE=4'b0000;
    defparam counter_633_add_4_2_lut_LC_17_15_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_633_add_4_2_lut_LC_17_15_0 (
            .in0(_gnd_net_),
            .in1(N__42785),
            .in2(N__43183),
            .in3(N__40752),
            .lcout(n45),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(n10700),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_633__i1_LC_17_15_1.C_ON=1'b1;
    defparam counter_633__i1_LC_17_15_1.SEQ_MODE=4'b1000;
    defparam counter_633__i1_LC_17_15_1.LUT_INIT=16'b1100101000111010;
    LogicCell40 counter_633__i1_LC_17_15_1 (
            .in0(N__42878),
            .in1(N__42756),
            .in2(N__42433),
            .in3(N__40749),
            .lcout(counter_1),
            .ltout(),
            .carryin(n10700),
            .carryout(n10701),
            .clk(N__46899),
            .ce(N__45981),
            .sr(_gnd_net_));
    defparam counter_633__i2_LC_17_15_2.C_ON=1'b1;
    defparam counter_633__i2_LC_17_15_2.SEQ_MODE=4'b1000;
    defparam counter_633__i2_LC_17_15_2.LUT_INIT=16'b1110001000101110;
    LogicCell40 counter_633__i2_LC_17_15_2 (
            .in0(N__42874),
            .in1(N__42423),
            .in2(N__43092),
            .in3(N__40746),
            .lcout(counter_2),
            .ltout(),
            .carryin(n10701),
            .carryout(n10702),
            .clk(N__46899),
            .ce(N__45981),
            .sr(_gnd_net_));
    defparam counter_633__i3_LC_17_15_3.C_ON=1'b1;
    defparam counter_633__i3_LC_17_15_3.SEQ_MODE=4'b1000;
    defparam counter_633__i3_LC_17_15_3.LUT_INIT=16'b1100101000111010;
    LogicCell40 counter_633__i3_LC_17_15_3 (
            .in0(N__42879),
            .in1(N__43074),
            .in2(N__42434),
            .in3(N__40743),
            .lcout(counter_3),
            .ltout(),
            .carryin(n10702),
            .carryout(n10703),
            .clk(N__46899),
            .ce(N__45981),
            .sr(_gnd_net_));
    defparam counter_633__i4_LC_17_15_4.C_ON=1'b1;
    defparam counter_633__i4_LC_17_15_4.SEQ_MODE=4'b1000;
    defparam counter_633__i4_LC_17_15_4.LUT_INIT=16'b1110001000101110;
    LogicCell40 counter_633__i4_LC_17_15_4 (
            .in0(N__42875),
            .in1(N__42427),
            .in2(N__43119),
            .in3(N__42444),
            .lcout(counter_4),
            .ltout(),
            .carryin(n10703),
            .carryout(n10704),
            .clk(N__46899),
            .ce(N__45981),
            .sr(_gnd_net_));
    defparam counter_633__i5_LC_17_15_5.C_ON=1'b1;
    defparam counter_633__i5_LC_17_15_5.SEQ_MODE=4'b1000;
    defparam counter_633__i5_LC_17_15_5.LUT_INIT=16'b1100101000111010;
    LogicCell40 counter_633__i5_LC_17_15_5 (
            .in0(N__42880),
            .in1(N__43104),
            .in2(N__42435),
            .in3(N__42441),
            .lcout(counter_5),
            .ltout(),
            .carryin(n10704),
            .carryout(n10705),
            .clk(N__46899),
            .ce(N__45981),
            .sr(_gnd_net_));
    defparam counter_633__i6_LC_17_15_6.C_ON=1'b1;
    defparam counter_633__i6_LC_17_15_6.SEQ_MODE=4'b1000;
    defparam counter_633__i6_LC_17_15_6.LUT_INIT=16'b1110001000101110;
    LogicCell40 counter_633__i6_LC_17_15_6 (
            .in0(N__42876),
            .in1(N__42431),
            .in2(N__42771),
            .in3(N__42438),
            .lcout(counter_6),
            .ltout(),
            .carryin(n10705),
            .carryout(n10706),
            .clk(N__46899),
            .ce(N__45981),
            .sr(_gnd_net_));
    defparam counter_633__i7_LC_17_15_7.C_ON=1'b0;
    defparam counter_633__i7_LC_17_15_7.SEQ_MODE=4'b1000;
    defparam counter_633__i7_LC_17_15_7.LUT_INIT=16'b1110010001001110;
    LogicCell40 counter_633__i7_LC_17_15_7 (
            .in0(N__42432),
            .in1(N__42877),
            .in2(N__42801),
            .in3(N__42402),
            .lcout(counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46899),
            .ce(N__45981),
            .sr(_gnd_net_));
    defparam i9193_4_lut_4_lut_LC_17_16_2.C_ON=1'b0;
    defparam i9193_4_lut_4_lut_LC_17_16_2.SEQ_MODE=4'b0000;
    defparam i9193_4_lut_4_lut_LC_17_16_2.LUT_INIT=16'b0000001101110111;
    LogicCell40 i9193_4_lut_4_lut_LC_17_16_2 (
            .in0(N__43128),
            .in1(N__43874),
            .in2(N__47677),
            .in3(N__43641),
            .lcout(n7681),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_190_LC_17_16_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_190_LC_17_16_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_190_LC_17_16_3.LUT_INIT=16'b1100110011001000;
    LogicCell40 i1_2_lut_3_lut_4_lut_4_lut_adj_190_LC_17_16_3 (
            .in0(N__44964),
            .in1(N__47646),
            .in2(N__45569),
            .in3(N__44529),
            .lcout(n11824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7627_2_lut_3_lut_4_lut_4_lut_LC_17_16_6.C_ON=1'b0;
    defparam i7627_2_lut_3_lut_4_lut_4_lut_LC_17_16_6.SEQ_MODE=4'b0000;
    defparam i7627_2_lut_3_lut_4_lut_4_lut_LC_17_16_6.LUT_INIT=16'b1010101010101000;
    LogicCell40 i7627_2_lut_3_lut_4_lut_4_lut_LC_17_16_6 (
            .in0(N__47647),
            .in1(N__45106),
            .in2(N__44113),
            .in3(N__45466),
            .lcout(n11964),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_i0_i0_LC_17_17_0.C_ON=1'b1;
    defparam current_pin_i0_i0_LC_17_17_0.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i0_LC_17_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i0_LC_17_17_0 (
            .in0(_gnd_net_),
            .in1(N__46323),
            .in2(_gnd_net_),
            .in3(N__42369),
            .lcout(current_pin_0),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(n10575),
            .clk(N__46887),
            .ce(N__42456),
            .sr(N__42465));
    defparam current_pin_i0_i1_LC_17_17_1.C_ON=1'b1;
    defparam current_pin_i0_i1_LC_17_17_1.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i1_LC_17_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i1_LC_17_17_1 (
            .in0(_gnd_net_),
            .in1(N__46510),
            .in2(_gnd_net_),
            .in3(N__42366),
            .lcout(current_pin_1),
            .ltout(),
            .carryin(n10575),
            .carryout(n10576),
            .clk(N__46887),
            .ce(N__42456),
            .sr(N__42465));
    defparam current_pin_i0_i2_LC_17_17_2.C_ON=1'b1;
    defparam current_pin_i0_i2_LC_17_17_2.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i2_LC_17_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i2_LC_17_17_2 (
            .in0(_gnd_net_),
            .in1(N__45560),
            .in2(_gnd_net_),
            .in3(N__42519),
            .lcout(current_pin_2),
            .ltout(),
            .carryin(n10576),
            .carryout(n10577),
            .clk(N__46887),
            .ce(N__42456),
            .sr(N__42465));
    defparam current_pin_i0_i3_LC_17_17_3.C_ON=1'b1;
    defparam current_pin_i0_i3_LC_17_17_3.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i3_LC_17_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i3_LC_17_17_3 (
            .in0(_gnd_net_),
            .in1(N__45267),
            .in2(_gnd_net_),
            .in3(N__42516),
            .lcout(current_pin_3),
            .ltout(),
            .carryin(n10577),
            .carryout(n10578),
            .clk(N__46887),
            .ce(N__42456),
            .sr(N__42465));
    defparam current_pin_i0_i4_LC_17_17_4.C_ON=1'b1;
    defparam current_pin_i0_i4_LC_17_17_4.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i4_LC_17_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i4_LC_17_17_4 (
            .in0(_gnd_net_),
            .in1(N__43244),
            .in2(_gnd_net_),
            .in3(N__42513),
            .lcout(current_pin_4),
            .ltout(),
            .carryin(n10578),
            .carryout(n10579),
            .clk(N__46887),
            .ce(N__42456),
            .sr(N__42465));
    defparam current_pin_i0_i5_LC_17_17_5.C_ON=1'b1;
    defparam current_pin_i0_i5_LC_17_17_5.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i5_LC_17_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i5_LC_17_17_5 (
            .in0(_gnd_net_),
            .in1(N__42510),
            .in2(_gnd_net_),
            .in3(N__42498),
            .lcout(current_pin_5),
            .ltout(),
            .carryin(n10579),
            .carryout(n10580),
            .clk(N__46887),
            .ce(N__42456),
            .sr(N__42465));
    defparam current_pin_i0_i6_LC_17_17_6.C_ON=1'b1;
    defparam current_pin_i0_i6_LC_17_17_6.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i6_LC_17_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i6_LC_17_17_6 (
            .in0(_gnd_net_),
            .in1(N__42495),
            .in2(_gnd_net_),
            .in3(N__42483),
            .lcout(current_pin_6),
            .ltout(),
            .carryin(n10580),
            .carryout(n10581),
            .clk(N__46887),
            .ce(N__42456),
            .sr(N__42465));
    defparam current_pin_i0_i7_LC_17_17_7.C_ON=1'b0;
    defparam current_pin_i0_i7_LC_17_17_7.SEQ_MODE=4'b1000;
    defparam current_pin_i0_i7_LC_17_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 current_pin_i0_i7_LC_17_17_7 (
            .in0(_gnd_net_),
            .in1(N__42477),
            .in2(_gnd_net_),
            .in3(N__42480),
            .lcout(current_pin_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46887),
            .ce(N__42456),
            .sr(N__42465));
    defparam i4198_2_lut_3_lut_4_lut_LC_17_18_0.C_ON=1'b0;
    defparam i4198_2_lut_3_lut_4_lut_LC_17_18_0.SEQ_MODE=4'b0000;
    defparam i4198_2_lut_3_lut_4_lut_LC_17_18_0.LUT_INIT=16'b1111110100000000;
    LogicCell40 i4198_2_lut_3_lut_4_lut_LC_17_18_0 (
            .in0(N__43911),
            .in1(N__43640),
            .in2(N__47658),
            .in3(N__42455),
            .lcout(n7985),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9181_2_lut_4_lut_LC_17_18_3.C_ON=1'b0;
    defparam i9181_2_lut_4_lut_LC_17_18_3.SEQ_MODE=4'b0000;
    defparam i9181_2_lut_4_lut_LC_17_18_3.LUT_INIT=16'b0000001000000011;
    LogicCell40 i9181_2_lut_4_lut_LC_17_18_3 (
            .in0(N__43174),
            .in1(N__47586),
            .in2(N__43668),
            .in3(N__43910),
            .lcout(n7635),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_17_18_4.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_17_18_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_17_18_4.LUT_INIT=16'b1100110011101100;
    LogicCell40 i1_3_lut_4_lut_LC_17_18_4 (
            .in0(N__43414),
            .in1(N__44891),
            .in2(N__45597),
            .in3(N__42588),
            .lcout(),
            .ltout(n9_adj_824_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i7_LC_17_18_5.C_ON=1'b0;
    defparam pin_output_i0_i7_LC_17_18_5.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i7_LC_17_18_5.LUT_INIT=16'b0111111100100000;
    LogicCell40 pin_output_i0_i7_LC_17_18_5 (
            .in0(N__45971),
            .in1(N__46098),
            .in2(N__42741),
            .in3(N__42946),
            .lcout(pin_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46895),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_167_LC_17_18_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_167_LC_17_18_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_167_LC_17_18_6.LUT_INIT=16'b1100110011011100;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_167_LC_17_18_6 (
            .in0(N__44995),
            .in1(N__44890),
            .in2(N__45596),
            .in3(N__42587),
            .lcout(),
            .ltout(n8_adj_822_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i5_LC_17_18_7.C_ON=1'b0;
    defparam pin_output_i0_i5_LC_17_18_7.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i5_LC_17_18_7.LUT_INIT=16'b0111111100100000;
    LogicCell40 pin_output_i0_i5_LC_17_18_7 (
            .in0(N__45970),
            .in1(N__46097),
            .in2(N__42738),
            .in3(N__42724),
            .lcout(pin_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46895),
            .ce(),
            .sr(_gnd_net_));
    defparam i8962_3_lut_LC_17_19_3.C_ON=1'b0;
    defparam i8962_3_lut_LC_17_19_3.SEQ_MODE=4'b0000;
    defparam i8962_3_lut_LC_17_19_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 i8962_3_lut_LC_17_19_3 (
            .in0(N__46344),
            .in1(N__42728),
            .in2(_gnd_net_),
            .in3(N__42698),
            .lcout(),
            .ltout(n13357_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_1__bdd_4_lut_9236_LC_17_19_4.C_ON=1'b0;
    defparam current_pin_1__bdd_4_lut_9236_LC_17_19_4.SEQ_MODE=4'b0000;
    defparam current_pin_1__bdd_4_lut_9236_LC_17_19_4.LUT_INIT=16'b1110110001100100;
    LogicCell40 current_pin_1__bdd_4_lut_9236_LC_17_19_4 (
            .in0(N__45487),
            .in1(N__46511),
            .in2(N__42675),
            .in3(N__42894),
            .lcout(n13625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_234_i6_2_lut_LC_17_19_6.C_ON=1'b0;
    defparam equal_234_i6_2_lut_LC_17_19_6.SEQ_MODE=4'b0000;
    defparam equal_234_i6_2_lut_LC_17_19_6.LUT_INIT=16'b1111111100110011;
    LogicCell40 equal_234_i6_2_lut_LC_17_19_6 (
            .in0(_gnd_net_),
            .in1(N__46512),
            .in2(_gnd_net_),
            .in3(N__46345),
            .lcout(n6_adj_810),
            .ltout(n6_adj_810_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7543_2_lut_3_lut_4_lut_LC_17_19_7.C_ON=1'b0;
    defparam i7543_2_lut_3_lut_4_lut_LC_17_19_7.SEQ_MODE=4'b0000;
    defparam i7543_2_lut_3_lut_4_lut_LC_17_19_7.LUT_INIT=16'b1111110111111111;
    LogicCell40 i7543_2_lut_3_lut_4_lut_LC_17_19_7 (
            .in0(N__43248),
            .in1(N__45268),
            .in2(N__42666),
            .in3(N__45488),
            .lcout(n11874),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_188_LC_17_20_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_188_LC_17_20_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_188_LC_17_20_1.LUT_INIT=16'b1100110011001000;
    LogicCell40 i1_2_lut_3_lut_4_lut_4_lut_adj_188_LC_17_20_1 (
            .in0(N__44530),
            .in1(N__47636),
            .in2(N__44114),
            .in3(N__45507),
            .lcout(n11823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_168_LC_17_20_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_168_LC_17_20_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_168_LC_17_20_3.LUT_INIT=16'b1111000011110100;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_168_LC_17_20_3 (
            .in0(N__44388),
            .in1(N__45508),
            .in2(N__44909),
            .in3(N__42615),
            .lcout(),
            .ltout(n7_adj_823_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i6_LC_17_20_4.C_ON=1'b0;
    defparam pin_output_i0_i6_LC_17_20_4.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i6_LC_17_20_4.LUT_INIT=16'b0010101011101010;
    LogicCell40 pin_output_i0_i6_LC_17_20_4 (
            .in0(N__42908),
            .in1(N__45974),
            .in2(N__42993),
            .in3(N__46144),
            .lcout(pin_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46903),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i19_LC_17_20_5.C_ON=1'b0;
    defparam pin_output_enable__i19_LC_17_20_5.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i19_LC_17_20_5.LUT_INIT=16'b1101110010001100;
    LogicCell40 pin_output_enable__i19_LC_17_20_5 (
            .in0(N__43365),
            .in1(N__42977),
            .in2(N__47149),
            .in3(N__47637),
            .lcout(pin_oe_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46903),
            .ce(),
            .sr(_gnd_net_));
    defparam i8963_3_lut_LC_17_20_7.C_ON=1'b0;
    defparam i8963_3_lut_LC_17_20_7.SEQ_MODE=4'b0000;
    defparam i8963_3_lut_LC_17_20_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 i8963_3_lut_LC_17_20_7 (
            .in0(N__46343),
            .in1(N__42950),
            .in2(_gnd_net_),
            .in3(N__42907),
            .lcout(n13358),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_165_LC_17_21_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_165_LC_17_21_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_165_LC_17_21_3.LUT_INIT=16'b1100110011001101;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_165_LC_17_21_3 (
            .in0(N__44107),
            .in1(N__44907),
            .in2(N__45587),
            .in3(N__44531),
            .lcout(n8_adj_826),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_LC_18_14_2.C_ON=1'b0;
    defparam i2_3_lut_LC_18_14_2.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_18_14_2.LUT_INIT=16'b0000000001000100;
    LogicCell40 i2_3_lut_LC_18_14_2 (
            .in0(N__43824),
            .in1(N__47329),
            .in2(_gnd_net_),
            .in3(N__43588),
            .lcout(n3762),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i16_LC_18_14_5.C_ON=1'b0;
    defparam pin_output_enable__i16_LC_18_14_5.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i16_LC_18_14_5.LUT_INIT=16'b1011100010101010;
    LogicCell40 pin_output_enable__i16_LC_18_14_5 (
            .in0(N__42818),
            .in1(N__42843),
            .in2(N__47460),
            .in3(N__47122),
            .lcout(pin_oe_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46908),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_202_LC_18_15_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_202_LC_18_15_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_202_LC_18_15_2.LUT_INIT=16'b1010101010001010;
    LogicCell40 i1_2_lut_3_lut_4_lut_4_lut_adj_202_LC_18_15_2 (
            .in0(N__47479),
            .in1(N__44112),
            .in2(N__45642),
            .in3(N__44537),
            .lcout(n11820),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_18_15_5.C_ON=1'b0;
    defparam i2_2_lut_LC_18_15_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_18_15_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i2_2_lut_LC_18_15_5 (
            .in0(_gnd_net_),
            .in1(N__42797),
            .in2(_gnd_net_),
            .in3(N__42786),
            .lcout(),
            .ltout(n10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9165_4_lut_LC_18_15_6.C_ON=1'b0;
    defparam i9165_4_lut_LC_18_15_6.SEQ_MODE=4'b0000;
    defparam i9165_4_lut_LC_18_15_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i9165_4_lut_LC_18_15_6 (
            .in0(N__42767),
            .in1(N__42755),
            .in2(N__42744),
            .in3(N__43062),
            .lcout(state_7_N_167_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_179_LC_18_15_7.C_ON=1'b0;
    defparam i6_4_lut_adj_179_LC_18_15_7.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_179_LC_18_15_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_179_LC_18_15_7 (
            .in0(N__43115),
            .in1(N__43103),
            .in2(N__43091),
            .in3(N__43073),
            .lcout(n14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8975_3_lut_LC_18_16_0.C_ON=1'b0;
    defparam i8975_3_lut_LC_18_16_0.SEQ_MODE=4'b0000;
    defparam i8975_3_lut_LC_18_16_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i8975_3_lut_LC_18_16_0 (
            .in0(N__43042),
            .in1(N__43009),
            .in2(_gnd_net_),
            .in3(N__46320),
            .lcout(n13370),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i11_LC_18_16_3.C_ON=1'b0;
    defparam pin_output_i0_i11_LC_18_16_3.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i11_LC_18_16_3.LUT_INIT=16'b0101110011001100;
    LogicCell40 pin_output_i0_i11_LC_18_16_3 (
            .in0(N__46094),
            .in1(N__43043),
            .in2(N__44199),
            .in3(N__45994),
            .lcout(pin_out_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46900),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_163_LC_18_16_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_163_LC_18_16_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_163_LC_18_16_5.LUT_INIT=16'b1010101010101011;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_163_LC_18_16_5 (
            .in0(N__44854),
            .in1(N__44426),
            .in2(N__45643),
            .in3(N__44534),
            .lcout(),
            .ltout(n7_adj_827_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i10_LC_18_16_6.C_ON=1'b0;
    defparam pin_output_i0_i10_LC_18_16_6.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i10_LC_18_16_6.LUT_INIT=16'b0111111100100000;
    LogicCell40 pin_output_i0_i10_LC_18_16_6 (
            .in0(N__45993),
            .in1(N__46095),
            .in2(N__43029),
            .in3(N__43010),
            .lcout(pin_out_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46900),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_160_LC_18_16_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_160_LC_18_16_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_160_LC_18_16_7.LUT_INIT=16'b1010101010101110;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_160_LC_18_16_7 (
            .in0(N__44853),
            .in1(N__45461),
            .in2(N__44996),
            .in3(N__44533),
            .lcout(n7_adj_830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_161_LC_18_17_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_161_LC_18_17_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_161_LC_18_17_0.LUT_INIT=16'b1100110011001110;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_161_LC_18_17_0 (
            .in0(N__45556),
            .in1(N__44878),
            .in2(N__44111),
            .in3(N__44535),
            .lcout(n8_adj_829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5882_2_lut_3_lut_4_lut_LC_18_17_2.C_ON=1'b0;
    defparam i5882_2_lut_3_lut_4_lut_LC_18_17_2.SEQ_MODE=4'b0000;
    defparam i5882_2_lut_3_lut_4_lut_LC_18_17_2.LUT_INIT=16'b1111111111111011;
    LogicCell40 i5882_2_lut_3_lut_4_lut_LC_18_17_2 (
            .in0(N__47478),
            .in1(N__43891),
            .in2(N__43651),
            .in3(N__43302),
            .lcout(n9675),
            .ltout(n9675_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i15_LC_18_17_3.C_ON=1'b0;
    defparam pin_output_i0_i15_LC_18_17_3.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i15_LC_18_17_3.LUT_INIT=16'b0111111100001000;
    LogicCell40 pin_output_i0_i15_LC_18_17_3 (
            .in0(N__45979),
            .in1(N__43308),
            .in2(N__42996),
            .in3(N__45787),
            .lcout(pin_out_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46892),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_162_LC_18_17_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_162_LC_18_17_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_162_LC_18_17_4.LUT_INIT=16'b1100110011101100;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_162_LC_18_17_4 (
            .in0(N__43431),
            .in1(N__44879),
            .in2(N__45634),
            .in3(N__44536),
            .lcout(n8_adj_832),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_4_lut_LC_18_17_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_4_lut_LC_18_17_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_4_lut_LC_18_17_7.LUT_INIT=16'b1111000011100000;
    LogicCell40 i1_2_lut_3_lut_4_lut_4_lut_LC_18_17_7 (
            .in0(N__45462),
            .in1(N__44991),
            .in2(N__47600),
            .in3(N__45062),
            .lcout(n11822),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9145_4_lut_LC_18_18_0.C_ON=1'b0;
    defparam i9145_4_lut_LC_18_18_0.SEQ_MODE=4'b0000;
    defparam i9145_4_lut_LC_18_18_0.LUT_INIT=16'b0011000010111000;
    LogicCell40 i9145_4_lut_LC_18_18_0 (
            .in0(N__44676),
            .in1(N__43236),
            .in2(N__43257),
            .in3(N__45251),
            .lcout(pin_out_22__N_216),
            .ltout(pin_out_22__N_216_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9155_4_lut_LC_18_18_1.C_ON=1'b0;
    defparam i9155_4_lut_LC_18_18_1.SEQ_MODE=4'b0000;
    defparam i9155_4_lut_LC_18_18_1.LUT_INIT=16'b0010110101111000;
    LogicCell40 i9155_4_lut_LC_18_18_1 (
            .in0(N__43237),
            .in1(N__45201),
            .in2(N__43296),
            .in3(N__44124),
            .lcout(n13551),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13637_bdd_4_lut_LC_18_18_4.C_ON=1'b0;
    defparam n13637_bdd_4_lut_LC_18_18_4.SEQ_MODE=4'b0000;
    defparam n13637_bdd_4_lut_LC_18_18_4.LUT_INIT=16'b1110111001010000;
    LogicCell40 n13637_bdd_4_lut_LC_18_18_4 (
            .in0(N__45452),
            .in1(N__43293),
            .in2(N__43284),
            .in3(N__46206),
            .lcout(),
            .ltout(n13640_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9144_3_lut_LC_18_18_5.C_ON=1'b0;
    defparam i9144_3_lut_LC_18_18_5.SEQ_MODE=4'b0000;
    defparam i9144_3_lut_LC_18_18_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 i9144_3_lut_LC_18_18_5 (
            .in0(N__45250),
            .in1(_gnd_net_),
            .in2(N__43272),
            .in3(N__43269),
            .lcout(n13540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_224_i7_2_lut_LC_18_18_6.C_ON=1'b0;
    defparam equal_224_i7_2_lut_LC_18_18_6.SEQ_MODE=4'b0000;
    defparam equal_224_i7_2_lut_LC_18_18_6.LUT_INIT=16'b1111111100110011;
    LogicCell40 equal_224_i7_2_lut_LC_18_18_6 (
            .in0(_gnd_net_),
            .in1(N__43238),
            .in2(_gnd_net_),
            .in3(N__45252),
            .lcout(n7_adj_797),
            .ltout(n7_adj_797_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_199_LC_18_18_7.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_199_LC_18_18_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_199_LC_18_18_7.LUT_INIT=16'b1010101010101110;
    LogicCell40 i1_2_lut_4_lut_adj_199_LC_18_18_7 (
            .in0(N__44886),
            .in1(N__43424),
            .in2(N__43200),
            .in3(N__45453),
            .lcout(n8_adj_836),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i41_4_lut_LC_18_19_4.C_ON=1'b0;
    defparam i41_4_lut_LC_18_19_4.SEQ_MODE=4'b0000;
    defparam i41_4_lut_LC_18_19_4.LUT_INIT=16'b0000000110101011;
    LogicCell40 i41_4_lut_LC_18_19_4 (
            .in0(N__47583),
            .in1(N__43197),
            .in2(N__43185),
            .in3(N__43976),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_189_LC_18_19_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_189_LC_18_19_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_189_LC_18_19_5.LUT_INIT=16'b1100010011001100;
    LogicCell40 i1_2_lut_3_lut_4_lut_4_lut_adj_189_LC_18_19_5 (
            .in0(N__43430),
            .in1(N__47584),
            .in2(N__44544),
            .in3(N__45574),
            .lcout(),
            .ltout(n11825_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i15_LC_18_19_6.C_ON=1'b0;
    defparam pin_output_enable__i15_LC_18_19_6.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i15_LC_18_19_6.LUT_INIT=16'b1100101011001100;
    LogicCell40 pin_output_enable__i15_LC_18_19_6 (
            .in0(N__47585),
            .in1(N__43988),
            .in2(N__44007),
            .in3(N__47123),
            .lcout(pin_oe_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46904),
            .ce(),
            .sr(_gnd_net_));
    defparam i4262_2_lut_3_lut_4_lut_LC_18_19_7.C_ON=1'b0;
    defparam i4262_2_lut_3_lut_4_lut_LC_18_19_7.SEQ_MODE=4'b0000;
    defparam i4262_2_lut_3_lut_4_lut_LC_18_19_7.LUT_INIT=16'b0000000010000000;
    LogicCell40 i4262_2_lut_3_lut_4_lut_LC_18_19_7 (
            .in0(N__43977),
            .in1(N__47582),
            .in2(N__43912),
            .in3(N__43625),
            .lcout(n8025),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7617_2_lut_3_lut_4_lut_4_lut_LC_18_20_0.C_ON=1'b0;
    defparam i7617_2_lut_3_lut_4_lut_4_lut_LC_18_20_0.SEQ_MODE=4'b0000;
    defparam i7617_2_lut_3_lut_4_lut_4_lut_LC_18_20_0.LUT_INIT=16'b1110111100000000;
    LogicCell40 i7617_2_lut_3_lut_4_lut_4_lut_LC_18_20_0 (
            .in0(N__44105),
            .in1(N__45101),
            .in2(N__45641),
            .in3(N__47641),
            .lcout(),
            .ltout(n11954_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i20_LC_18_20_1.C_ON=1'b0;
    defparam pin_output_enable__i20_LC_18_20_1.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i20_LC_18_20_1.LUT_INIT=16'b1010110010101010;
    LogicCell40 pin_output_enable__i20_LC_18_20_1 (
            .in0(N__43442),
            .in1(N__47642),
            .in2(N__43458),
            .in3(N__47130),
            .lcout(pin_oe_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46909),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_4_lut_LC_18_20_5.C_ON=1'b0;
    defparam i1_2_lut_4_lut_4_lut_LC_18_20_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_4_lut_LC_18_20_5.LUT_INIT=16'b1111000011010000;
    LogicCell40 i1_2_lut_4_lut_4_lut_LC_18_20_5 (
            .in0(N__43428),
            .in1(N__45570),
            .in2(N__47676),
            .in3(N__45091),
            .lcout(n11821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_177_LC_18_21_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_177_LC_18_21_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_177_LC_18_21_6.LUT_INIT=16'b1100110111001100;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_177_LC_18_21_6 (
            .in0(N__45100),
            .in1(N__44908),
            .in2(N__44115),
            .in3(N__45668),
            .lcout(n7_adj_837),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i8_LC_18_22_5.C_ON=1'b0;
    defparam pin_output_i0_i8_LC_18_22_5.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i8_LC_18_22_5.LUT_INIT=16'b0111001011110000;
    LogicCell40 pin_output_i0_i8_LC_18_22_5 (
            .in0(N__43359),
            .in1(N__46141),
            .in2(N__43336),
            .in3(N__45980),
            .lcout(pin_out_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46919),
            .ce(),
            .sr(_gnd_net_));
    defparam i7625_2_lut_3_lut_4_lut_4_lut_LC_19_15_6.C_ON=1'b0;
    defparam i7625_2_lut_3_lut_4_lut_4_lut_LC_19_15_6.SEQ_MODE=4'b0000;
    defparam i7625_2_lut_3_lut_4_lut_4_lut_LC_19_15_6.LUT_INIT=16'b1100110010001100;
    LogicCell40 i7625_2_lut_3_lut_4_lut_4_lut_LC_19_15_6 (
            .in0(N__44431),
            .in1(N__47481),
            .in2(N__45669),
            .in3(N__44539),
            .lcout(),
            .ltout(n11962_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i14_LC_19_15_7.C_ON=1'b0;
    defparam pin_output_enable__i14_LC_19_15_7.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i14_LC_19_15_7.LUT_INIT=16'b1100101011001100;
    LogicCell40 pin_output_enable__i14_LC_19_15_7 (
            .in0(N__47482),
            .in1(N__44231),
            .in2(N__44250),
            .in3(N__47119),
            .lcout(pin_oe_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46910),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_198_LC_19_16_4.C_ON=1'b0;
    defparam i1_2_lut_adj_198_LC_19_16_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_198_LC_19_16_4.LUT_INIT=16'b1111111100110011;
    LogicCell40 i1_2_lut_adj_198_LC_19_16_4 (
            .in0(_gnd_net_),
            .in1(N__44220),
            .in2(_gnd_net_),
            .in3(N__44871),
            .lcout(n8_adj_828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7621_2_lut_3_lut_4_lut_4_lut_LC_19_16_5.C_ON=1'b0;
    defparam i7621_2_lut_3_lut_4_lut_4_lut_LC_19_16_5.SEQ_MODE=4'b0000;
    defparam i7621_2_lut_3_lut_4_lut_4_lut_LC_19_16_5.LUT_INIT=16'b1100110010001100;
    LogicCell40 i7621_2_lut_3_lut_4_lut_4_lut_LC_19_16_5 (
            .in0(N__44981),
            .in1(N__47483),
            .in2(N__45670),
            .in3(N__45105),
            .lcout(),
            .ltout(n11958_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i21_LC_19_16_6.C_ON=1'b0;
    defparam pin_output_enable__i21_LC_19_16_6.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i21_LC_19_16_6.LUT_INIT=16'b1100101011001100;
    LogicCell40 pin_output_enable__i21_LC_19_16_6 (
            .in0(N__47484),
            .in1(N__44168),
            .in2(N__44190),
            .in3(N__47124),
            .lcout(pin_oe_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46905),
            .ce(),
            .sr(_gnd_net_));
    defparam i9140_3_lut_LC_19_17_1.C_ON=1'b0;
    defparam i9140_3_lut_LC_19_17_1.SEQ_MODE=4'b0000;
    defparam i9140_3_lut_LC_19_17_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i9140_3_lut_LC_19_17_1 (
            .in0(N__45534),
            .in1(N__45117),
            .in2(_gnd_net_),
            .in3(N__44157),
            .lcout(),
            .ltout(n13536_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9146_3_lut_LC_19_17_2.C_ON=1'b0;
    defparam i9146_3_lut_LC_19_17_2.SEQ_MODE=4'b0000;
    defparam i9146_3_lut_LC_19_17_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 i9146_3_lut_LC_19_17_2 (
            .in0(_gnd_net_),
            .in1(N__45261),
            .in2(N__44139),
            .in3(N__44136),
            .lcout(n13542),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_LC_19_17_3.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_19_17_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_19_17_3.LUT_INIT=16'b1111111100010000;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_19_17_3 (
            .in0(N__44538),
            .in1(N__44422),
            .in2(N__45615),
            .in3(N__44902),
            .lcout(),
            .ltout(n7_adj_831_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i14_LC_19_17_4.C_ON=1'b0;
    defparam pin_output_i0_i14_LC_19_17_4.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i14_LC_19_17_4.LUT_INIT=16'b0111111100100000;
    LogicCell40 pin_output_i0_i14_LC_19_17_4 (
            .in0(N__45995),
            .in1(N__46137),
            .in2(N__44118),
            .in3(N__45752),
            .lcout(pin_out_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46896),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_201_LC_19_17_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_201_LC_19_17_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_201_LC_19_17_6.LUT_INIT=16'b1111000011110001;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_201_LC_19_17_6 (
            .in0(N__45090),
            .in1(N__44095),
            .in2(N__44912),
            .in3(N__45538),
            .lcout(),
            .ltout(n7_adj_833_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i16_LC_19_17_7.C_ON=1'b0;
    defparam pin_output_i0_i16_LC_19_17_7.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i16_LC_19_17_7.LUT_INIT=16'b0111111101000000;
    LogicCell40 pin_output_i0_i16_LC_19_17_7 (
            .in0(N__46136),
            .in1(N__45996),
            .in2(N__44553),
            .in3(N__44698),
            .lcout(pin_out_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46896),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i19_LC_19_18_5.C_ON=1'b0;
    defparam pin_output_i0_i19_LC_19_18_5.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i19_LC_19_18_5.LUT_INIT=16'b0111001011110000;
    LogicCell40 pin_output_i0_i19_LC_19_18_5 (
            .in0(N__44550),
            .in1(N__46096),
            .in2(N__44278),
            .in3(N__45959),
            .lcout(pin_out_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46906),
            .ce(),
            .sr(_gnd_net_));
    defparam i7619_2_lut_3_lut_4_lut_4_lut_LC_19_18_7.C_ON=1'b0;
    defparam i7619_2_lut_3_lut_4_lut_4_lut_LC_19_18_7.SEQ_MODE=4'b0000;
    defparam i7619_2_lut_3_lut_4_lut_4_lut_LC_19_18_7.LUT_INIT=16'b1110111100000000;
    LogicCell40 i7619_2_lut_3_lut_4_lut_4_lut_LC_19_18_7 (
            .in0(N__44540),
            .in1(N__45010),
            .in2(N__45652),
            .in3(N__47480),
            .lcout(n11956),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_178_LC_19_19_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_178_LC_19_19_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_178_LC_19_19_6.LUT_INIT=16'b1010101010101011;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_178_LC_19_19_6 (
            .in0(N__44903),
            .in1(N__44405),
            .in2(N__45654),
            .in3(N__45089),
            .lcout(),
            .ltout(n7_adj_835_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i18_LC_19_19_7.C_ON=1'b0;
    defparam pin_output_i0_i18_LC_19_19_7.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i18_LC_19_19_7.LUT_INIT=16'b0011101010101010;
    LogicCell40 pin_output_i0_i18_LC_19_19_7 (
            .in0(N__44309),
            .in1(N__46110),
            .in2(N__44442),
            .in3(N__45960),
            .lcout(pin_out_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46911),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_19_20_2.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_19_20_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_19_20_2.LUT_INIT=16'b1111000111110000;
    LogicCell40 i1_2_lut_4_lut_LC_19_20_2 (
            .in0(N__44421),
            .in1(N__45099),
            .in2(N__44910),
            .in3(N__45611),
            .lcout(),
            .ltout(n7_adj_839_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i22_LC_19_20_3.C_ON=1'b0;
    defparam pin_output_i0_i22_LC_19_20_3.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i22_LC_19_20_3.LUT_INIT=16'b0111111100100000;
    LogicCell40 pin_output_i0_i22_LC_19_20_3 (
            .in0(N__45956),
            .in1(N__46111),
            .in2(N__44328),
            .in3(N__44581),
            .lcout(pin_out_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46914),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_0__bdd_4_lut_9241_LC_19_20_4.C_ON=1'b0;
    defparam current_pin_0__bdd_4_lut_9241_LC_19_20_4.SEQ_MODE=4'b0000;
    defparam current_pin_0__bdd_4_lut_9241_LC_19_20_4.LUT_INIT=16'b1111001110001000;
    LogicCell40 current_pin_0__bdd_4_lut_9241_LC_19_20_4 (
            .in0(N__44308),
            .in1(N__46559),
            .in2(N__44282),
            .in3(N__46392),
            .lcout(n13631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_176_LC_19_20_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_176_LC_19_20_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_176_LC_19_20_5.LUT_INIT=16'b1111111100010000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_176_LC_19_20_5 (
            .in0(N__45098),
            .in1(N__45006),
            .in2(N__45653),
            .in3(N__44892),
            .lcout(n7_adj_838),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_200_LC_19_21_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_200_LC_19_21_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_200_LC_19_21_1.LUT_INIT=16'b1111111100000001;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_200_LC_19_21_1 (
            .in0(N__45108),
            .in1(N__45019),
            .in2(N__45650),
            .in3(N__44911),
            .lcout(),
            .ltout(n8_adj_834_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i17_LC_19_21_2.C_ON=1'b0;
    defparam pin_output_i0_i17_LC_19_21_2.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i17_LC_19_21_2.LUT_INIT=16'b0100110011101100;
    LogicCell40 pin_output_i0_i17_LC_19_21_2 (
            .in0(N__45957),
            .in1(N__44738),
            .in2(N__44754),
            .in3(N__46139),
            .lcout(pin_out_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46920),
            .ce(),
            .sr(_gnd_net_));
    defparam n13631_bdd_4_lut_LC_19_21_3.C_ON=1'b0;
    defparam n13631_bdd_4_lut_LC_19_21_3.SEQ_MODE=4'b0000;
    defparam n13631_bdd_4_lut_LC_19_21_3.LUT_INIT=16'b1100110010111000;
    LogicCell40 n13631_bdd_4_lut_LC_19_21_3 (
            .in0(N__44737),
            .in1(N__44724),
            .in2(N__44708),
            .in3(N__46563),
            .lcout(),
            .ltout(n13634_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8994_3_lut_LC_19_21_4.C_ON=1'b0;
    defparam i8994_3_lut_LC_19_21_4.SEQ_MODE=4'b0000;
    defparam i8994_3_lut_LC_19_21_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 i8994_3_lut_LC_19_21_4 (
            .in0(_gnd_net_),
            .in1(N__45598),
            .in2(N__44679),
            .in3(N__44559),
            .lcout(n13389),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i21_LC_19_21_7.C_ON=1'b0;
    defparam pin_output_i0_i21_LC_19_21_7.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i21_LC_19_21_7.LUT_INIT=16'b0111010011110000;
    LogicCell40 pin_output_i0_i21_LC_19_21_7 (
            .in0(N__46138),
            .in1(N__44667),
            .in2(N__44642),
            .in3(N__45958),
            .lcout(pin_out_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46920),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i20_LC_19_22_0.C_ON=1'b0;
    defparam pin_output_i0_i20_LC_19_22_0.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i20_LC_19_22_0.LUT_INIT=16'b0111000011111000;
    LogicCell40 pin_output_i0_i20_LC_19_22_0 (
            .in0(N__45952),
            .in1(N__44661),
            .in2(N__44615),
            .in3(N__46140),
            .lcout(pin_out_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46922),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_4__I_0_i19_3_lut_LC_19_22_1.C_ON=1'b0;
    defparam current_pin_4__I_0_i19_3_lut_LC_19_22_1.SEQ_MODE=4'b0000;
    defparam current_pin_4__I_0_i19_3_lut_LC_19_22_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 current_pin_4__I_0_i19_3_lut_LC_19_22_1 (
            .in0(N__44635),
            .in1(N__44608),
            .in2(_gnd_net_),
            .in3(N__46408),
            .lcout(),
            .ltout(n19_adj_790_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8993_4_lut_LC_19_22_2.C_ON=1'b0;
    defparam i8993_4_lut_LC_19_22_2.SEQ_MODE=4'b0000;
    defparam i8993_4_lut_LC_19_22_2.LUT_INIT=16'b0100010011110000;
    LogicCell40 i8993_4_lut_LC_19_22_2 (
            .in0(N__46409),
            .in1(N__44585),
            .in2(N__44562),
            .in3(N__46571),
            .lcout(n13388),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8980_3_lut_LC_20_17_0.C_ON=1'b0;
    defparam i8980_3_lut_LC_20_17_0.SEQ_MODE=4'b0000;
    defparam i8980_3_lut_LC_20_17_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 i8980_3_lut_LC_20_17_0 (
            .in0(N__45811),
            .in1(N__46165),
            .in2(_gnd_net_),
            .in3(N__46336),
            .lcout(),
            .ltout(n13375_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_1__bdd_4_lut_LC_20_17_1.C_ON=1'b0;
    defparam current_pin_1__bdd_4_lut_LC_20_17_1.SEQ_MODE=4'b0000;
    defparam current_pin_1__bdd_4_lut_LC_20_17_1.LUT_INIT=16'b1110110001100100;
    LogicCell40 current_pin_1__bdd_4_lut_LC_20_17_1 (
            .in0(N__45492),
            .in1(N__46513),
            .in2(N__46209),
            .in3(N__45735),
            .lcout(n13637),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i12_LC_20_17_2.C_ON=1'b0;
    defparam pin_output_i0_i12_LC_20_17_2.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i12_LC_20_17_2.LUT_INIT=16'b0100111011001100;
    LogicCell40 pin_output_i0_i12_LC_20_17_2 (
            .in0(N__46194),
            .in1(N__46166),
            .in2(N__46151),
            .in3(N__45978),
            .lcout(pin_out_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46901),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_i0_i13_LC_20_17_3.C_ON=1'b0;
    defparam pin_output_i0_i13_LC_20_17_3.SEQ_MODE=4'b1000;
    defparam pin_output_i0_i13_LC_20_17_3.LUT_INIT=16'b0111111101000000;
    LogicCell40 pin_output_i0_i13_LC_20_17_3 (
            .in0(N__46132),
            .in1(N__46008),
            .in2(N__45992),
            .in3(N__45812),
            .lcout(pin_out_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46901),
            .ce(),
            .sr(_gnd_net_));
    defparam i8981_3_lut_LC_20_17_6.C_ON=1'b0;
    defparam i8981_3_lut_LC_20_17_6.SEQ_MODE=4'b0000;
    defparam i8981_3_lut_LC_20_17_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i8981_3_lut_LC_20_17_6 (
            .in0(N__45788),
            .in1(N__45751),
            .in2(_gnd_net_),
            .in3(N__46335),
            .lcout(n13376),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i13_LC_20_18_0.C_ON=1'b0;
    defparam pin_output_enable__i13_LC_20_18_0.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i13_LC_20_18_0.LUT_INIT=16'b1101100011001100;
    LogicCell40 pin_output_enable__i13_LC_20_18_0 (
            .in0(N__45729),
            .in1(N__45707),
            .in2(N__47659),
            .in3(N__47147),
            .lcout(pin_oe_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46912),
            .ce(),
            .sr(_gnd_net_));
    defparam i9075_4_lut_LC_20_21_3.C_ON=1'b0;
    defparam i9075_4_lut_LC_20_21_3.SEQ_MODE=4'b0000;
    defparam i9075_4_lut_LC_20_21_3.LUT_INIT=16'b0000000010101100;
    LogicCell40 i9075_4_lut_LC_20_21_3 (
            .in0(N__46656),
            .in1(N__46605),
            .in2(N__45651),
            .in3(N__45269),
            .lcout(n13465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_0__bdd_4_lut_9246_LC_21_17_1.C_ON=1'b0;
    defparam current_pin_0__bdd_4_lut_9246_LC_21_17_1.SEQ_MODE=4'b0000;
    defparam current_pin_0__bdd_4_lut_9246_LC_21_17_1.LUT_INIT=16'b1011100011001100;
    LogicCell40 current_pin_0__bdd_4_lut_9246_LC_21_17_1 (
            .in0(N__45189),
            .in1(N__46337),
            .in2(N__45174),
            .in3(N__46522),
            .lcout(),
            .ltout(n13643_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13643_bdd_4_lut_LC_21_17_2.C_ON=1'b0;
    defparam n13643_bdd_4_lut_LC_21_17_2.SEQ_MODE=4'b0000;
    defparam n13643_bdd_4_lut_LC_21_17_2.LUT_INIT=16'b1110010111100000;
    LogicCell40 n13643_bdd_4_lut_LC_21_17_2 (
            .in0(N__46523),
            .in1(N__45150),
            .in2(N__45138),
            .in3(N__45135),
            .lcout(n13646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pin_output_enable__i17_LC_21_17_4.C_ON=1'b0;
    defparam pin_output_enable__i17_LC_21_17_4.SEQ_MODE=4'b1000;
    defparam pin_output_enable__i17_LC_21_17_4.LUT_INIT=16'b1101100011001100;
    LogicCell40 pin_output_enable__i17_LC_21_17_4 (
            .in0(N__47706),
            .in1(N__46934),
            .in2(N__47663),
            .in3(N__47148),
            .lcout(pin_oe_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46907),
            .ce(),
            .sr(_gnd_net_));
    defparam i8957_4_lut_LC_23_32_1.C_ON=1'b0;
    defparam i8957_4_lut_LC_23_32_1.SEQ_MODE=4'b0000;
    defparam i8957_4_lut_LC_23_32_1.LUT_INIT=16'b0010111000100010;
    LogicCell40 i8957_4_lut_LC_23_32_1 (
            .in0(N__46215),
            .in1(N__46572),
            .in2(N__46419),
            .in3(N__46662),
            .lcout(n13352),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n13607_bdd_4_lut_LC_24_27_6.C_ON=1'b0;
    defparam n13607_bdd_4_lut_LC_24_27_6.SEQ_MODE=4'b0000;
    defparam n13607_bdd_4_lut_LC_24_27_6.LUT_INIT=16'b1100110010111000;
    LogicCell40 n13607_bdd_4_lut_LC_24_27_6 (
            .in0(N__46644),
            .in1(N__46428),
            .in2(N__46632),
            .in3(N__46555),
            .lcout(n13610),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam current_pin_0__bdd_4_lut_9231_LC_24_32_0.C_ON=1'b0;
    defparam current_pin_0__bdd_4_lut_9231_LC_24_32_0.SEQ_MODE=4'b0000;
    defparam current_pin_0__bdd_4_lut_9231_LC_24_32_0.LUT_INIT=16'b1101100010101010;
    LogicCell40 current_pin_0__bdd_4_lut_9231_LC_24_32_0 (
            .in0(N__46411),
            .in1(N__46593),
            .in2(N__46587),
            .in3(N__46567),
            .lcout(n13607),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Mux_82_i19_3_lut_LC_24_32_2.C_ON=1'b0;
    defparam Mux_82_i19_3_lut_LC_24_32_2.SEQ_MODE=4'b0000;
    defparam Mux_82_i19_3_lut_LC_24_32_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 Mux_82_i19_3_lut_LC_24_32_2 (
            .in0(N__46412),
            .in1(N__46233),
            .in2(_gnd_net_),
            .in3(N__46227),
            .lcout(n19_adj_789),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
